magic
tech sky130A
magscale 1 2
timestamp 1625353099
<< obsli1 >>
rect 1104 2159 238987 158831
<< obsm1 >>
rect 474 1844 239278 158840
<< metal2 >>
rect 2318 159200 2374 160000
rect 4618 159200 4674 160000
rect 7378 159200 7434 160000
rect 10138 159200 10194 160000
rect 12438 159200 12494 160000
rect 15198 159200 15254 160000
rect 17958 159200 18014 160000
rect 20258 159200 20314 160000
rect 23018 159200 23074 160000
rect 25778 159200 25834 160000
rect 28078 159200 28134 160000
rect 30838 159200 30894 160000
rect 33598 159200 33654 160000
rect 35898 159200 35954 160000
rect 38658 159200 38714 160000
rect 41418 159200 41474 160000
rect 43718 159200 43774 160000
rect 46478 159200 46534 160000
rect 49238 159200 49294 160000
rect 51538 159200 51594 160000
rect 54298 159200 54354 160000
rect 57058 159200 57114 160000
rect 59358 159200 59414 160000
rect 62118 159200 62174 160000
rect 64878 159200 64934 160000
rect 67178 159200 67234 160000
rect 69938 159200 69994 160000
rect 72698 159200 72754 160000
rect 74998 159200 75054 160000
rect 77758 159200 77814 160000
rect 80518 159200 80574 160000
rect 82818 159200 82874 160000
rect 85578 159200 85634 160000
rect 88338 159200 88394 160000
rect 90638 159200 90694 160000
rect 93398 159200 93454 160000
rect 96158 159200 96214 160000
rect 98458 159200 98514 160000
rect 101218 159200 101274 160000
rect 103978 159200 104034 160000
rect 106278 159200 106334 160000
rect 109038 159200 109094 160000
rect 111798 159200 111854 160000
rect 114098 159200 114154 160000
rect 116858 159200 116914 160000
rect 119618 159200 119674 160000
rect 121918 159200 121974 160000
rect 124678 159200 124734 160000
rect 127438 159200 127494 160000
rect 129738 159200 129794 160000
rect 132498 159200 132554 160000
rect 135258 159200 135314 160000
rect 137558 159200 137614 160000
rect 140318 159200 140374 160000
rect 143078 159200 143134 160000
rect 145378 159200 145434 160000
rect 148138 159200 148194 160000
rect 150898 159200 150954 160000
rect 153198 159200 153254 160000
rect 155958 159200 156014 160000
rect 158718 159200 158774 160000
rect 161018 159200 161074 160000
rect 163778 159200 163834 160000
rect 166538 159200 166594 160000
rect 168838 159200 168894 160000
rect 171598 159200 171654 160000
rect 174358 159200 174414 160000
rect 176658 159200 176714 160000
rect 179418 159200 179474 160000
rect 182178 159200 182234 160000
rect 184478 159200 184534 160000
rect 187238 159200 187294 160000
rect 189998 159200 190054 160000
rect 192298 159200 192354 160000
rect 195058 159200 195114 160000
rect 197818 159200 197874 160000
rect 200118 159200 200174 160000
rect 202878 159200 202934 160000
rect 205638 159200 205694 160000
rect 207938 159200 207994 160000
rect 210698 159200 210754 160000
rect 213458 159200 213514 160000
rect 215758 159200 215814 160000
rect 218518 159200 218574 160000
rect 221278 159200 221334 160000
rect 223578 159200 223634 160000
rect 226338 159200 226394 160000
rect 229098 159200 229154 160000
rect 231398 159200 231454 160000
rect 234158 159200 234214 160000
rect 236918 159200 236974 160000
rect 239218 159200 239274 160000
rect 478 0 534 800
rect 2778 0 2834 800
rect 5538 0 5594 800
rect 8298 0 8354 800
rect 10598 0 10654 800
rect 13358 0 13414 800
rect 16118 0 16174 800
rect 18418 0 18474 800
rect 21178 0 21234 800
rect 23938 0 23994 800
rect 26238 0 26294 800
rect 28998 0 29054 800
rect 31758 0 31814 800
rect 34058 0 34114 800
rect 36818 0 36874 800
rect 39578 0 39634 800
rect 41878 0 41934 800
rect 44638 0 44694 800
rect 47398 0 47454 800
rect 49698 0 49754 800
rect 52458 0 52514 800
rect 55218 0 55274 800
rect 57518 0 57574 800
rect 60278 0 60334 800
rect 63038 0 63094 800
rect 65338 0 65394 800
rect 68098 0 68154 800
rect 70858 0 70914 800
rect 73158 0 73214 800
rect 75918 0 75974 800
rect 78678 0 78734 800
rect 80978 0 81034 800
rect 83738 0 83794 800
rect 86498 0 86554 800
rect 88798 0 88854 800
rect 91558 0 91614 800
rect 94318 0 94374 800
rect 96618 0 96674 800
rect 99378 0 99434 800
rect 102138 0 102194 800
rect 104438 0 104494 800
rect 107198 0 107254 800
rect 109958 0 110014 800
rect 112258 0 112314 800
rect 115018 0 115074 800
rect 117778 0 117834 800
rect 120078 0 120134 800
rect 122838 0 122894 800
rect 125598 0 125654 800
rect 127898 0 127954 800
rect 130658 0 130714 800
rect 133418 0 133474 800
rect 135718 0 135774 800
rect 138478 0 138534 800
rect 141238 0 141294 800
rect 143538 0 143594 800
rect 146298 0 146354 800
rect 149058 0 149114 800
rect 151358 0 151414 800
rect 154118 0 154174 800
rect 156878 0 156934 800
rect 159178 0 159234 800
rect 161938 0 161994 800
rect 164698 0 164754 800
rect 166998 0 167054 800
rect 169758 0 169814 800
rect 172518 0 172574 800
rect 174818 0 174874 800
rect 177578 0 177634 800
rect 180338 0 180394 800
rect 182638 0 182694 800
rect 185398 0 185454 800
rect 188158 0 188214 800
rect 190458 0 190514 800
rect 193218 0 193274 800
rect 195978 0 196034 800
rect 198278 0 198334 800
rect 201038 0 201094 800
rect 203798 0 203854 800
rect 206098 0 206154 800
rect 208858 0 208914 800
rect 211618 0 211674 800
rect 213918 0 213974 800
rect 216678 0 216734 800
rect 219438 0 219494 800
rect 221738 0 221794 800
rect 224498 0 224554 800
rect 227258 0 227314 800
rect 229558 0 229614 800
rect 232318 0 232374 800
rect 235078 0 235134 800
rect 237378 0 237434 800
<< obsm2 >>
rect 480 159144 2262 159200
rect 2430 159144 4562 159200
rect 4730 159144 7322 159200
rect 7490 159144 10082 159200
rect 10250 159144 12382 159200
rect 12550 159144 15142 159200
rect 15310 159144 17902 159200
rect 18070 159144 20202 159200
rect 20370 159144 22962 159200
rect 23130 159144 25722 159200
rect 25890 159144 28022 159200
rect 28190 159144 30782 159200
rect 30950 159144 33542 159200
rect 33710 159144 35842 159200
rect 36010 159144 38602 159200
rect 38770 159144 41362 159200
rect 41530 159144 43662 159200
rect 43830 159144 46422 159200
rect 46590 159144 49182 159200
rect 49350 159144 51482 159200
rect 51650 159144 54242 159200
rect 54410 159144 57002 159200
rect 57170 159144 59302 159200
rect 59470 159144 62062 159200
rect 62230 159144 64822 159200
rect 64990 159144 67122 159200
rect 67290 159144 69882 159200
rect 70050 159144 72642 159200
rect 72810 159144 74942 159200
rect 75110 159144 77702 159200
rect 77870 159144 80462 159200
rect 80630 159144 82762 159200
rect 82930 159144 85522 159200
rect 85690 159144 88282 159200
rect 88450 159144 90582 159200
rect 90750 159144 93342 159200
rect 93510 159144 96102 159200
rect 96270 159144 98402 159200
rect 98570 159144 101162 159200
rect 101330 159144 103922 159200
rect 104090 159144 106222 159200
rect 106390 159144 108982 159200
rect 109150 159144 111742 159200
rect 111910 159144 114042 159200
rect 114210 159144 116802 159200
rect 116970 159144 119562 159200
rect 119730 159144 121862 159200
rect 122030 159144 124622 159200
rect 124790 159144 127382 159200
rect 127550 159144 129682 159200
rect 129850 159144 132442 159200
rect 132610 159144 135202 159200
rect 135370 159144 137502 159200
rect 137670 159144 140262 159200
rect 140430 159144 143022 159200
rect 143190 159144 145322 159200
rect 145490 159144 148082 159200
rect 148250 159144 150842 159200
rect 151010 159144 153142 159200
rect 153310 159144 155902 159200
rect 156070 159144 158662 159200
rect 158830 159144 160962 159200
rect 161130 159144 163722 159200
rect 163890 159144 166482 159200
rect 166650 159144 168782 159200
rect 168950 159144 171542 159200
rect 171710 159144 174302 159200
rect 174470 159144 176602 159200
rect 176770 159144 179362 159200
rect 179530 159144 182122 159200
rect 182290 159144 184422 159200
rect 184590 159144 187182 159200
rect 187350 159144 189942 159200
rect 190110 159144 192242 159200
rect 192410 159144 195002 159200
rect 195170 159144 197762 159200
rect 197930 159144 200062 159200
rect 200230 159144 202822 159200
rect 202990 159144 205582 159200
rect 205750 159144 207882 159200
rect 208050 159144 210642 159200
rect 210810 159144 213402 159200
rect 213570 159144 215702 159200
rect 215870 159144 218462 159200
rect 218630 159144 221222 159200
rect 221390 159144 223522 159200
rect 223690 159144 226282 159200
rect 226450 159144 229042 159200
rect 229210 159144 231342 159200
rect 231510 159144 234102 159200
rect 234270 159144 236862 159200
rect 237030 159144 239162 159200
rect 480 856 239272 159144
rect 590 800 2722 856
rect 2890 800 5482 856
rect 5650 800 8242 856
rect 8410 800 10542 856
rect 10710 800 13302 856
rect 13470 800 16062 856
rect 16230 800 18362 856
rect 18530 800 21122 856
rect 21290 800 23882 856
rect 24050 800 26182 856
rect 26350 800 28942 856
rect 29110 800 31702 856
rect 31870 800 34002 856
rect 34170 800 36762 856
rect 36930 800 39522 856
rect 39690 800 41822 856
rect 41990 800 44582 856
rect 44750 800 47342 856
rect 47510 800 49642 856
rect 49810 800 52402 856
rect 52570 800 55162 856
rect 55330 800 57462 856
rect 57630 800 60222 856
rect 60390 800 62982 856
rect 63150 800 65282 856
rect 65450 800 68042 856
rect 68210 800 70802 856
rect 70970 800 73102 856
rect 73270 800 75862 856
rect 76030 800 78622 856
rect 78790 800 80922 856
rect 81090 800 83682 856
rect 83850 800 86442 856
rect 86610 800 88742 856
rect 88910 800 91502 856
rect 91670 800 94262 856
rect 94430 800 96562 856
rect 96730 800 99322 856
rect 99490 800 102082 856
rect 102250 800 104382 856
rect 104550 800 107142 856
rect 107310 800 109902 856
rect 110070 800 112202 856
rect 112370 800 114962 856
rect 115130 800 117722 856
rect 117890 800 120022 856
rect 120190 800 122782 856
rect 122950 800 125542 856
rect 125710 800 127842 856
rect 128010 800 130602 856
rect 130770 800 133362 856
rect 133530 800 135662 856
rect 135830 800 138422 856
rect 138590 800 141182 856
rect 141350 800 143482 856
rect 143650 800 146242 856
rect 146410 800 149002 856
rect 149170 800 151302 856
rect 151470 800 154062 856
rect 154230 800 156822 856
rect 156990 800 159122 856
rect 159290 800 161882 856
rect 162050 800 164642 856
rect 164810 800 166942 856
rect 167110 800 169702 856
rect 169870 800 172462 856
rect 172630 800 174762 856
rect 174930 800 177522 856
rect 177690 800 180282 856
rect 180450 800 182582 856
rect 182750 800 185342 856
rect 185510 800 188102 856
rect 188270 800 190402 856
rect 190570 800 193162 856
rect 193330 800 195922 856
rect 196090 800 198222 856
rect 198390 800 200982 856
rect 201150 800 203742 856
rect 203910 800 206042 856
rect 206210 800 208802 856
rect 208970 800 211562 856
rect 211730 800 213862 856
rect 214030 800 216622 856
rect 216790 800 219382 856
rect 219550 800 221682 856
rect 221850 800 224442 856
rect 224610 800 227202 856
rect 227370 800 229502 856
rect 229670 800 232262 856
rect 232430 800 235022 856
rect 235190 800 237322 856
rect 237490 800 239272 856
<< metal3 >>
rect 0 158448 800 158568
rect 239200 155728 240000 155848
rect 0 154368 800 154488
rect 239200 151648 240000 151768
rect 0 150968 800 151088
rect 239200 147568 240000 147688
rect 0 146888 800 147008
rect 239200 144168 240000 144288
rect 0 142808 800 142928
rect 239200 140088 240000 140208
rect 0 139408 800 139528
rect 239200 136008 240000 136128
rect 0 135328 800 135448
rect 239200 132608 240000 132728
rect 0 131248 800 131368
rect 239200 128528 240000 128648
rect 0 127848 800 127968
rect 239200 124448 240000 124568
rect 0 123768 800 123888
rect 239200 121048 240000 121168
rect 0 119688 800 119808
rect 239200 116968 240000 117088
rect 0 116288 800 116408
rect 239200 112888 240000 113008
rect 0 112208 800 112328
rect 239200 109488 240000 109608
rect 0 108128 800 108248
rect 239200 105408 240000 105528
rect 0 104728 800 104848
rect 239200 101328 240000 101448
rect 0 100648 800 100768
rect 239200 97928 240000 98048
rect 0 96568 800 96688
rect 239200 93848 240000 93968
rect 0 93168 800 93288
rect 239200 89768 240000 89888
rect 0 89088 800 89208
rect 239200 86368 240000 86488
rect 0 85008 800 85128
rect 239200 82288 240000 82408
rect 0 81608 800 81728
rect 239200 78208 240000 78328
rect 0 77528 800 77648
rect 239200 74808 240000 74928
rect 0 73448 800 73568
rect 239200 70728 240000 70848
rect 0 70048 800 70168
rect 239200 66648 240000 66768
rect 0 65968 800 66088
rect 239200 63248 240000 63368
rect 0 61888 800 62008
rect 239200 59168 240000 59288
rect 0 58488 800 58608
rect 239200 55088 240000 55208
rect 0 54408 800 54528
rect 239200 51688 240000 51808
rect 0 50328 800 50448
rect 239200 47608 240000 47728
rect 0 46928 800 47048
rect 239200 43528 240000 43648
rect 0 42848 800 42968
rect 239200 40128 240000 40248
rect 0 38768 800 38888
rect 239200 36048 240000 36168
rect 0 35368 800 35488
rect 239200 31968 240000 32088
rect 0 31288 800 31408
rect 239200 28568 240000 28688
rect 0 27208 800 27328
rect 239200 24488 240000 24608
rect 0 23808 800 23928
rect 239200 20408 240000 20528
rect 0 19728 800 19848
rect 239200 17008 240000 17128
rect 0 15648 800 15768
rect 239200 12928 240000 13048
rect 0 12248 800 12368
rect 239200 8848 240000 8968
rect 0 8168 800 8288
rect 239200 5448 240000 5568
rect 0 4088 800 4208
rect 239200 1368 240000 1488
<< obsm3 >>
rect 880 158368 239200 158541
rect 800 155928 239200 158368
rect 800 155648 239120 155928
rect 800 154568 239200 155648
rect 880 154288 239200 154568
rect 800 151848 239200 154288
rect 800 151568 239120 151848
rect 800 151168 239200 151568
rect 880 150888 239200 151168
rect 800 147768 239200 150888
rect 800 147488 239120 147768
rect 800 147088 239200 147488
rect 880 146808 239200 147088
rect 800 144368 239200 146808
rect 800 144088 239120 144368
rect 800 143008 239200 144088
rect 880 142728 239200 143008
rect 800 140288 239200 142728
rect 800 140008 239120 140288
rect 800 139608 239200 140008
rect 880 139328 239200 139608
rect 800 136208 239200 139328
rect 800 135928 239120 136208
rect 800 135528 239200 135928
rect 880 135248 239200 135528
rect 800 132808 239200 135248
rect 800 132528 239120 132808
rect 800 131448 239200 132528
rect 880 131168 239200 131448
rect 800 128728 239200 131168
rect 800 128448 239120 128728
rect 800 128048 239200 128448
rect 880 127768 239200 128048
rect 800 124648 239200 127768
rect 800 124368 239120 124648
rect 800 123968 239200 124368
rect 880 123688 239200 123968
rect 800 121248 239200 123688
rect 800 120968 239120 121248
rect 800 119888 239200 120968
rect 880 119608 239200 119888
rect 800 117168 239200 119608
rect 800 116888 239120 117168
rect 800 116488 239200 116888
rect 880 116208 239200 116488
rect 800 113088 239200 116208
rect 800 112808 239120 113088
rect 800 112408 239200 112808
rect 880 112128 239200 112408
rect 800 109688 239200 112128
rect 800 109408 239120 109688
rect 800 108328 239200 109408
rect 880 108048 239200 108328
rect 800 105608 239200 108048
rect 800 105328 239120 105608
rect 800 104928 239200 105328
rect 880 104648 239200 104928
rect 800 101528 239200 104648
rect 800 101248 239120 101528
rect 800 100848 239200 101248
rect 880 100568 239200 100848
rect 800 98128 239200 100568
rect 800 97848 239120 98128
rect 800 96768 239200 97848
rect 880 96488 239200 96768
rect 800 94048 239200 96488
rect 800 93768 239120 94048
rect 800 93368 239200 93768
rect 880 93088 239200 93368
rect 800 89968 239200 93088
rect 800 89688 239120 89968
rect 800 89288 239200 89688
rect 880 89008 239200 89288
rect 800 86568 239200 89008
rect 800 86288 239120 86568
rect 800 85208 239200 86288
rect 880 84928 239200 85208
rect 800 82488 239200 84928
rect 800 82208 239120 82488
rect 800 81808 239200 82208
rect 880 81528 239200 81808
rect 800 78408 239200 81528
rect 800 78128 239120 78408
rect 800 77728 239200 78128
rect 880 77448 239200 77728
rect 800 75008 239200 77448
rect 800 74728 239120 75008
rect 800 73648 239200 74728
rect 880 73368 239200 73648
rect 800 70928 239200 73368
rect 800 70648 239120 70928
rect 800 70248 239200 70648
rect 880 69968 239200 70248
rect 800 66848 239200 69968
rect 800 66568 239120 66848
rect 800 66168 239200 66568
rect 880 65888 239200 66168
rect 800 63448 239200 65888
rect 800 63168 239120 63448
rect 800 62088 239200 63168
rect 880 61808 239200 62088
rect 800 59368 239200 61808
rect 800 59088 239120 59368
rect 800 58688 239200 59088
rect 880 58408 239200 58688
rect 800 55288 239200 58408
rect 800 55008 239120 55288
rect 800 54608 239200 55008
rect 880 54328 239200 54608
rect 800 51888 239200 54328
rect 800 51608 239120 51888
rect 800 50528 239200 51608
rect 880 50248 239200 50528
rect 800 47808 239200 50248
rect 800 47528 239120 47808
rect 800 47128 239200 47528
rect 880 46848 239200 47128
rect 800 43728 239200 46848
rect 800 43448 239120 43728
rect 800 43048 239200 43448
rect 880 42768 239200 43048
rect 800 40328 239200 42768
rect 800 40048 239120 40328
rect 800 38968 239200 40048
rect 880 38688 239200 38968
rect 800 36248 239200 38688
rect 800 35968 239120 36248
rect 800 35568 239200 35968
rect 880 35288 239200 35568
rect 800 32168 239200 35288
rect 800 31888 239120 32168
rect 800 31488 239200 31888
rect 880 31208 239200 31488
rect 800 28768 239200 31208
rect 800 28488 239120 28768
rect 800 27408 239200 28488
rect 880 27128 239200 27408
rect 800 24688 239200 27128
rect 800 24408 239120 24688
rect 800 24008 239200 24408
rect 880 23728 239200 24008
rect 800 20608 239200 23728
rect 800 20328 239120 20608
rect 800 19928 239200 20328
rect 880 19648 239200 19928
rect 800 17208 239200 19648
rect 800 16928 239120 17208
rect 800 15848 239200 16928
rect 880 15568 239200 15848
rect 800 13128 239200 15568
rect 800 12848 239120 13128
rect 800 12448 239200 12848
rect 880 12168 239200 12448
rect 800 9048 239200 12168
rect 800 8768 239120 9048
rect 800 8368 239200 8768
rect 880 8088 239200 8368
rect 800 5648 239200 8088
rect 800 5368 239120 5648
rect 800 4288 239200 5368
rect 880 4008 239200 4288
rect 800 1568 239200 4008
rect 800 1395 239120 1568
<< metal4 >>
rect 4208 2128 4528 157808
rect 9208 2128 9528 157808
rect 14208 95452 14528 157808
rect 19208 95452 19528 157808
rect 24208 95452 24528 157808
rect 29208 95452 29528 157808
rect 34208 95452 34528 157808
rect 39208 95452 39528 157808
rect 44208 95452 44528 157808
rect 49208 95452 49528 157808
rect 54208 95452 54528 157808
rect 59208 95452 59528 157808
rect 64208 95452 64528 157808
rect 69208 95452 69528 157808
rect 74208 95452 74528 157808
rect 79208 95452 79528 157808
rect 84208 95452 84528 157808
rect 89208 95452 89528 157808
rect 94208 95452 94528 157808
rect 99208 95452 99528 157808
rect 104208 95452 104528 157808
rect 109208 95452 109528 157808
rect 14208 2128 14528 14048
rect 19208 2128 19528 14048
rect 24208 2128 24528 14048
rect 29208 2128 29528 14048
rect 34208 2128 34528 14048
rect 39208 2128 39528 14048
rect 44208 2128 44528 14048
rect 49208 2128 49528 14048
rect 54208 2128 54528 14048
rect 59208 2128 59528 14048
rect 64208 2128 64528 14048
rect 69208 2128 69528 14048
rect 74208 2128 74528 14048
rect 79208 2128 79528 14048
rect 84208 2128 84528 14048
rect 89208 2128 89528 14048
rect 94208 2128 94528 14048
rect 99208 2128 99528 14048
rect 104208 2128 104528 14048
rect 109208 2128 109528 14048
rect 114208 2128 114528 157808
rect 119208 2128 119528 157808
rect 124208 2128 124528 157808
rect 129208 2128 129528 157808
rect 134208 2128 134528 157808
rect 139208 2128 139528 157808
rect 144208 2128 144528 157808
rect 149208 2128 149528 157808
rect 154208 2128 154528 157808
rect 159208 2128 159528 157808
rect 164208 2128 164528 157808
rect 169208 2128 169528 157808
rect 174208 2128 174528 157808
rect 179208 2128 179528 157808
rect 184208 2128 184528 157808
rect 189208 2128 189528 157808
rect 194208 2128 194528 157808
rect 199208 2128 199528 157808
rect 204208 2128 204528 157808
rect 209208 2128 209528 157808
rect 214208 2128 214528 157808
rect 219208 2128 219528 157808
rect 224208 2128 224528 157808
rect 229208 2128 229528 157808
rect 234208 2128 234528 157808
<< obsm4 >>
rect 1998 2347 4128 157589
rect 4608 2347 9128 157589
rect 9608 95372 14128 157589
rect 14608 95372 19128 157589
rect 19608 95372 24128 157589
rect 24608 95372 29128 157589
rect 29608 95372 34128 157589
rect 34608 95372 39128 157589
rect 39608 95372 44128 157589
rect 44608 95372 49128 157589
rect 49608 95372 54128 157589
rect 54608 95372 59128 157589
rect 59608 95372 64128 157589
rect 64608 95372 69128 157589
rect 69608 95372 74128 157589
rect 74608 95372 79128 157589
rect 79608 95372 84128 157589
rect 84608 95372 89128 157589
rect 89608 95372 94128 157589
rect 94608 95372 99128 157589
rect 99608 95372 104128 157589
rect 104608 95372 109128 157589
rect 109608 95372 114128 157589
rect 9608 14128 114128 95372
rect 9608 2347 14128 14128
rect 14608 2347 19128 14128
rect 19608 2347 24128 14128
rect 24608 2347 29128 14128
rect 29608 2347 34128 14128
rect 34608 2347 39128 14128
rect 39608 2347 44128 14128
rect 44608 2347 49128 14128
rect 49608 2347 54128 14128
rect 54608 2347 59128 14128
rect 59608 2347 64128 14128
rect 64608 2347 69128 14128
rect 69608 2347 74128 14128
rect 74608 2347 79128 14128
rect 79608 2347 84128 14128
rect 84608 2347 89128 14128
rect 89608 2347 94128 14128
rect 94608 2347 99128 14128
rect 99608 2347 104128 14128
rect 104608 2347 109128 14128
rect 109608 2347 114128 14128
rect 114608 2347 119128 157589
rect 119608 2347 124128 157589
rect 124608 2347 129128 157589
rect 129608 2347 134128 157589
rect 134608 2347 139128 157589
rect 139608 2347 144128 157589
rect 144608 2347 149128 157589
rect 149608 2347 154128 157589
rect 154608 2347 159128 157589
rect 159608 2347 164128 157589
rect 164608 2347 169128 157589
rect 169608 2347 174128 157589
rect 174608 2347 179128 157589
rect 179608 2347 184128 157589
rect 184608 2347 189128 157589
rect 189608 2347 194128 157589
rect 194608 2347 199128 157589
rect 199608 2347 204128 157589
rect 204608 2347 209128 157589
rect 209608 2347 214128 157589
rect 214608 2347 219128 157589
rect 219608 2347 224128 157589
rect 224608 2347 229128 157589
rect 229608 2347 234128 157589
rect 234608 2347 236098 157589
<< metal5 >>
rect 1104 143160 238832 143480
rect 1104 127842 238832 128162
rect 1104 112524 238832 112844
rect 1104 97206 238832 97526
rect 1104 81888 238832 82208
rect 1104 66570 238832 66890
rect 1104 51252 238832 51572
rect 1104 35934 238832 36254
rect 1104 20616 238832 20936
rect 1104 5298 238832 5618
<< obsm5 >>
rect 1956 82528 236140 95020
rect 1956 67210 236140 81568
rect 1956 51892 236140 66250
rect 1956 36574 236140 50932
rect 1956 21256 236140 35614
rect 1956 14460 236140 20296
<< labels >>
rlabel metal2 s 232318 0 232374 800 6 clk_i
port 1 nsew signal input
rlabel metal3 s 239200 147568 240000 147688 6 debug_req_i
port 2 nsew signal input
rlabel metal2 s 205638 159200 205694 160000 6 eFPGA_delay_o[0]
port 3 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 eFPGA_delay_o[1]
port 4 nsew signal output
rlabel metal2 s 224498 0 224554 800 6 eFPGA_delay_o[2]
port 5 nsew signal output
rlabel metal2 s 148138 159200 148194 160000 6 eFPGA_delay_o[3]
port 6 nsew signal output
rlabel metal2 s 69938 159200 69994 160000 6 eFPGA_en_o
port 7 nsew signal output
rlabel metal2 s 96618 0 96674 800 6 eFPGA_fpga_done_i
port 8 nsew signal input
rlabel metal3 s 239200 140088 240000 140208 6 eFPGA_operand_a_o[0]
port 9 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 eFPGA_operand_a_o[10]
port 10 nsew signal output
rlabel metal3 s 0 131248 800 131368 6 eFPGA_operand_a_o[11]
port 11 nsew signal output
rlabel metal2 s 219438 0 219494 800 6 eFPGA_operand_a_o[12]
port 12 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 eFPGA_operand_a_o[13]
port 13 nsew signal output
rlabel metal2 s 138478 0 138534 800 6 eFPGA_operand_a_o[14]
port 14 nsew signal output
rlabel metal2 s 200118 159200 200174 160000 6 eFPGA_operand_a_o[15]
port 15 nsew signal output
rlabel metal3 s 239200 74808 240000 74928 6 eFPGA_operand_a_o[16]
port 16 nsew signal output
rlabel metal2 s 176658 159200 176714 160000 6 eFPGA_operand_a_o[17]
port 17 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 eFPGA_operand_a_o[18]
port 18 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 eFPGA_operand_a_o[19]
port 19 nsew signal output
rlabel metal2 s 2318 159200 2374 160000 6 eFPGA_operand_a_o[1]
port 20 nsew signal output
rlabel metal2 s 46478 159200 46534 160000 6 eFPGA_operand_a_o[20]
port 21 nsew signal output
rlabel metal3 s 239200 124448 240000 124568 6 eFPGA_operand_a_o[21]
port 22 nsew signal output
rlabel metal3 s 239200 8848 240000 8968 6 eFPGA_operand_a_o[22]
port 23 nsew signal output
rlabel metal3 s 239200 20408 240000 20528 6 eFPGA_operand_a_o[23]
port 24 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 eFPGA_operand_a_o[24]
port 25 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 eFPGA_operand_a_o[25]
port 26 nsew signal output
rlabel metal2 s 234158 159200 234214 160000 6 eFPGA_operand_a_o[26]
port 27 nsew signal output
rlabel metal2 s 239218 159200 239274 160000 6 eFPGA_operand_a_o[27]
port 28 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 eFPGA_operand_a_o[28]
port 29 nsew signal output
rlabel metal2 s 143078 159200 143134 160000 6 eFPGA_operand_a_o[29]
port 30 nsew signal output
rlabel metal3 s 239200 36048 240000 36168 6 eFPGA_operand_a_o[2]
port 31 nsew signal output
rlabel metal2 s 188158 0 188214 800 6 eFPGA_operand_a_o[30]
port 32 nsew signal output
rlabel metal2 s 121918 159200 121974 160000 6 eFPGA_operand_a_o[31]
port 33 nsew signal output
rlabel metal2 s 213918 0 213974 800 6 eFPGA_operand_a_o[3]
port 34 nsew signal output
rlabel metal2 s 195058 159200 195114 160000 6 eFPGA_operand_a_o[4]
port 35 nsew signal output
rlabel metal3 s 0 42848 800 42968 6 eFPGA_operand_a_o[5]
port 36 nsew signal output
rlabel metal2 s 74998 159200 75054 160000 6 eFPGA_operand_a_o[6]
port 37 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 eFPGA_operand_a_o[7]
port 38 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 eFPGA_operand_a_o[8]
port 39 nsew signal output
rlabel metal2 s 90638 159200 90694 160000 6 eFPGA_operand_a_o[9]
port 40 nsew signal output
rlabel metal2 s 229098 159200 229154 160000 6 eFPGA_operand_b_o[0]
port 41 nsew signal output
rlabel metal2 s 223578 159200 223634 160000 6 eFPGA_operand_b_o[10]
port 42 nsew signal output
rlabel metal2 s 109038 159200 109094 160000 6 eFPGA_operand_b_o[11]
port 43 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 eFPGA_operand_b_o[12]
port 44 nsew signal output
rlabel metal3 s 0 146888 800 147008 6 eFPGA_operand_b_o[13]
port 45 nsew signal output
rlabel metal2 s 127438 159200 127494 160000 6 eFPGA_operand_b_o[14]
port 46 nsew signal output
rlabel metal2 s 67178 159200 67234 160000 6 eFPGA_operand_b_o[15]
port 47 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 eFPGA_operand_b_o[16]
port 48 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 eFPGA_operand_b_o[17]
port 49 nsew signal output
rlabel metal2 s 208858 0 208914 800 6 eFPGA_operand_b_o[18]
port 50 nsew signal output
rlabel metal2 s 25778 159200 25834 160000 6 eFPGA_operand_b_o[19]
port 51 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 eFPGA_operand_b_o[1]
port 52 nsew signal output
rlabel metal2 s 80978 0 81034 800 6 eFPGA_operand_b_o[20]
port 53 nsew signal output
rlabel metal3 s 239200 86368 240000 86488 6 eFPGA_operand_b_o[21]
port 54 nsew signal output
rlabel metal2 s 135258 159200 135314 160000 6 eFPGA_operand_b_o[22]
port 55 nsew signal output
rlabel metal2 s 93398 159200 93454 160000 6 eFPGA_operand_b_o[23]
port 56 nsew signal output
rlabel metal2 s 182178 159200 182234 160000 6 eFPGA_operand_b_o[24]
port 57 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 eFPGA_operand_b_o[25]
port 58 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 eFPGA_operand_b_o[26]
port 59 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 eFPGA_operand_b_o[27]
port 60 nsew signal output
rlabel metal2 s 15198 159200 15254 160000 6 eFPGA_operand_b_o[28]
port 61 nsew signal output
rlabel metal2 s 156878 0 156934 800 6 eFPGA_operand_b_o[29]
port 62 nsew signal output
rlabel metal3 s 239200 112888 240000 113008 6 eFPGA_operand_b_o[2]
port 63 nsew signal output
rlabel metal3 s 239200 40128 240000 40248 6 eFPGA_operand_b_o[30]
port 64 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 eFPGA_operand_b_o[31]
port 65 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 eFPGA_operand_b_o[3]
port 66 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 eFPGA_operand_b_o[4]
port 67 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 eFPGA_operand_b_o[5]
port 68 nsew signal output
rlabel metal2 s 132498 159200 132554 160000 6 eFPGA_operand_b_o[6]
port 69 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 eFPGA_operand_b_o[7]
port 70 nsew signal output
rlabel metal2 s 161018 159200 161074 160000 6 eFPGA_operand_b_o[8]
port 71 nsew signal output
rlabel metal2 s 177578 0 177634 800 6 eFPGA_operand_b_o[9]
port 72 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 eFPGA_operator_o[0]
port 73 nsew signal output
rlabel metal3 s 239200 109488 240000 109608 6 eFPGA_operator_o[1]
port 74 nsew signal output
rlabel metal2 s 41418 159200 41474 160000 6 eFPGA_result_a_i[0]
port 75 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 eFPGA_result_a_i[10]
port 76 nsew signal input
rlabel metal2 s 129738 159200 129794 160000 6 eFPGA_result_a_i[11]
port 77 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 eFPGA_result_a_i[12]
port 78 nsew signal input
rlabel metal2 s 226338 159200 226394 160000 6 eFPGA_result_a_i[13]
port 79 nsew signal input
rlabel metal2 s 35898 159200 35954 160000 6 eFPGA_result_a_i[14]
port 80 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 eFPGA_result_a_i[15]
port 81 nsew signal input
rlabel metal2 s 158718 159200 158774 160000 6 eFPGA_result_a_i[16]
port 82 nsew signal input
rlabel metal2 s 72698 159200 72754 160000 6 eFPGA_result_a_i[17]
port 83 nsew signal input
rlabel metal2 s 38658 159200 38714 160000 6 eFPGA_result_a_i[18]
port 84 nsew signal input
rlabel metal3 s 239200 121048 240000 121168 6 eFPGA_result_a_i[19]
port 85 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 eFPGA_result_a_i[1]
port 86 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 eFPGA_result_a_i[20]
port 87 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 eFPGA_result_a_i[21]
port 88 nsew signal input
rlabel metal2 s 235078 0 235134 800 6 eFPGA_result_a_i[22]
port 89 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 eFPGA_result_a_i[23]
port 90 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 eFPGA_result_a_i[24]
port 91 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 eFPGA_result_a_i[25]
port 92 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 eFPGA_result_a_i[26]
port 93 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 eFPGA_result_a_i[27]
port 94 nsew signal input
rlabel metal2 s 98458 159200 98514 160000 6 eFPGA_result_a_i[28]
port 95 nsew signal input
rlabel metal2 s 146298 0 146354 800 6 eFPGA_result_a_i[29]
port 96 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 eFPGA_result_a_i[2]
port 97 nsew signal input
rlabel metal3 s 239200 151648 240000 151768 6 eFPGA_result_a_i[30]
port 98 nsew signal input
rlabel metal2 s 96158 159200 96214 160000 6 eFPGA_result_a_i[31]
port 99 nsew signal input
rlabel metal2 s 163778 159200 163834 160000 6 eFPGA_result_a_i[3]
port 100 nsew signal input
rlabel metal2 s 82818 159200 82874 160000 6 eFPGA_result_a_i[4]
port 101 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 eFPGA_result_a_i[5]
port 102 nsew signal input
rlabel metal2 s 171598 159200 171654 160000 6 eFPGA_result_a_i[6]
port 103 nsew signal input
rlabel metal2 s 70858 0 70914 800 6 eFPGA_result_a_i[7]
port 104 nsew signal input
rlabel metal2 s 189998 159200 190054 160000 6 eFPGA_result_a_i[8]
port 105 nsew signal input
rlabel metal2 s 85578 159200 85634 160000 6 eFPGA_result_a_i[9]
port 106 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 eFPGA_result_b_i[0]
port 107 nsew signal input
rlabel metal3 s 239200 82288 240000 82408 6 eFPGA_result_b_i[10]
port 108 nsew signal input
rlabel metal2 s 174358 159200 174414 160000 6 eFPGA_result_b_i[11]
port 109 nsew signal input
rlabel metal3 s 239200 70728 240000 70848 6 eFPGA_result_b_i[12]
port 110 nsew signal input
rlabel metal2 s 80518 159200 80574 160000 6 eFPGA_result_b_i[13]
port 111 nsew signal input
rlabel metal2 s 119618 159200 119674 160000 6 eFPGA_result_b_i[14]
port 112 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 eFPGA_result_b_i[15]
port 113 nsew signal input
rlabel metal2 s 221278 159200 221334 160000 6 eFPGA_result_b_i[16]
port 114 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 eFPGA_result_b_i[17]
port 115 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 eFPGA_result_b_i[18]
port 116 nsew signal input
rlabel metal2 s 155958 159200 156014 160000 6 eFPGA_result_b_i[19]
port 117 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 eFPGA_result_b_i[1]
port 118 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 eFPGA_result_b_i[20]
port 119 nsew signal input
rlabel metal2 s 116858 159200 116914 160000 6 eFPGA_result_b_i[21]
port 120 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 eFPGA_result_b_i[22]
port 121 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 eFPGA_result_b_i[23]
port 122 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 eFPGA_result_b_i[24]
port 123 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 eFPGA_result_b_i[25]
port 124 nsew signal input
rlabel metal2 s 103978 159200 104034 160000 6 eFPGA_result_b_i[26]
port 125 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 eFPGA_result_b_i[27]
port 126 nsew signal input
rlabel metal3 s 239200 155728 240000 155848 6 eFPGA_result_b_i[28]
port 127 nsew signal input
rlabel metal2 s 236918 159200 236974 160000 6 eFPGA_result_b_i[29]
port 128 nsew signal input
rlabel metal2 s 30838 159200 30894 160000 6 eFPGA_result_b_i[2]
port 129 nsew signal input
rlabel metal3 s 0 154368 800 154488 6 eFPGA_result_b_i[30]
port 130 nsew signal input
rlabel metal2 s 193218 0 193274 800 6 eFPGA_result_b_i[31]
port 131 nsew signal input
rlabel metal2 s 192298 159200 192354 160000 6 eFPGA_result_b_i[3]
port 132 nsew signal input
rlabel metal2 s 231398 159200 231454 160000 6 eFPGA_result_b_i[4]
port 133 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 eFPGA_result_b_i[5]
port 134 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 eFPGA_result_b_i[6]
port 135 nsew signal input
rlabel metal2 s 229558 0 229614 800 6 eFPGA_result_b_i[7]
port 136 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 eFPGA_result_b_i[8]
port 137 nsew signal input
rlabel metal2 s 77758 159200 77814 160000 6 eFPGA_result_b_i[9]
port 138 nsew signal input
rlabel metal2 s 111798 159200 111854 160000 6 eFPGA_result_c_i[0]
port 139 nsew signal input
rlabel metal2 s 153198 159200 153254 160000 6 eFPGA_result_c_i[10]
port 140 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 eFPGA_result_c_i[11]
port 141 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 eFPGA_result_c_i[12]
port 142 nsew signal input
rlabel metal2 s 195978 0 196034 800 6 eFPGA_result_c_i[13]
port 143 nsew signal input
rlabel metal2 s 124678 159200 124734 160000 6 eFPGA_result_c_i[14]
port 144 nsew signal input
rlabel metal3 s 239200 17008 240000 17128 6 eFPGA_result_c_i[15]
port 145 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 eFPGA_result_c_i[16]
port 146 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 eFPGA_result_c_i[17]
port 147 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 eFPGA_result_c_i[18]
port 148 nsew signal input
rlabel metal2 s 180338 0 180394 800 6 eFPGA_result_c_i[19]
port 149 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 eFPGA_result_c_i[1]
port 150 nsew signal input
rlabel metal3 s 239200 1368 240000 1488 6 eFPGA_result_c_i[20]
port 151 nsew signal input
rlabel metal3 s 239200 28568 240000 28688 6 eFPGA_result_c_i[21]
port 152 nsew signal input
rlabel metal2 s 478 0 534 800 6 eFPGA_result_c_i[22]
port 153 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 eFPGA_result_c_i[23]
port 154 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 eFPGA_result_c_i[24]
port 155 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 eFPGA_result_c_i[25]
port 156 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 eFPGA_result_c_i[26]
port 157 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 eFPGA_result_c_i[27]
port 158 nsew signal input
rlabel metal2 s 54298 159200 54354 160000 6 eFPGA_result_c_i[28]
port 159 nsew signal input
rlabel metal2 s 17958 159200 18014 160000 6 eFPGA_result_c_i[29]
port 160 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 eFPGA_result_c_i[2]
port 161 nsew signal input
rlabel metal2 s 187238 159200 187294 160000 6 eFPGA_result_c_i[30]
port 162 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 eFPGA_result_c_i[31]
port 163 nsew signal input
rlabel metal2 s 10138 159200 10194 160000 6 eFPGA_result_c_i[3]
port 164 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 eFPGA_result_c_i[4]
port 165 nsew signal input
rlabel metal3 s 239200 66648 240000 66768 6 eFPGA_result_c_i[5]
port 166 nsew signal input
rlabel metal2 s 114098 159200 114154 160000 6 eFPGA_result_c_i[6]
port 167 nsew signal input
rlabel metal2 s 207938 159200 207994 160000 6 eFPGA_result_c_i[7]
port 168 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 eFPGA_result_c_i[8]
port 169 nsew signal input
rlabel metal3 s 239200 55088 240000 55208 6 eFPGA_result_c_i[9]
port 170 nsew signal input
rlabel metal2 s 59358 159200 59414 160000 6 eFPGA_write_strobe_o
port 171 nsew signal output
rlabel metal2 s 216678 0 216734 800 6 ext_data_addr_i[0]
port 172 nsew signal input
rlabel metal2 s 213458 159200 213514 160000 6 ext_data_addr_i[1]
port 173 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 ext_data_addr_i[2]
port 174 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 ext_data_addr_i[3]
port 175 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 ext_data_addr_i[4]
port 176 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 ext_data_addr_i[5]
port 177 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 ext_data_addr_i[6]
port 178 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 ext_data_addr_i[7]
port 179 nsew signal input
rlabel metal2 s 62118 159200 62174 160000 6 ext_data_addr_i[8]
port 180 nsew signal input
rlabel metal2 s 190458 0 190514 800 6 ext_data_addr_i[9]
port 181 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 ext_data_be_i[0]
port 182 nsew signal input
rlabel metal3 s 239200 89768 240000 89888 6 ext_data_be_i[1]
port 183 nsew signal input
rlabel metal2 s 4618 159200 4674 160000 6 ext_data_be_i[2]
port 184 nsew signal input
rlabel metal3 s 239200 132608 240000 132728 6 ext_data_be_i[3]
port 185 nsew signal input
rlabel metal2 s 51538 159200 51594 160000 6 ext_data_rdata_o[0]
port 186 nsew signal output
rlabel metal3 s 239200 31968 240000 32088 6 ext_data_rdata_o[10]
port 187 nsew signal output
rlabel metal2 s 198278 0 198334 800 6 ext_data_rdata_o[11]
port 188 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 ext_data_rdata_o[12]
port 189 nsew signal output
rlabel metal2 s 215758 159200 215814 160000 6 ext_data_rdata_o[13]
port 190 nsew signal output
rlabel metal2 s 33598 159200 33654 160000 6 ext_data_rdata_o[14]
port 191 nsew signal output
rlabel metal2 s 145378 159200 145434 160000 6 ext_data_rdata_o[15]
port 192 nsew signal output
rlabel metal2 s 166538 159200 166594 160000 6 ext_data_rdata_o[16]
port 193 nsew signal output
rlabel metal2 s 185398 0 185454 800 6 ext_data_rdata_o[17]
port 194 nsew signal output
rlabel metal2 s 64878 159200 64934 160000 6 ext_data_rdata_o[18]
port 195 nsew signal output
rlabel metal2 s 88338 159200 88394 160000 6 ext_data_rdata_o[19]
port 196 nsew signal output
rlabel metal2 s 43718 159200 43774 160000 6 ext_data_rdata_o[1]
port 197 nsew signal output
rlabel metal2 s 197818 159200 197874 160000 6 ext_data_rdata_o[20]
port 198 nsew signal output
rlabel metal3 s 239200 5448 240000 5568 6 ext_data_rdata_o[21]
port 199 nsew signal output
rlabel metal2 s 28078 159200 28134 160000 6 ext_data_rdata_o[22]
port 200 nsew signal output
rlabel metal2 s 57058 159200 57114 160000 6 ext_data_rdata_o[23]
port 201 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 ext_data_rdata_o[24]
port 202 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 ext_data_rdata_o[25]
port 203 nsew signal output
rlabel metal2 s 12438 159200 12494 160000 6 ext_data_rdata_o[26]
port 204 nsew signal output
rlabel metal2 s 237378 0 237434 800 6 ext_data_rdata_o[27]
port 205 nsew signal output
rlabel metal3 s 0 158448 800 158568 6 ext_data_rdata_o[28]
port 206 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 ext_data_rdata_o[29]
port 207 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 ext_data_rdata_o[2]
port 208 nsew signal output
rlabel metal2 s 206098 0 206154 800 6 ext_data_rdata_o[30]
port 209 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 ext_data_rdata_o[31]
port 210 nsew signal output
rlabel metal3 s 239200 116968 240000 117088 6 ext_data_rdata_o[3]
port 211 nsew signal output
rlabel metal2 s 101218 159200 101274 160000 6 ext_data_rdata_o[4]
port 212 nsew signal output
rlabel metal3 s 239200 128528 240000 128648 6 ext_data_rdata_o[5]
port 213 nsew signal output
rlabel metal3 s 239200 24488 240000 24608 6 ext_data_rdata_o[6]
port 214 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 ext_data_rdata_o[7]
port 215 nsew signal output
rlabel metal3 s 239200 144168 240000 144288 6 ext_data_rdata_o[8]
port 216 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 ext_data_rdata_o[9]
port 217 nsew signal output
rlabel metal3 s 239200 59168 240000 59288 6 ext_data_req_i
port 218 nsew signal input
rlabel metal3 s 239200 101328 240000 101448 6 ext_data_rvalid_o
port 219 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 ext_data_wdata_i[0]
port 220 nsew signal input
rlabel metal2 s 227258 0 227314 800 6 ext_data_wdata_i[10]
port 221 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 ext_data_wdata_i[11]
port 222 nsew signal input
rlabel metal3 s 239200 43528 240000 43648 6 ext_data_wdata_i[12]
port 223 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 ext_data_wdata_i[13]
port 224 nsew signal input
rlabel metal2 s 168838 159200 168894 160000 6 ext_data_wdata_i[14]
port 225 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 ext_data_wdata_i[15]
port 226 nsew signal input
rlabel metal2 s 23018 159200 23074 160000 6 ext_data_wdata_i[16]
port 227 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 ext_data_wdata_i[17]
port 228 nsew signal input
rlabel metal2 s 210698 159200 210754 160000 6 ext_data_wdata_i[18]
port 229 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 ext_data_wdata_i[19]
port 230 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 ext_data_wdata_i[1]
port 231 nsew signal input
rlabel metal2 s 7378 159200 7434 160000 6 ext_data_wdata_i[20]
port 232 nsew signal input
rlabel metal3 s 239200 12928 240000 13048 6 ext_data_wdata_i[21]
port 233 nsew signal input
rlabel metal3 s 239200 105408 240000 105528 6 ext_data_wdata_i[22]
port 234 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 ext_data_wdata_i[23]
port 235 nsew signal input
rlabel metal3 s 239200 47608 240000 47728 6 ext_data_wdata_i[24]
port 236 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 ext_data_wdata_i[25]
port 237 nsew signal input
rlabel metal2 s 150898 159200 150954 160000 6 ext_data_wdata_i[26]
port 238 nsew signal input
rlabel metal2 s 140318 159200 140374 160000 6 ext_data_wdata_i[27]
port 239 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 ext_data_wdata_i[28]
port 240 nsew signal input
rlabel metal2 s 49238 159200 49294 160000 6 ext_data_wdata_i[29]
port 241 nsew signal input
rlabel metal2 s 20258 159200 20314 160000 6 ext_data_wdata_i[2]
port 242 nsew signal input
rlabel metal2 s 218518 159200 218574 160000 6 ext_data_wdata_i[30]
port 243 nsew signal input
rlabel metal2 s 143538 0 143594 800 6 ext_data_wdata_i[31]
port 244 nsew signal input
rlabel metal3 s 239200 78208 240000 78328 6 ext_data_wdata_i[3]
port 245 nsew signal input
rlabel metal3 s 239200 51688 240000 51808 6 ext_data_wdata_i[4]
port 246 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 ext_data_wdata_i[5]
port 247 nsew signal input
rlabel metal2 s 109958 0 110014 800 6 ext_data_wdata_i[6]
port 248 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 ext_data_wdata_i[7]
port 249 nsew signal input
rlabel metal2 s 182638 0 182694 800 6 ext_data_wdata_i[8]
port 250 nsew signal input
rlabel metal3 s 239200 97928 240000 98048 6 ext_data_wdata_i[9]
port 251 nsew signal input
rlabel metal2 s 179418 159200 179474 160000 6 ext_data_we_i
port 252 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 fetch_enable_i
port 253 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 irq_ack_o
port 254 nsew signal output
rlabel metal3 s 239200 136008 240000 136128 6 irq_i
port 255 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 irq_id_i[0]
port 256 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 irq_id_i[1]
port 257 nsew signal input
rlabel metal2 s 202878 159200 202934 160000 6 irq_id_i[2]
port 258 nsew signal input
rlabel metal2 s 137558 159200 137614 160000 6 irq_id_i[3]
port 259 nsew signal input
rlabel metal2 s 106278 159200 106334 160000 6 irq_id_i[4]
port 260 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 irq_id_o[0]
port 261 nsew signal output
rlabel metal3 s 239200 93848 240000 93968 6 irq_id_o[1]
port 262 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 irq_id_o[2]
port 263 nsew signal output
rlabel metal3 s 239200 63248 240000 63368 6 irq_id_o[3]
port 264 nsew signal output
rlabel metal2 s 184478 159200 184534 160000 6 irq_id_o[4]
port 265 nsew signal output
rlabel metal2 s 78678 0 78734 800 6 reset
port 266 nsew signal input
rlabel metal4 s 234208 2128 234528 157808 6 VPWR
port 267 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 157808 6 VPWR
port 268 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 157808 6 VPWR
port 269 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 157808 6 VPWR
port 270 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 157808 6 VPWR
port 271 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 157808 6 VPWR
port 272 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 157808 6 VPWR
port 273 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 157808 6 VPWR
port 274 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 157808 6 VPWR
port 275 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 157808 6 VPWR
port 276 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 157808 6 VPWR
port 277 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 157808 6 VPWR
port 278 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 157808 6 VPWR
port 279 nsew power bidirectional
rlabel metal4 s 104208 95452 104528 157808 6 VPWR
port 280 nsew power bidirectional
rlabel metal4 s 94208 95452 94528 157808 6 VPWR
port 281 nsew power bidirectional
rlabel metal4 s 84208 95452 84528 157808 6 VPWR
port 282 nsew power bidirectional
rlabel metal4 s 74208 95452 74528 157808 6 VPWR
port 283 nsew power bidirectional
rlabel metal4 s 64208 95452 64528 157808 6 VPWR
port 284 nsew power bidirectional
rlabel metal4 s 54208 95452 54528 157808 6 VPWR
port 285 nsew power bidirectional
rlabel metal4 s 44208 95452 44528 157808 6 VPWR
port 286 nsew power bidirectional
rlabel metal4 s 34208 95452 34528 157808 6 VPWR
port 287 nsew power bidirectional
rlabel metal4 s 24208 95452 24528 157808 6 VPWR
port 288 nsew power bidirectional
rlabel metal4 s 14208 95452 14528 157808 6 VPWR
port 289 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 157808 6 VPWR
port 290 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 14048 6 VPWR
port 291 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 14048 6 VPWR
port 292 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 14048 6 VPWR
port 293 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 14048 6 VPWR
port 294 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 14048 6 VPWR
port 295 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 14048 6 VPWR
port 296 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 14048 6 VPWR
port 297 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 14048 6 VPWR
port 298 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 14048 6 VPWR
port 299 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 14048 6 VPWR
port 300 nsew power bidirectional
rlabel metal5 s 1104 127842 238832 128162 6 VPWR
port 301 nsew power bidirectional
rlabel metal5 s 1104 97206 238832 97526 6 VPWR
port 302 nsew power bidirectional
rlabel metal5 s 1104 66570 238832 66890 6 VPWR
port 303 nsew power bidirectional
rlabel metal5 s 1104 35934 238832 36254 6 VPWR
port 304 nsew power bidirectional
rlabel metal5 s 1104 5298 238832 5618 6 VPWR
port 305 nsew power bidirectional
rlabel metal4 s 229208 2128 229528 157808 6 VGND
port 306 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 157808 6 VGND
port 307 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 157808 6 VGND
port 308 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 157808 6 VGND
port 309 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 157808 6 VGND
port 310 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 157808 6 VGND
port 311 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 157808 6 VGND
port 312 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 157808 6 VGND
port 313 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 157808 6 VGND
port 314 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 157808 6 VGND
port 315 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 157808 6 VGND
port 316 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 157808 6 VGND
port 317 nsew ground bidirectional
rlabel metal4 s 109208 95452 109528 157808 6 VGND
port 318 nsew ground bidirectional
rlabel metal4 s 99208 95452 99528 157808 6 VGND
port 319 nsew ground bidirectional
rlabel metal4 s 89208 95452 89528 157808 6 VGND
port 320 nsew ground bidirectional
rlabel metal4 s 79208 95452 79528 157808 6 VGND
port 321 nsew ground bidirectional
rlabel metal4 s 69208 95452 69528 157808 6 VGND
port 322 nsew ground bidirectional
rlabel metal4 s 59208 95452 59528 157808 6 VGND
port 323 nsew ground bidirectional
rlabel metal4 s 49208 95452 49528 157808 6 VGND
port 324 nsew ground bidirectional
rlabel metal4 s 39208 95452 39528 157808 6 VGND
port 325 nsew ground bidirectional
rlabel metal4 s 29208 95452 29528 157808 6 VGND
port 326 nsew ground bidirectional
rlabel metal4 s 19208 95452 19528 157808 6 VGND
port 327 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 157808 6 VGND
port 328 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 14048 6 VGND
port 329 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 14048 6 VGND
port 330 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 14048 6 VGND
port 331 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 14048 6 VGND
port 332 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 14048 6 VGND
port 333 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 14048 6 VGND
port 334 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 14048 6 VGND
port 335 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 14048 6 VGND
port 336 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 14048 6 VGND
port 337 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 14048 6 VGND
port 338 nsew ground bidirectional
rlabel metal5 s 1104 143160 238832 143480 6 VGND
port 339 nsew ground bidirectional
rlabel metal5 s 1104 112524 238832 112844 6 VGND
port 340 nsew ground bidirectional
rlabel metal5 s 1104 81888 238832 82208 6 VGND
port 341 nsew ground bidirectional
rlabel metal5 s 1104 51252 238832 51572 6 VGND
port 342 nsew ground bidirectional
rlabel metal5 s 1104 20616 238832 20936 6 VGND
port 343 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 240000 160000
string LEFview TRUE
string GDS_FILE /project/openlane/core_sram/runs/core_sram/results/magic/core_sram.gds
string GDS_END 67478202
string GDS_START 10607422
<< end >>

