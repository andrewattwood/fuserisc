magic
tech sky130A
magscale 1 2
timestamp 1624390264
<< obsli1 >>
rect 1104 1717 58880 27761
<< obsm1 >>
rect 474 1504 59418 28144
<< metal2 >>
rect 938 29200 994 30000
rect 1398 29200 1454 30000
rect 2318 29200 2374 30000
rect 2778 29200 2834 30000
rect 3238 29200 3294 30000
rect 4158 29200 4214 30000
rect 4618 29200 4674 30000
rect 5538 29200 5594 30000
rect 5998 29200 6054 30000
rect 6458 29200 6514 30000
rect 7378 29200 7434 30000
rect 7838 29200 7894 30000
rect 8758 29200 8814 30000
rect 9218 29200 9274 30000
rect 9678 29200 9734 30000
rect 10598 29200 10654 30000
rect 11058 29200 11114 30000
rect 11978 29200 12034 30000
rect 12438 29200 12494 30000
rect 12898 29200 12954 30000
rect 13818 29200 13874 30000
rect 14278 29200 14334 30000
rect 14738 29200 14794 30000
rect 15658 29200 15714 30000
rect 16118 29200 16174 30000
rect 17038 29200 17094 30000
rect 17498 29200 17554 30000
rect 17958 29200 18014 30000
rect 18878 29200 18934 30000
rect 19338 29200 19394 30000
rect 20258 29200 20314 30000
rect 20718 29200 20774 30000
rect 21178 29200 21234 30000
rect 22098 29200 22154 30000
rect 22558 29200 22614 30000
rect 23478 29200 23534 30000
rect 23938 29200 23994 30000
rect 24398 29200 24454 30000
rect 25318 29200 25374 30000
rect 25778 29200 25834 30000
rect 26698 29200 26754 30000
rect 27158 29200 27214 30000
rect 27618 29200 27674 30000
rect 28538 29200 28594 30000
rect 28998 29200 29054 30000
rect 29918 29200 29974 30000
rect 30378 29200 30434 30000
rect 30838 29200 30894 30000
rect 31758 29200 31814 30000
rect 32218 29200 32274 30000
rect 33138 29200 33194 30000
rect 33598 29200 33654 30000
rect 34058 29200 34114 30000
rect 34978 29200 35034 30000
rect 35438 29200 35494 30000
rect 36358 29200 36414 30000
rect 36818 29200 36874 30000
rect 37278 29200 37334 30000
rect 38198 29200 38254 30000
rect 38658 29200 38714 30000
rect 39578 29200 39634 30000
rect 40038 29200 40094 30000
rect 40498 29200 40554 30000
rect 41418 29200 41474 30000
rect 41878 29200 41934 30000
rect 42798 29200 42854 30000
rect 43258 29200 43314 30000
rect 43718 29200 43774 30000
rect 44638 29200 44694 30000
rect 45098 29200 45154 30000
rect 45558 29200 45614 30000
rect 46478 29200 46534 30000
rect 46938 29200 46994 30000
rect 47858 29200 47914 30000
rect 48318 29200 48374 30000
rect 48778 29200 48834 30000
rect 49698 29200 49754 30000
rect 50158 29200 50214 30000
rect 51078 29200 51134 30000
rect 51538 29200 51594 30000
rect 51998 29200 52054 30000
rect 52918 29200 52974 30000
rect 53378 29200 53434 30000
rect 54298 29200 54354 30000
rect 54758 29200 54814 30000
rect 55218 29200 55274 30000
rect 56138 29200 56194 30000
rect 56598 29200 56654 30000
rect 57518 29200 57574 30000
rect 57978 29200 58034 30000
rect 58438 29200 58494 30000
rect 59358 29200 59414 30000
rect 478 0 534 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57518 0 57574 800
rect 57978 0 58034 800
rect 58898 0 58954 800
rect 59358 0 59414 800
<< obsm2 >>
rect 480 29144 882 29200
rect 1050 29144 1342 29200
rect 1510 29144 2262 29200
rect 2430 29144 2722 29200
rect 2890 29144 3182 29200
rect 3350 29144 4102 29200
rect 4270 29144 4562 29200
rect 4730 29144 5482 29200
rect 5650 29144 5942 29200
rect 6110 29144 6402 29200
rect 6570 29144 7322 29200
rect 7490 29144 7782 29200
rect 7950 29144 8702 29200
rect 8870 29144 9162 29200
rect 9330 29144 9622 29200
rect 9790 29144 10542 29200
rect 10710 29144 11002 29200
rect 11170 29144 11922 29200
rect 12090 29144 12382 29200
rect 12550 29144 12842 29200
rect 13010 29144 13762 29200
rect 13930 29144 14222 29200
rect 14390 29144 14682 29200
rect 14850 29144 15602 29200
rect 15770 29144 16062 29200
rect 16230 29144 16982 29200
rect 17150 29144 17442 29200
rect 17610 29144 17902 29200
rect 18070 29144 18822 29200
rect 18990 29144 19282 29200
rect 19450 29144 20202 29200
rect 20370 29144 20662 29200
rect 20830 29144 21122 29200
rect 21290 29144 22042 29200
rect 22210 29144 22502 29200
rect 22670 29144 23422 29200
rect 23590 29144 23882 29200
rect 24050 29144 24342 29200
rect 24510 29144 25262 29200
rect 25430 29144 25722 29200
rect 25890 29144 26642 29200
rect 26810 29144 27102 29200
rect 27270 29144 27562 29200
rect 27730 29144 28482 29200
rect 28650 29144 28942 29200
rect 29110 29144 29862 29200
rect 30030 29144 30322 29200
rect 30490 29144 30782 29200
rect 30950 29144 31702 29200
rect 31870 29144 32162 29200
rect 32330 29144 33082 29200
rect 33250 29144 33542 29200
rect 33710 29144 34002 29200
rect 34170 29144 34922 29200
rect 35090 29144 35382 29200
rect 35550 29144 36302 29200
rect 36470 29144 36762 29200
rect 36930 29144 37222 29200
rect 37390 29144 38142 29200
rect 38310 29144 38602 29200
rect 38770 29144 39522 29200
rect 39690 29144 39982 29200
rect 40150 29144 40442 29200
rect 40610 29144 41362 29200
rect 41530 29144 41822 29200
rect 41990 29144 42742 29200
rect 42910 29144 43202 29200
rect 43370 29144 43662 29200
rect 43830 29144 44582 29200
rect 44750 29144 45042 29200
rect 45210 29144 45502 29200
rect 45670 29144 46422 29200
rect 46590 29144 46882 29200
rect 47050 29144 47802 29200
rect 47970 29144 48262 29200
rect 48430 29144 48722 29200
rect 48890 29144 49642 29200
rect 49810 29144 50102 29200
rect 50270 29144 51022 29200
rect 51190 29144 51482 29200
rect 51650 29144 51942 29200
rect 52110 29144 52862 29200
rect 53030 29144 53322 29200
rect 53490 29144 54242 29200
rect 54410 29144 54702 29200
rect 54870 29144 55162 29200
rect 55330 29144 56082 29200
rect 56250 29144 56542 29200
rect 56710 29144 57462 29200
rect 57630 29144 57922 29200
rect 58090 29144 58382 29200
rect 58550 29144 59302 29200
rect 480 856 59412 29144
rect 590 711 882 856
rect 1050 711 1342 856
rect 1510 711 2262 856
rect 2430 711 2722 856
rect 2890 711 3182 856
rect 3350 711 4102 856
rect 4270 711 4562 856
rect 4730 711 5482 856
rect 5650 711 5942 856
rect 6110 711 6402 856
rect 6570 711 7322 856
rect 7490 711 7782 856
rect 7950 711 8702 856
rect 8870 711 9162 856
rect 9330 711 9622 856
rect 9790 711 10542 856
rect 10710 711 11002 856
rect 11170 711 11922 856
rect 12090 711 12382 856
rect 12550 711 12842 856
rect 13010 711 13762 856
rect 13930 711 14222 856
rect 14390 711 15142 856
rect 15310 711 15602 856
rect 15770 711 16062 856
rect 16230 711 16982 856
rect 17150 711 17442 856
rect 17610 711 18362 856
rect 18530 711 18822 856
rect 18990 711 19282 856
rect 19450 711 20202 856
rect 20370 711 20662 856
rect 20830 711 21582 856
rect 21750 711 22042 856
rect 22210 711 22502 856
rect 22670 711 23422 856
rect 23590 711 23882 856
rect 24050 711 24802 856
rect 24970 711 25262 856
rect 25430 711 25722 856
rect 25890 711 26642 856
rect 26810 711 27102 856
rect 27270 711 28022 856
rect 28190 711 28482 856
rect 28650 711 28942 856
rect 29110 711 29862 856
rect 30030 711 30322 856
rect 30490 711 31242 856
rect 31410 711 31702 856
rect 31870 711 32162 856
rect 32330 711 33082 856
rect 33250 711 33542 856
rect 33710 711 34002 856
rect 34170 711 34922 856
rect 35090 711 35382 856
rect 35550 711 36302 856
rect 36470 711 36762 856
rect 36930 711 37222 856
rect 37390 711 38142 856
rect 38310 711 38602 856
rect 38770 711 39522 856
rect 39690 711 39982 856
rect 40150 711 40442 856
rect 40610 711 41362 856
rect 41530 711 41822 856
rect 41990 711 42742 856
rect 42910 711 43202 856
rect 43370 711 43662 856
rect 43830 711 44582 856
rect 44750 711 45042 856
rect 45210 711 45962 856
rect 46130 711 46422 856
rect 46590 711 46882 856
rect 47050 711 47802 856
rect 47970 711 48262 856
rect 48430 711 49182 856
rect 49350 711 49642 856
rect 49810 711 50102 856
rect 50270 711 51022 856
rect 51190 711 51482 856
rect 51650 711 52402 856
rect 52570 711 52862 856
rect 53030 711 53322 856
rect 53490 711 54242 856
rect 54410 711 54702 856
rect 54870 711 55622 856
rect 55790 711 56082 856
rect 56250 711 56542 856
rect 56710 711 57462 856
rect 57630 711 57922 856
rect 58090 711 58842 856
rect 59010 711 59302 856
<< metal3 >>
rect 0 28568 800 28688
rect 59200 28568 60000 28688
rect 0 27888 800 28008
rect 0 27208 800 27328
rect 59200 27208 60000 27328
rect 59200 26528 60000 26648
rect 0 25848 800 25968
rect 59200 25848 60000 25968
rect 0 25168 800 25288
rect 59200 24488 60000 24608
rect 0 23808 800 23928
rect 59200 23808 60000 23928
rect 0 23128 800 23248
rect 0 22448 800 22568
rect 59200 22448 60000 22568
rect 59200 21768 60000 21888
rect 0 21088 800 21208
rect 59200 21088 60000 21208
rect 0 20408 800 20528
rect 59200 19728 60000 19848
rect 0 19048 800 19168
rect 59200 19048 60000 19168
rect 0 18368 800 18488
rect 0 17688 800 17808
rect 59200 17688 60000 17808
rect 59200 17008 60000 17128
rect 0 16328 800 16448
rect 59200 16328 60000 16448
rect 0 15648 800 15768
rect 59200 14968 60000 15088
rect 0 14288 800 14408
rect 59200 14288 60000 14408
rect 0 13608 800 13728
rect 0 12928 800 13048
rect 59200 12928 60000 13048
rect 59200 12248 60000 12368
rect 0 11568 800 11688
rect 59200 11568 60000 11688
rect 0 10888 800 11008
rect 59200 10208 60000 10328
rect 0 9528 800 9648
rect 59200 9528 60000 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
rect 59200 8168 60000 8288
rect 59200 7488 60000 7608
rect 0 6808 800 6928
rect 59200 6808 60000 6928
rect 0 6128 800 6248
rect 59200 5448 60000 5568
rect 0 4768 800 4888
rect 59200 4768 60000 4888
rect 0 4088 800 4208
rect 59200 4088 60000 4208
rect 0 3408 800 3528
rect 59200 2728 60000 2848
rect 0 2048 800 2168
rect 59200 2048 60000 2168
rect 0 1368 800 1488
rect 59200 688 60000 808
<< obsm3 >>
rect 880 28488 59120 28661
rect 800 28088 59200 28488
rect 880 27808 59200 28088
rect 800 27408 59200 27808
rect 880 27128 59120 27408
rect 800 26728 59200 27128
rect 800 26448 59120 26728
rect 800 26048 59200 26448
rect 880 25768 59120 26048
rect 800 25368 59200 25768
rect 880 25088 59200 25368
rect 800 24688 59200 25088
rect 800 24408 59120 24688
rect 800 24008 59200 24408
rect 880 23728 59120 24008
rect 800 23328 59200 23728
rect 880 23048 59200 23328
rect 800 22648 59200 23048
rect 880 22368 59120 22648
rect 800 21968 59200 22368
rect 800 21688 59120 21968
rect 800 21288 59200 21688
rect 880 21008 59120 21288
rect 800 20608 59200 21008
rect 880 20328 59200 20608
rect 800 19928 59200 20328
rect 800 19648 59120 19928
rect 800 19248 59200 19648
rect 880 18968 59120 19248
rect 800 18568 59200 18968
rect 880 18288 59200 18568
rect 800 17888 59200 18288
rect 880 17608 59120 17888
rect 800 17208 59200 17608
rect 800 16928 59120 17208
rect 800 16528 59200 16928
rect 880 16248 59120 16528
rect 800 15848 59200 16248
rect 880 15568 59200 15848
rect 800 15168 59200 15568
rect 800 14888 59120 15168
rect 800 14488 59200 14888
rect 880 14208 59120 14488
rect 800 13808 59200 14208
rect 880 13528 59200 13808
rect 800 13128 59200 13528
rect 880 12848 59120 13128
rect 800 12448 59200 12848
rect 800 12168 59120 12448
rect 800 11768 59200 12168
rect 880 11488 59120 11768
rect 800 11088 59200 11488
rect 880 10808 59200 11088
rect 800 10408 59200 10808
rect 800 10128 59120 10408
rect 800 9728 59200 10128
rect 880 9448 59120 9728
rect 800 9048 59200 9448
rect 880 8768 59200 9048
rect 800 8368 59200 8768
rect 880 8088 59120 8368
rect 800 7688 59200 8088
rect 800 7408 59120 7688
rect 800 7008 59200 7408
rect 880 6728 59120 7008
rect 800 6328 59200 6728
rect 880 6048 59200 6328
rect 800 5648 59200 6048
rect 800 5368 59120 5648
rect 800 4968 59200 5368
rect 880 4688 59120 4968
rect 800 4288 59200 4688
rect 880 4008 59120 4288
rect 800 3608 59200 4008
rect 880 3328 59200 3608
rect 800 2928 59200 3328
rect 800 2648 59120 2928
rect 800 2248 59200 2648
rect 880 1968 59120 2248
rect 800 1568 59200 1968
rect 880 1288 59200 1568
rect 800 888 59200 1288
rect 800 715 59120 888
<< metal4 >>
rect 10576 2128 10896 27792
rect 20208 2128 20528 27792
rect 29840 2128 30160 27792
rect 39472 2128 39792 27792
rect 49104 2128 49424 27792
<< metal5 >>
rect 1104 23341 58880 23661
rect 1104 19067 58880 19387
rect 1104 14792 58880 15112
rect 1104 10517 58880 10837
rect 1104 6243 58880 6563
<< obsm5 >>
rect 1104 15432 58880 18747
rect 1104 11157 58880 14472
rect 1104 6883 58880 10197
<< labels >>
rlabel metal3 s 0 23808 800 23928 6 core_a_data_addr_o[0]
port 1 nsew signal output
rlabel metal2 s 54298 29200 54354 30000 6 core_a_data_addr_o[1]
port 2 nsew signal output
rlabel metal2 s 43718 29200 43774 30000 6 core_a_data_addr_o[2]
port 3 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 core_a_data_addr_o[3]
port 4 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 core_a_data_addr_o[4]
port 5 nsew signal output
rlabel metal2 s 29918 29200 29974 30000 6 core_a_data_addr_o[5]
port 6 nsew signal output
rlabel metal2 s 10598 29200 10654 30000 6 core_a_data_addr_o[6]
port 7 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 core_a_data_addr_o[7]
port 8 nsew signal output
rlabel metal2 s 55218 29200 55274 30000 6 core_a_data_addr_o[8]
port 9 nsew signal output
rlabel metal3 s 59200 9528 60000 9648 6 core_a_data_addr_o[9]
port 10 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 core_a_data_be_o[0]
port 11 nsew signal output
rlabel metal2 s 23938 29200 23994 30000 6 core_a_data_be_o[1]
port 12 nsew signal output
rlabel metal2 s 13818 29200 13874 30000 6 core_a_data_be_o[2]
port 13 nsew signal output
rlabel metal3 s 59200 19048 60000 19168 6 core_a_data_be_o[3]
port 14 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 core_a_data_rdata_i[0]
port 15 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 core_a_data_rdata_i[10]
port 16 nsew signal input
rlabel metal3 s 59200 22448 60000 22568 6 core_a_data_rdata_i[11]
port 17 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 core_a_data_rdata_i[12]
port 18 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 core_a_data_rdata_i[13]
port 19 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 core_a_data_rdata_i[14]
port 20 nsew signal input
rlabel metal2 s 51998 29200 52054 30000 6 core_a_data_rdata_i[15]
port 21 nsew signal input
rlabel metal2 s 57978 29200 58034 30000 6 core_a_data_rdata_i[16]
port 22 nsew signal input
rlabel metal3 s 59200 2728 60000 2848 6 core_a_data_rdata_i[17]
port 23 nsew signal input
rlabel metal3 s 59200 26528 60000 26648 6 core_a_data_rdata_i[18]
port 24 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 core_a_data_rdata_i[19]
port 25 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 core_a_data_rdata_i[1]
port 26 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 core_a_data_rdata_i[20]
port 27 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 core_a_data_rdata_i[21]
port 28 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 core_a_data_rdata_i[22]
port 29 nsew signal input
rlabel metal2 s 28538 29200 28594 30000 6 core_a_data_rdata_i[23]
port 30 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 core_a_data_rdata_i[24]
port 31 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 core_a_data_rdata_i[25]
port 32 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 core_a_data_rdata_i[26]
port 33 nsew signal input
rlabel metal2 s 31758 29200 31814 30000 6 core_a_data_rdata_i[27]
port 34 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 core_a_data_rdata_i[28]
port 35 nsew signal input
rlabel metal2 s 41418 29200 41474 30000 6 core_a_data_rdata_i[29]
port 36 nsew signal input
rlabel metal2 s 11978 29200 12034 30000 6 core_a_data_rdata_i[2]
port 37 nsew signal input
rlabel metal2 s 38658 29200 38714 30000 6 core_a_data_rdata_i[30]
port 38 nsew signal input
rlabel metal2 s 26698 29200 26754 30000 6 core_a_data_rdata_i[31]
port 39 nsew signal input
rlabel metal2 s 15658 29200 15714 30000 6 core_a_data_rdata_i[3]
port 40 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 core_a_data_rdata_i[4]
port 41 nsew signal input
rlabel metal3 s 59200 14288 60000 14408 6 core_a_data_rdata_i[5]
port 42 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 core_a_data_rdata_i[6]
port 43 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 core_a_data_rdata_i[7]
port 44 nsew signal input
rlabel metal2 s 45098 29200 45154 30000 6 core_a_data_rdata_i[8]
port 45 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 core_a_data_rdata_i[9]
port 46 nsew signal input
rlabel metal2 s 24398 29200 24454 30000 6 core_a_data_req_o
port 47 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 core_a_data_rvalid_i
port 48 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 core_a_data_wdata_o[0]
port 49 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 core_a_data_wdata_o[10]
port 50 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 core_a_data_wdata_o[11]
port 51 nsew signal output
rlabel metal2 s 35438 29200 35494 30000 6 core_a_data_wdata_o[12]
port 52 nsew signal output
rlabel metal2 s 9678 29200 9734 30000 6 core_a_data_wdata_o[13]
port 53 nsew signal output
rlabel metal2 s 12438 29200 12494 30000 6 core_a_data_wdata_o[14]
port 54 nsew signal output
rlabel metal2 s 43258 29200 43314 30000 6 core_a_data_wdata_o[15]
port 55 nsew signal output
rlabel metal2 s 46478 29200 46534 30000 6 core_a_data_wdata_o[16]
port 56 nsew signal output
rlabel metal3 s 59200 16328 60000 16448 6 core_a_data_wdata_o[17]
port 57 nsew signal output
rlabel metal2 s 19338 29200 19394 30000 6 core_a_data_wdata_o[18]
port 58 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 core_a_data_wdata_o[19]
port 59 nsew signal output
rlabel metal2 s 54758 29200 54814 30000 6 core_a_data_wdata_o[1]
port 60 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 core_a_data_wdata_o[20]
port 61 nsew signal output
rlabel metal2 s 57518 29200 57574 30000 6 core_a_data_wdata_o[21]
port 62 nsew signal output
rlabel metal2 s 3238 29200 3294 30000 6 core_a_data_wdata_o[22]
port 63 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 core_a_data_wdata_o[23]
port 64 nsew signal output
rlabel metal3 s 59200 10208 60000 10328 6 core_a_data_wdata_o[24]
port 65 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 core_a_data_wdata_o[25]
port 66 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 core_a_data_wdata_o[26]
port 67 nsew signal output
rlabel metal3 s 59200 19728 60000 19848 6 core_a_data_wdata_o[27]
port 68 nsew signal output
rlabel metal2 s 25778 29200 25834 30000 6 core_a_data_wdata_o[28]
port 69 nsew signal output
rlabel metal2 s 37278 29200 37334 30000 6 core_a_data_wdata_o[29]
port 70 nsew signal output
rlabel metal2 s 4158 0 4214 800 6 core_a_data_wdata_o[2]
port 71 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 core_a_data_wdata_o[30]
port 72 nsew signal output
rlabel metal2 s 45558 29200 45614 30000 6 core_a_data_wdata_o[31]
port 73 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 core_a_data_wdata_o[3]
port 74 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 core_a_data_wdata_o[4]
port 75 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 core_a_data_wdata_o[5]
port 76 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 core_a_data_wdata_o[6]
port 77 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 core_a_data_wdata_o[7]
port 78 nsew signal output
rlabel metal2 s 48778 29200 48834 30000 6 core_a_data_wdata_o[8]
port 79 nsew signal output
rlabel metal2 s 17958 29200 18014 30000 6 core_a_data_wdata_o[9]
port 80 nsew signal output
rlabel metal3 s 59200 8168 60000 8288 6 core_a_data_we_o
port 81 nsew signal output
rlabel metal2 s 2318 0 2374 800 6 core_b_data_addr_o[0]
port 82 nsew signal output
rlabel metal2 s 32218 29200 32274 30000 6 core_b_data_addr_o[1]
port 83 nsew signal output
rlabel metal2 s 2778 29200 2834 30000 6 core_b_data_addr_o[2]
port 84 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 core_b_data_addr_o[3]
port 85 nsew signal output
rlabel metal2 s 56138 29200 56194 30000 6 core_b_data_addr_o[4]
port 86 nsew signal output
rlabel metal2 s 36818 29200 36874 30000 6 core_b_data_addr_o[5]
port 87 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 core_b_data_addr_o[6]
port 88 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 core_b_data_addr_o[7]
port 89 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 core_b_data_addr_o[8]
port 90 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 core_b_data_addr_o[9]
port 91 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 core_b_data_be_o[0]
port 92 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 core_b_data_be_o[1]
port 93 nsew signal output
rlabel metal2 s 5538 29200 5594 30000 6 core_b_data_be_o[2]
port 94 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 core_b_data_be_o[3]
port 95 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 core_b_data_rdata_i[0]
port 96 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 core_b_data_rdata_i[10]
port 97 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 core_b_data_rdata_i[11]
port 98 nsew signal input
rlabel metal2 s 17038 29200 17094 30000 6 core_b_data_rdata_i[12]
port 99 nsew signal input
rlabel metal2 s 53378 29200 53434 30000 6 core_b_data_rdata_i[13]
port 100 nsew signal input
rlabel metal2 s 33598 29200 33654 30000 6 core_b_data_rdata_i[14]
port 101 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 core_b_data_rdata_i[15]
port 102 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 core_b_data_rdata_i[16]
port 103 nsew signal input
rlabel metal3 s 59200 25848 60000 25968 6 core_b_data_rdata_i[17]
port 104 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 core_b_data_rdata_i[18]
port 105 nsew signal input
rlabel metal2 s 40038 29200 40094 30000 6 core_b_data_rdata_i[19]
port 106 nsew signal input
rlabel metal2 s 938 29200 994 30000 6 core_b_data_rdata_i[1]
port 107 nsew signal input
rlabel metal3 s 59200 2048 60000 2168 6 core_b_data_rdata_i[20]
port 108 nsew signal input
rlabel metal3 s 59200 4088 60000 4208 6 core_b_data_rdata_i[21]
port 109 nsew signal input
rlabel metal2 s 36358 29200 36414 30000 6 core_b_data_rdata_i[22]
port 110 nsew signal input
rlabel metal3 s 59200 17688 60000 17808 6 core_b_data_rdata_i[23]
port 111 nsew signal input
rlabel metal2 s 12898 29200 12954 30000 6 core_b_data_rdata_i[24]
port 112 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 core_b_data_rdata_i[25]
port 113 nsew signal input
rlabel metal2 s 46938 29200 46994 30000 6 core_b_data_rdata_i[26]
port 114 nsew signal input
rlabel metal2 s 4618 29200 4674 30000 6 core_b_data_rdata_i[27]
port 115 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 core_b_data_rdata_i[28]
port 116 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 core_b_data_rdata_i[29]
port 117 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 core_b_data_rdata_i[2]
port 118 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 core_b_data_rdata_i[30]
port 119 nsew signal input
rlabel metal2 s 11058 29200 11114 30000 6 core_b_data_rdata_i[31]
port 120 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 core_b_data_rdata_i[3]
port 121 nsew signal input
rlabel metal2 s 48318 29200 48374 30000 6 core_b_data_rdata_i[4]
port 122 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 core_b_data_rdata_i[5]
port 123 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 core_b_data_rdata_i[6]
port 124 nsew signal input
rlabel metal3 s 59200 4768 60000 4888 6 core_b_data_rdata_i[7]
port 125 nsew signal input
rlabel metal2 s 34058 29200 34114 30000 6 core_b_data_rdata_i[8]
port 126 nsew signal input
rlabel metal3 s 59200 21088 60000 21208 6 core_b_data_rdata_i[9]
port 127 nsew signal input
rlabel metal2 s 52918 29200 52974 30000 6 core_b_data_req_o
port 128 nsew signal output
rlabel metal2 s 51538 29200 51594 30000 6 core_b_data_rvalid_i
port 129 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 core_b_data_wdata_o[0]
port 130 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 core_b_data_wdata_o[10]
port 131 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 core_b_data_wdata_o[11]
port 132 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 core_b_data_wdata_o[12]
port 133 nsew signal output
rlabel metal2 s 50158 29200 50214 30000 6 core_b_data_wdata_o[13]
port 134 nsew signal output
rlabel metal2 s 41878 0 41934 800 6 core_b_data_wdata_o[14]
port 135 nsew signal output
rlabel metal2 s 39578 0 39634 800 6 core_b_data_wdata_o[15]
port 136 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 core_b_data_wdata_o[16]
port 137 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 core_b_data_wdata_o[17]
port 138 nsew signal output
rlabel metal2 s 20718 29200 20774 30000 6 core_b_data_wdata_o[18]
port 139 nsew signal output
rlabel metal2 s 30838 29200 30894 30000 6 core_b_data_wdata_o[19]
port 140 nsew signal output
rlabel metal2 s 5998 29200 6054 30000 6 core_b_data_wdata_o[1]
port 141 nsew signal output
rlabel metal2 s 27618 29200 27674 30000 6 core_b_data_wdata_o[20]
port 142 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 core_b_data_wdata_o[21]
port 143 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 core_b_data_wdata_o[22]
port 144 nsew signal output
rlabel metal2 s 28998 29200 29054 30000 6 core_b_data_wdata_o[23]
port 145 nsew signal output
rlabel metal2 s 22558 29200 22614 30000 6 core_b_data_wdata_o[24]
port 146 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 core_b_data_wdata_o[25]
port 147 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 core_b_data_wdata_o[26]
port 148 nsew signal output
rlabel metal3 s 59200 21768 60000 21888 6 core_b_data_wdata_o[27]
port 149 nsew signal output
rlabel metal3 s 59200 28568 60000 28688 6 core_b_data_wdata_o[28]
port 150 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 core_b_data_wdata_o[29]
port 151 nsew signal output
rlabel metal2 s 49698 29200 49754 30000 6 core_b_data_wdata_o[2]
port 152 nsew signal output
rlabel metal2 s 42798 29200 42854 30000 6 core_b_data_wdata_o[30]
port 153 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 core_b_data_wdata_o[31]
port 154 nsew signal output
rlabel metal2 s 56598 29200 56654 30000 6 core_b_data_wdata_o[3]
port 155 nsew signal output
rlabel metal2 s 16118 29200 16174 30000 6 core_b_data_wdata_o[4]
port 156 nsew signal output
rlabel metal2 s 51078 0 51134 800 6 core_b_data_wdata_o[5]
port 157 nsew signal output
rlabel metal2 s 44638 29200 44694 30000 6 core_b_data_wdata_o[6]
port 158 nsew signal output
rlabel metal2 s 27158 29200 27214 30000 6 core_b_data_wdata_o[7]
port 159 nsew signal output
rlabel metal2 s 6458 29200 6514 30000 6 core_b_data_wdata_o[8]
port 160 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 core_b_data_wdata_o[9]
port 161 nsew signal output
rlabel metal2 s 51078 29200 51134 30000 6 core_b_data_we_o
port 162 nsew signal output
rlabel metal3 s 59200 12248 60000 12368 6 wb_data_addr_i[0]
port 163 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_data_addr_i[10]
port 164 nsew signal input
rlabel metal2 s 2318 29200 2374 30000 6 wb_data_addr_i[1]
port 165 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wb_data_addr_i[2]
port 166 nsew signal input
rlabel metal3 s 59200 14968 60000 15088 6 wb_data_addr_i[3]
port 167 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wb_data_addr_i[4]
port 168 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wb_data_addr_i[5]
port 169 nsew signal input
rlabel metal2 s 7378 29200 7434 30000 6 wb_data_addr_i[6]
port 170 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wb_data_addr_i[7]
port 171 nsew signal input
rlabel metal2 s 7838 29200 7894 30000 6 wb_data_addr_i[8]
port 172 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wb_data_addr_i[9]
port 173 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wb_data_be_i[0]
port 174 nsew signal input
rlabel metal2 s 8758 29200 8814 30000 6 wb_data_be_i[1]
port 175 nsew signal input
rlabel metal2 s 17498 29200 17554 30000 6 wb_data_be_i[2]
port 176 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wb_data_be_i[3]
port 177 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wb_data_rdata_o[0]
port 178 nsew signal output
rlabel metal2 s 14738 29200 14794 30000 6 wb_data_rdata_o[10]
port 179 nsew signal output
rlabel metal3 s 59200 11568 60000 11688 6 wb_data_rdata_o[11]
port 180 nsew signal output
rlabel metal2 s 58438 29200 58494 30000 6 wb_data_rdata_o[12]
port 181 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 wb_data_rdata_o[13]
port 182 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 wb_data_rdata_o[14]
port 183 nsew signal output
rlabel metal2 s 24858 0 24914 800 6 wb_data_rdata_o[15]
port 184 nsew signal output
rlabel metal2 s 1398 0 1454 800 6 wb_data_rdata_o[16]
port 185 nsew signal output
rlabel metal2 s 39578 29200 39634 30000 6 wb_data_rdata_o[17]
port 186 nsew signal output
rlabel metal2 s 20258 29200 20314 30000 6 wb_data_rdata_o[18]
port 187 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 wb_data_rdata_o[19]
port 188 nsew signal output
rlabel metal3 s 59200 5448 60000 5568 6 wb_data_rdata_o[1]
port 189 nsew signal output
rlabel metal2 s 41878 29200 41934 30000 6 wb_data_rdata_o[20]
port 190 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 wb_data_rdata_o[21]
port 191 nsew signal output
rlabel metal2 s 1398 29200 1454 30000 6 wb_data_rdata_o[22]
port 192 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 wb_data_rdata_o[23]
port 193 nsew signal output
rlabel metal2 s 21178 29200 21234 30000 6 wb_data_rdata_o[24]
port 194 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 wb_data_rdata_o[25]
port 195 nsew signal output
rlabel metal2 s 9218 29200 9274 30000 6 wb_data_rdata_o[26]
port 196 nsew signal output
rlabel metal2 s 478 0 534 800 6 wb_data_rdata_o[27]
port 197 nsew signal output
rlabel metal2 s 4158 29200 4214 30000 6 wb_data_rdata_o[28]
port 198 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 wb_data_rdata_o[29]
port 199 nsew signal output
rlabel metal2 s 33138 29200 33194 30000 6 wb_data_rdata_o[2]
port 200 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 wb_data_rdata_o[30]
port 201 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wb_data_rdata_o[31]
port 202 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 wb_data_rdata_o[3]
port 203 nsew signal output
rlabel metal2 s 4618 0 4674 800 6 wb_data_rdata_o[4]
port 204 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 wb_data_rdata_o[5]
port 205 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 wb_data_rdata_o[6]
port 206 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wb_data_rdata_o[7]
port 207 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 wb_data_rdata_o[8]
port 208 nsew signal output
rlabel metal2 s 47858 29200 47914 30000 6 wb_data_rdata_o[9]
port 209 nsew signal output
rlabel metal2 s 44638 0 44694 800 6 wb_data_rvalid_o
port 210 nsew signal output
rlabel metal3 s 59200 17008 60000 17128 6 wb_data_wdata_i[0]
port 211 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wb_data_wdata_i[10]
port 212 nsew signal input
rlabel metal3 s 59200 7488 60000 7608 6 wb_data_wdata_i[11]
port 213 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wb_data_wdata_i[12]
port 214 nsew signal input
rlabel metal2 s 14278 29200 14334 30000 6 wb_data_wdata_i[13]
port 215 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wb_data_wdata_i[14]
port 216 nsew signal input
rlabel metal3 s 59200 688 60000 808 6 wb_data_wdata_i[15]
port 217 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wb_data_wdata_i[16]
port 218 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 wb_data_wdata_i[17]
port 219 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_data_wdata_i[18]
port 220 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wb_data_wdata_i[19]
port 221 nsew signal input
rlabel metal3 s 59200 23808 60000 23928 6 wb_data_wdata_i[1]
port 222 nsew signal input
rlabel metal2 s 25318 29200 25374 30000 6 wb_data_wdata_i[20]
port 223 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wb_data_wdata_i[21]
port 224 nsew signal input
rlabel metal2 s 23478 29200 23534 30000 6 wb_data_wdata_i[22]
port 225 nsew signal input
rlabel metal2 s 34978 29200 35034 30000 6 wb_data_wdata_i[23]
port 226 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wb_data_wdata_i[24]
port 227 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wb_data_wdata_i[25]
port 228 nsew signal input
rlabel metal2 s 40498 29200 40554 30000 6 wb_data_wdata_i[26]
port 229 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wb_data_wdata_i[27]
port 230 nsew signal input
rlabel metal3 s 59200 12928 60000 13048 6 wb_data_wdata_i[28]
port 231 nsew signal input
rlabel metal2 s 22098 29200 22154 30000 6 wb_data_wdata_i[29]
port 232 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wb_data_wdata_i[2]
port 233 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wb_data_wdata_i[30]
port 234 nsew signal input
rlabel metal3 s 59200 24488 60000 24608 6 wb_data_wdata_i[31]
port 235 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wb_data_wdata_i[3]
port 236 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wb_data_wdata_i[4]
port 237 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wb_data_wdata_i[5]
port 238 nsew signal input
rlabel metal3 s 59200 6808 60000 6928 6 wb_data_wdata_i[6]
port 239 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wb_data_wdata_i[7]
port 240 nsew signal input
rlabel metal2 s 30378 29200 30434 30000 6 wb_data_wdata_i[8]
port 241 nsew signal input
rlabel metal2 s 38198 29200 38254 30000 6 wb_data_wdata_i[9]
port 242 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 wb_data_we_i
port 243 nsew signal input
rlabel metal2 s 18878 29200 18934 30000 6 wbs_cyc_i
port 244 nsew signal input
rlabel metal2 s 59358 29200 59414 30000 6 wbs_stb_i
port 245 nsew signal input
rlabel metal4 s 49104 2128 49424 27792 6 VPWR
port 246 nsew power bidirectional
rlabel metal4 s 29840 2128 30160 27792 6 VPWR
port 247 nsew power bidirectional
rlabel metal4 s 10576 2128 10896 27792 6 VPWR
port 248 nsew power bidirectional
rlabel metal5 s 1104 23341 58880 23661 6 VPWR
port 249 nsew power bidirectional
rlabel metal5 s 1104 14792 58880 15112 6 VPWR
port 250 nsew power bidirectional
rlabel metal5 s 1104 6243 58880 6563 6 VPWR
port 251 nsew power bidirectional
rlabel metal4 s 39472 2128 39792 27792 6 VGND
port 252 nsew ground bidirectional
rlabel metal4 s 20208 2128 20528 27792 6 VGND
port 253 nsew ground bidirectional
rlabel metal5 s 1104 19067 58880 19387 6 VGND
port 254 nsew ground bidirectional
rlabel metal5 s 1104 10517 58880 10837 6 VGND
port 255 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 60000 30000
string LEFview TRUE
string GDS_FILE /project/openlane/wb_mem_split/runs/wb_mem_split/results/magic/wb_mem_split.gds
string GDS_END 1514626
string GDS_START 128132
<< end >>

