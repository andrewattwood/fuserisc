##
## LEF for PtnCells ;
## created by Innovus v15.20-p005_1 on Sat Jul 17 12:09:20 2021
##

VERSION 5.7 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO eFPGA_CPU_top
  CLASS BLOCK ;
  SIZE 3370.4200 BY 2569.7200 ;
  FOREIGN eFPGA_CPU_top 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.4954 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 243.104 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 10.4123 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 49.4167 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2539.5500 0.8000 2539.8500 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.8654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.744 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 231.256 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1234.3 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2529.1800 0.8000 2529.4800 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.7144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 174.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2518.2000 0.8000 2518.5000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.1164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 192.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2507.2200 0.8000 2507.5200 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 80.1384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 422.896 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2496.2400 0.8000 2496.5400 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.9612 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 254.527 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.048 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 648.7600 0.0000 648.9000 0.4850 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 50.0449 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 247.404 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 505.7000 0.0000 505.8400 0.4850 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.8908 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 174.293 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 2.539 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 15.4908 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 83.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 518.5800 0.0000 518.7200 0.4850 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4754 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 23.864 LAYER met4  ;
    PORT
      LAYER met4 ;
        RECT 648.4500 0.0000 648.7500 0.8000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1004 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2485.2600 0.8000 2485.5600 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.3504 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 145.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2474.8900 0.8000 2475.1900 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.9064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 191.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2463.9100 0.8000 2464.2100 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.8824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 197.168 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.0468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 16.72 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2452.9300 0.8000 2453.2300 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.1604 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.184 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2441.9500 0.8000 2442.2500 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.1964 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.376 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2430.9700 0.8000 2431.2700 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.145 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 246.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2420.6000 0.8000 2420.9000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.6873 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2409.6200 0.8000 2409.9200 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.4904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 167.944 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2398.6400 0.8000 2398.9400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.7164 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 195.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2387.6600 0.8000 2387.9600 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.026 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 230.408 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2376.6800 0.8000 2376.9800 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.0784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 187.08 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2366.3100 0.8000 2366.6100 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.3892 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 179.008 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 29.4468 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 157.52 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2355.3300 0.8000 2355.6300 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.9744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 181.192 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2344.3500 0.8000 2344.6500 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.6178 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 56.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2333.3700 0.8000 2333.6700 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.731 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 282.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2322.3900 0.8000 2322.6900 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.2354 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 172.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.6088 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 30.384 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2312.0200 0.8000 2312.3200 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.6624 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.528 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2301.0400 0.8000 2301.3400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.7684 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 190.76 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2290.0600 0.8000 2290.3600 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.2144 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2279.0800 0.8000 2279.3800 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.4794 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.352 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.3148 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 12.816 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2268.1000 0.8000 2268.4000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.0084 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 176.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2257.7300 0.8000 2258.0300 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.5734 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.72 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2246.7500 0.8000 2247.0500 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 37.6672 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 201.824 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 250.829 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 1338.22 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2235.7700 0.8000 2236.0700 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.4224 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 178.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2224.7900 0.8000 2225.0900 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 35.4784 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 189.68 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.9618 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 21.6 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2213.8100 0.8000 2214.1100 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 40.8072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 218.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2203.4400 0.8000 2203.7400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 47.7552 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 255.16 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2192.4600 0.8000 2192.7600 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.8712 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.672 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2181.4800 0.8000 2181.7800 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 34.5264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 184.136 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2170.5000 0.8000 2170.8000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5018 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.56 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2159.5200 0.8000 2159.8200 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.158 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.672 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2149.1500 0.8000 2149.4500 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2138.1700 0.8000 2138.4700 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2127.1900 0.8000 2127.4900 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2116.2100 0.8000 2116.5100 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2105.2300 0.8000 2105.5300 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2094.8600 0.8000 2095.1600 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2083.8800 0.8000 2084.1800 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2072.9000 0.8000 2073.2000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2061.9200 0.8000 2062.2200 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2050.9400 0.8000 2051.2400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2040.5700 0.8000 2040.8700 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2029.5900 0.8000 2029.8900 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2018.6100 0.8000 2018.9100 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 2007.6300 0.8000 2007.9300 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1996.6500 0.8000 1996.9500 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1986.2800 0.8000 1986.5800 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1975.3000 0.8000 1975.6000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1964.3200 0.8000 1964.6200 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1953.3400 0.8000 1953.6400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1942.3600 0.8000 1942.6600 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1931.9900 0.8000 1932.2900 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1921.0100 0.8000 1921.3100 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.1384 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1910.0300 0.8000 1910.3300 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.8432 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1899.0500 0.8000 1899.3500 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.6904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 94.344 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1888.0700 0.8000 1888.3700 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.2254 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 171.864 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1877.7000 0.8000 1878.0000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.4704 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 98.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1866.7200 0.8000 1867.0200 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.4824 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 82.568 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1855.7400 0.8000 1856.0400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.38 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1844.7600 0.8000 1845.0600 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.482 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 275.4 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1833.7800 0.8000 1834.0800 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.1622 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 225.224 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1823.4100 0.8000 1823.7100 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.0454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 90.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1812.4300 0.8000 1812.7300 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.5064 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 125.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1801.4500 0.8000 1801.7500 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.5326 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 117.502 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 4.6728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 25.392 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 668.0800 0.0000 668.2200 0.4850 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 15.8134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 84.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 5.7918 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 31.36 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1790.4700 0.8000 1790.7700 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.4594 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.912 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.3768 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.48 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1779.4900 0.8000 1779.7900 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.9694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 170.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1769.1200 0.8000 1769.4200 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.2682 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 97.896 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1758.1400 0.8000 1758.4400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.5974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1747.1600 0.8000 1747.4600 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.2104 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.784 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1736.1800 0.8000 1736.4800 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.5152 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 200.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1725.2000 0.8000 1725.5000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.4974 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 130.648 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1714.8300 0.8000 1715.1300 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.0072 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 144.504 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1703.8500 0.8000 1704.1500 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.9454 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 127.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1692.8700 0.8000 1693.1700 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 22.8414 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 121.816 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1681.8900 0.8000 1682.1900 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.3124 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1670.9100 0.8000 1671.2100 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.9154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 175.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1660.5400 0.8000 1660.8400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.1174 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 123.288 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1649.5600 0.8000 1649.8600 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 25.0494 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.592 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1638.5800 0.8000 1638.8800 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.6874 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 89.8848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 479.856 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1627.6000 0.8000 1627.9000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.1579 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 139.952 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 50.9058 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 271.968 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1616.6200 0.8000 1616.9200 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 31.5894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 163.032 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1606.2500 0.8000 1606.5500 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.5142 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 147.208 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1595.2700 0.8000 1595.5700 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.0474 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 112.248 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1584.2900 0.8000 1584.5900 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.6022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.904 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1573.3100 0.8000 1573.6100 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 23.6694 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 126.232 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1562.3300 0.8000 1562.6300 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.3012 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 114.072 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1551.9600 0.8000 1552.2600 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.0154 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 138.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1540.9800 0.8000 1541.2800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 45.2298 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 242.632 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1530.0000 0.8000 1530.3000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.6894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 115.672 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1519.0200 0.8000 1519.3200 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 26.6214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 136.536 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1508.0400 0.8000 1508.3400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 28.1134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 150.4 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 86.6388 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 462.544 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1497.6700 0.8000 1497.9700 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 32.8764 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 169.896 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1486.6900 0.8000 1486.9900 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.8394 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 100.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1475.7100 0.8000 1476.0100 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 29.4016 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 156.8 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.8048 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 42.096 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1464.7300 0.8000 1465.0300 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 24.9564 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 133.096 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1453.7500 0.8000 1454.0500 ;
    END
  END wbs_dat_o[0]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 13.4574 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 71.768 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1443.3800 0.8000 1443.6800 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 16.9894 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 91.552 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 9.0627 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 44.9921 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1432.4000 0.8000 1432.7000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 55.5252 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 296.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1421.4200 0.8000 1421.7200 ;
    END
  END la_data_out[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1410.4400 0.8000 1410.7400 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1399.4600 0.8000 1399.7600 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1389.0900 0.8000 1389.3900 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1378.1100 0.8000 1378.4100 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1367.1300 0.8000 1367.4300 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1356.1500 0.8000 1356.4500 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1345.1700 0.8000 1345.4700 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1334.8000 0.8000 1335.1000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1323.8200 0.8000 1324.1200 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1312.8400 0.8000 1313.1400 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1301.8600 0.8000 1302.1600 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1290.8800 0.8000 1291.1800 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1280.5100 0.8000 1280.8100 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1269.5300 0.8000 1269.8300 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1258.5500 0.8000 1258.8500 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1247.5700 0.8000 1247.8700 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1236.5900 0.8000 1236.8900 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1225.6100 0.8000 1225.9100 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1215.2400 0.8000 1215.5400 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1204.2600 0.8000 1204.5600 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1193.2800 0.8000 1193.5800 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1182.3000 0.8000 1182.6000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1171.3200 0.8000 1171.6200 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1160.9500 0.8000 1161.2500 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1149.9700 0.8000 1150.2700 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1138.9900 0.8000 1139.2900 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1128.0100 0.8000 1128.3100 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1117.0300 0.8000 1117.3300 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1106.6600 0.8000 1106.9600 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1095.6800 0.8000 1095.9800 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1084.7000 0.8000 1085.0000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1073.7200 0.8000 1074.0200 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1062.7400 0.8000 1063.0400 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1052.3700 0.8000 1052.6700 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1041.3900 0.8000 1041.6900 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1030.4100 0.8000 1030.7100 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1019.4300 0.8000 1019.7300 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 1008.4500 0.8000 1008.7500 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 998.0800 0.8000 998.3800 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 987.1000 0.8000 987.4000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 976.1200 0.8000 976.4200 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 965.1400 0.8000 965.4400 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 954.1600 0.8000 954.4600 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 943.7900 0.8000 944.0900 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 932.8100 0.8000 933.1100 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 921.8300 0.8000 922.1300 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 910.8500 0.8000 911.1500 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 899.8700 0.8000 900.1700 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 889.5000 0.8000 889.8000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 878.5200 0.8000 878.8200 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 867.5400 0.8000 867.8400 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 856.5600 0.8000 856.8600 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 845.5800 0.8000 845.8800 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 835.2100 0.8000 835.5100 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 824.2300 0.8000 824.5300 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 813.2500 0.8000 813.5500 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 802.2700 0.8000 802.5700 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 791.2900 0.8000 791.5900 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 780.9200 0.8000 781.2200 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 769.9400 0.8000 770.2400 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 758.9600 0.8000 759.2600 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 747.9800 0.8000 748.2800 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 737.0000 0.8000 737.3000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 726.6300 0.8000 726.9300 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 715.6500 0.8000 715.9500 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 704.6700 0.8000 704.9700 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 693.6900 0.8000 693.9900 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 682.7100 0.8000 683.0100 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 672.3400 0.8000 672.6400 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 661.3600 0.8000 661.6600 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 650.3800 0.8000 650.6800 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 639.4000 0.8000 639.7000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 628.4200 0.8000 628.7200 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 618.0500 0.8000 618.3500 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 607.0700 0.8000 607.3700 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 596.0900 0.8000 596.3900 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 585.1100 0.8000 585.4100 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 574.1300 0.8000 574.4300 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 563.7600 0.8000 564.0600 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 552.7800 0.8000 553.0800 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 541.8000 0.8000 542.1000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 530.8200 0.8000 531.1200 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 519.8400 0.8000 520.1400 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 509.4700 0.8000 509.7700 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 498.4900 0.8000 498.7900 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 487.5100 0.8000 487.8100 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 476.5300 0.8000 476.8300 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 465.5500 0.8000 465.8500 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 455.1800 0.8000 455.4800 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 444.2000 0.8000 444.5000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 433.2200 0.8000 433.5200 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 422.2400 0.8000 422.5400 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 411.2600 0.8000 411.5600 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 400.8900 0.8000 401.1900 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 389.9100 0.8000 390.2100 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 378.9300 0.8000 379.2300 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 367.9500 0.8000 368.2500 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 356.9700 0.8000 357.2700 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 346.6000 0.8000 346.9000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 335.6200 0.8000 335.9200 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 324.6400 0.8000 324.9400 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 313.6600 0.8000 313.9600 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 302.6800 0.8000 302.9800 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 292.3100 0.8000 292.6100 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 281.3300 0.8000 281.6300 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 270.3500 0.8000 270.6500 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 259.3700 0.8000 259.6700 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 248.3900 0.8000 248.6900 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 238.0200 0.8000 238.3200 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 227.0400 0.8000 227.3400 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 216.0600 0.8000 216.3600 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 205.0800 0.8000 205.3800 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 194.1000 0.8000 194.4000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 183.7300 0.8000 184.0300 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 172.7500 0.8000 173.0500 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 161.7700 0.8000 162.0700 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 150.7900 0.8000 151.0900 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 139.8100 0.8000 140.1100 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 129.4400 0.8000 129.7400 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 118.4600 0.8000 118.7600 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 107.4800 0.8000 107.7800 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 96.5000 0.8000 96.8000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 85.5200 0.8000 85.8200 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 75.1500 0.8000 75.4500 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 64.1700 0.8000 64.4700 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.0000 53.1900 0.8000 53.4900 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8724 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.448 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 141.944 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 757.504 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 42.2100 0.8000 42.5100 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 71.602 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 377.368 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 7.6218 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 41.12 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 31.2300 0.8000 31.5300 ;
    END
  END la_data_in[0]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 169.466 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 846.699 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 32.4325 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 153.9 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2847.5600 0.0000 2847.7000 0.4850 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 217.035 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1084.88 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.5328 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 25.6992 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 120.234 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2618.4800 0.0000 2618.6200 0.4850 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 338.107 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1690.14 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 7.4778 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.352 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 29.6738 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 160.127 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2389.4000 0.0000 2389.5400 0.4850 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 241.951 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1209.01 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 3.4608 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 18.928 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 35.8362 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 175.058 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 2160.7800 0.0000 2160.9200 0.4850 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 155.416 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 776.566 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4278 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 2.752 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 31.5203 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 151.496 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.55873 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 1931.7000 0.0000 1931.8400 0.4850 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0532 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 70.105 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 6.3096 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.592 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met3  ;
    ANTENNAMAXAREACAR 40.7845 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 203.833 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.566667 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1702.6200 0.0000 1702.7600 0.4850 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.0000 0.0000 1474.1400 0.4850 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 201.573 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1007.18 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.08 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 17.1094 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 92.192 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.4848 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 3.056 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 3.84762 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 24.254 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 1244.9200 0.0000 1245.0600 0.4850 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 36.236 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 180.901 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 7.5119 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 32.619 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1015.8400 0.0000 1015.9800 0.4850 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 38.9968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 194.705 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.2568 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.84 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met3  ;
    ANTENNAMAXAREACAR 5.74127 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 23.7222 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.725397 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 787.2200 0.0000 787.3600 0.4850 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 74.2654 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 370.93 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.1448 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 22.576 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 57.2171 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 281.948 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521429 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 558.1400 0.0000 558.2800 0.4850 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 77.8786 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 388.878 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.1249 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.136 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 2.6808 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 14.768 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.252 LAYER met4  ;
    ANTENNAMAXAREACAR 46.5075 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 226.464 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.521429 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 329.0600 0.0000 329.2000 0.4850 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 85.2472 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 425.957 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.262 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.864 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 0.6678 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 4.032 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 10.4302 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 50.7063 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 100.4400 0.0000 100.5800 0.4850 ;
    END
  END io_in[0]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 102.024 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 510.009 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2923.9200 0.0000 2924.0600 0.4850 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 156.205 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 780.797 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2694.8400 0.0000 2694.9800 0.4850 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 268.919 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1344.37 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2465.7600 0.0000 2465.9000 0.4850 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9056 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.33 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.9488 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.864 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2237.1400 0.0000 2237.2800 0.4850 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.8356 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 94.017 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7288 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.024 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2008.0600 0.0000 2008.2000 0.4850 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 19.9892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 99.785 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 25.0776 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 134.688 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1778.9800 0.0000 1779.1200 0.4850 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.564 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 74.6482 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 372.883 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 3.564 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.3948 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.576 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.7425 LAYER met3  ;
    ANTENNAMAXAREACAR 1.11987 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 5.08754 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.123098 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1549.9000 0.0000 1550.0400 0.4850 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 155.338 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 776.465 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1321.2800 0.0000 1321.4200 0.4850 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 152.258 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 761.065 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1092.2000 0.0000 1092.3400 0.4850 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 154.508 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 772.313 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 863.1200 0.0000 863.2600 0.4850 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 154.003 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 769.786 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 634.5000 0.0000 634.6400 0.4850 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3886 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 6.664 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 165.148 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 881.728 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 405.4200 0.0000 405.5600 0.4850 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 153.435 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 766.948 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 176.3400 0.0000 176.4800 0.4850 ;
    END
  END io_out[0]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 158.992 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 794.444 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.6388 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.544 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2999.8200 0.0000 2999.9600 0.4850 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 101.577 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 507.605 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.676 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.072 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 1.782 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 13.2948 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 71.376 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 2771.2000 0.0000 2771.3400 0.4850 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 103.382 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 516.747 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 9.8688 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 53.104 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2542.1200 0.0000 2542.2600 0.4850 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 27.011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 134.54 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 4.0728 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 22.192 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2313.0400 0.0000 2313.1800 0.4850 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.8303 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 103.926 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2084.4200 0.0000 2084.5600 0.4850 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 217.968 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1089.5 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1855.3400 0.0000 1855.4800 0.4850 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 514.031 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2741.97 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1626.2600 0.0000 1626.4000 0.4850 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.133 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.504 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 63.1848 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 337.456 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 1397.6400 0.0000 1397.7800 0.4850 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 158.373 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 791.641 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1168.5600 0.0000 1168.7000 0.4850 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 150.2 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 750.722 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 1.782 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 2.8788 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.824 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 939.4800 0.0000 939.6200 0.4850 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 159.07 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 795.127 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 710.8600 0.0000 711.0000 0.4850 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 156.083 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 780.188 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 481.7800 0.0000 481.9200 0.4850 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 156.905 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 784.297 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 252.7000 0.0000 252.8400 0.4850 ;
    END
  END io_oeb[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6283 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 19.816 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 4.5588 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 24.784 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.126 LAYER met4  ;
    ANTENNAMAXAREACAR 115.115 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 576.294 LAYER met4  ;
    ANTENNAMAXCUTCAR 1.04286 LAYER via4  ;
    PORT
      LAYER met3 ;
        RECT 0.0000 20.2500 0.8000 20.5500 ;
    END
  END user_clock2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 6.0000 6.0000 3364.4200 9.0000 ;
        RECT 1285.9400 176.0000 2448.7800 177.6000 ;
        RECT 1285.9400 135.7400 2388.6400 137.3400 ;
        RECT 1285.9400 405.6400 1948.2000 407.2400 ;
        RECT 1285.9400 864.9200 1948.2000 866.5200 ;
        RECT 1285.9400 635.2800 2448.7800 636.8800 ;
        RECT 1285.9400 1094.5600 2448.7800 1096.1600 ;
        RECT 6.0000 176.2600 1287.6800 177.8600 ;
        RECT 656.8450 405.9000 1067.4600 407.5000 ;
        RECT 6.0000 405.9000 516.5150 407.5000 ;
        RECT 1063.0600 6.0000 1064.6600 10.6000 ;
        RECT 1065.8600 136.0000 1287.6800 137.6000 ;
        RECT 1002.9200 186.3900 1010.9200 187.9900 ;
        RECT 1065.8600 144.7700 1071.0600 146.3700 ;
        RECT 1063.0600 174.6600 1064.6600 177.8600 ;
        RECT 1065.8600 169.1000 1071.0600 170.7000 ;
        RECT 1065.8600 186.2900 1071.0600 187.8900 ;
        RECT 1059.4600 186.3900 1067.4600 187.9900 ;
        RECT 1002.9200 397.8900 1010.9200 399.4900 ;
        RECT 1002.9200 416.0300 1010.9200 417.6300 ;
        RECT 1059.4600 397.8900 1067.4600 399.4900 ;
        RECT 1059.4600 416.0300 1067.4600 417.6300 ;
        RECT 1285.9400 144.5100 1291.1400 146.1100 ;
        RECT 1285.9400 168.8400 1291.1400 170.4400 ;
        RECT 1279.6800 169.1000 1287.6800 170.7000 ;
        RECT 1285.9400 186.0300 1291.1400 187.6300 ;
        RECT 1279.6800 186.2900 1287.6800 187.8900 ;
        RECT 1499.7600 144.5100 1507.7600 146.1100 ;
        RECT 1506.1600 144.5100 1511.3600 146.1100 ;
        RECT 1506.1600 168.8400 1511.3600 170.4400 ;
        RECT 1499.7600 168.8400 1507.7600 170.4400 ;
        RECT 1506.1600 186.0300 1511.3600 187.6300 ;
        RECT 1285.9400 397.7300 1291.1400 399.3300 ;
        RECT 1285.9400 415.6700 1291.1400 417.2700 ;
        RECT 1506.1600 415.6700 1511.3600 417.2700 ;
        RECT 1506.1600 397.7300 1511.3600 399.3300 ;
        RECT 1499.7600 397.7300 1507.7600 399.3300 ;
        RECT 6.0000 635.5400 1287.6800 637.1400 ;
        RECT 6.0000 865.1800 167.1150 866.7800 ;
        RECT 6.0000 1094.8200 167.1150 1096.4200 ;
        RECT 1002.9200 627.5300 1010.9200 629.1300 ;
        RECT 1002.9200 645.6700 1010.9200 647.2700 ;
        RECT 1065.8600 628.6800 1071.0600 630.2800 ;
        RECT 1063.0600 633.9400 1064.6600 637.1400 ;
        RECT 1059.4600 627.5300 1061.3600 629.1300 ;
        RECT 1059.4600 645.6700 1067.4600 647.2700 ;
        RECT 1065.8600 645.5700 1071.0600 647.1700 ;
        RECT 1002.9200 857.1700 1010.9200 858.7700 ;
        RECT 1059.4600 857.1700 1067.4600 858.7700 ;
        RECT 1285.9400 627.3700 1291.1400 628.9700 ;
        RECT 1285.9400 645.3100 1291.1400 646.9100 ;
        RECT 1279.6800 645.5700 1287.6800 647.1700 ;
        RECT 1279.6800 628.6800 1287.6800 630.2800 ;
        RECT 1499.7600 627.3700 1507.7600 628.9700 ;
        RECT 1499.7600 645.3100 1507.7600 646.9100 ;
        RECT 1506.1600 627.3700 1511.3600 628.9700 ;
        RECT 1506.1600 645.3100 1511.3600 646.9100 ;
        RECT 1499.7600 857.0100 1507.7600 858.6100 ;
        RECT 1506.1600 857.0100 1511.3600 858.6100 ;
        RECT 1285.9400 857.0100 1291.1400 858.6100 ;
        RECT 953.4450 1094.8200 1287.6800 1096.4200 ;
        RECT 953.4450 865.1800 1067.4600 866.7800 ;
        RECT 1002.9200 875.3100 1010.9200 876.9100 ;
        RECT 1059.4600 875.3100 1067.4600 876.9100 ;
        RECT 1002.9200 1104.9500 1010.9200 1106.5500 ;
        RECT 1002.9200 1086.8100 1010.9200 1088.4100 ;
        RECT 1059.4600 1086.8100 1061.3600 1088.4100 ;
        RECT 1065.8600 1087.9600 1071.0600 1089.5600 ;
        RECT 1063.0600 1093.2200 1064.6600 1096.4200 ;
        RECT 1059.4600 1104.9500 1067.4600 1106.5500 ;
        RECT 1065.8600 1104.8500 1071.0600 1106.4500 ;
        RECT 1285.9400 874.9500 1291.1400 876.5500 ;
        RECT 1499.7600 874.9500 1507.7600 876.5500 ;
        RECT 1506.1600 874.9500 1511.3600 876.5500 ;
        RECT 1285.9400 1086.6500 1291.1400 1088.2500 ;
        RECT 1279.6800 1087.9600 1287.6800 1089.5600 ;
        RECT 1285.9400 1104.5900 1291.1400 1106.1900 ;
        RECT 1279.6800 1104.8500 1287.6800 1106.4500 ;
        RECT 1506.1600 1086.6500 1511.3600 1088.2500 ;
        RECT 1499.7600 1086.6500 1507.7600 1088.2500 ;
        RECT 1506.1600 1104.5900 1511.3600 1106.1900 ;
        RECT 1726.3800 144.5100 1731.5800 146.1100 ;
        RECT 1726.3800 168.8400 1731.5800 170.4400 ;
        RECT 1719.9800 168.8400 1727.9800 170.4400 ;
        RECT 1726.3800 186.0300 1731.5800 187.6300 ;
        RECT 1946.6000 144.5100 1951.8000 146.1100 ;
        RECT 1946.6000 168.8400 1951.8000 170.4400 ;
        RECT 1940.2000 168.8400 1948.2000 170.4400 ;
        RECT 1946.6000 186.0300 1951.8000 187.6300 ;
        RECT 1726.3800 397.7300 1731.5800 399.3300 ;
        RECT 1719.9800 397.7300 1727.9800 399.3300 ;
        RECT 1726.3800 415.6700 1731.5800 417.2700 ;
        RECT 1719.9800 415.6700 1727.9800 417.2700 ;
        RECT 1940.2000 397.7300 1948.2000 399.3300 ;
        RECT 1940.2000 415.6700 1948.2000 417.2700 ;
        RECT 2166.8200 144.5100 2172.0200 146.1100 ;
        RECT 2160.4200 144.5100 2168.4200 146.1100 ;
        RECT 2166.8200 168.8400 2172.0200 170.4400 ;
        RECT 2160.4200 168.8400 2168.4200 170.4400 ;
        RECT 2166.8200 186.0300 2172.0200 187.6300 ;
        RECT 2380.6400 168.8400 2388.6400 170.4400 ;
        RECT 2387.0400 186.0300 2392.2400 187.6300 ;
        RECT 2166.8200 405.6400 2448.7800 407.2400 ;
        RECT 2166.8200 397.7300 2172.0200 399.3300 ;
        RECT 2166.8200 415.6700 2172.0200 417.2700 ;
        RECT 2387.0400 397.7300 2392.2400 399.3300 ;
        RECT 2380.6400 397.7300 2388.6400 399.3300 ;
        RECT 2387.0400 415.6700 2392.2400 417.2700 ;
        RECT 2380.6400 415.6700 2388.6400 417.2700 ;
        RECT 2440.7800 415.6700 2448.7800 417.2700 ;
        RECT 2440.7800 397.7300 2448.7800 399.3300 ;
        RECT 1719.9800 627.3700 1727.9800 628.9700 ;
        RECT 1726.3800 645.3100 1731.5800 646.9100 ;
        RECT 1726.3800 627.3700 1731.5800 628.9700 ;
        RECT 1719.9800 645.3100 1727.9800 646.9100 ;
        RECT 1946.6000 645.3100 1951.8000 646.9100 ;
        RECT 1946.6000 628.4200 1951.8000 630.0200 ;
        RECT 1940.2000 627.3700 1942.1000 628.9700 ;
        RECT 1943.8000 633.6800 1945.4000 636.8800 ;
        RECT 1940.2000 645.3100 1948.2000 646.9100 ;
        RECT 1726.3800 857.0100 1731.5800 858.6100 ;
        RECT 1940.2000 857.0100 1948.2000 858.6100 ;
        RECT 1719.9800 857.0100 1727.9800 858.6100 ;
        RECT 2166.8200 645.3100 2172.0200 646.9100 ;
        RECT 2160.4200 628.4200 2168.4200 630.0200 ;
        RECT 2166.8200 627.3700 2172.0200 628.9700 ;
        RECT 2387.0400 627.3700 2392.2400 628.9700 ;
        RECT 2387.0400 645.3100 2392.2400 646.9100 ;
        RECT 2380.6400 645.3100 2388.6400 646.9100 ;
        RECT 2380.6400 627.3700 2388.6400 628.9700 ;
        RECT 2440.7800 627.3700 2448.7800 628.9700 ;
        RECT 2440.7800 645.3100 2448.7800 646.9100 ;
        RECT 2166.8200 857.0100 2172.0200 858.6100 ;
        RECT 2387.0400 857.0100 2392.2400 858.6100 ;
        RECT 2440.7800 857.0100 2448.7800 858.6100 ;
        RECT 2380.6400 857.0100 2388.6400 858.6100 ;
        RECT 1726.3800 874.9500 1731.5800 876.5500 ;
        RECT 1719.9800 874.9500 1727.9800 876.5500 ;
        RECT 1940.2000 874.9500 1948.2000 876.5500 ;
        RECT 1719.9800 1086.6500 1727.9800 1088.2500 ;
        RECT 1726.3800 1086.6500 1731.5800 1088.2500 ;
        RECT 1726.3800 1104.5900 1731.5800 1106.1900 ;
        RECT 1719.9800 1104.5900 1727.9800 1106.1900 ;
        RECT 1946.6000 1104.5900 1951.8000 1106.1900 ;
        RECT 1946.6000 1087.7000 1951.8000 1089.3000 ;
        RECT 1940.2000 1086.6500 1942.1000 1088.2500 ;
        RECT 1943.8000 1092.9600 1945.4000 1096.1600 ;
        RECT 1940.2000 1104.5900 1948.2000 1106.1900 ;
        RECT 2166.8200 864.9200 2448.7800 866.5200 ;
        RECT 2166.8200 874.9500 2172.0200 876.5500 ;
        RECT 2387.0400 874.9500 2392.2400 876.5500 ;
        RECT 2440.7800 874.9500 2448.7800 876.5500 ;
        RECT 2380.6400 874.9500 2388.6400 876.5500 ;
        RECT 2160.4200 1087.7000 2168.4200 1089.3000 ;
        RECT 2166.8200 1086.6500 2172.0200 1088.2500 ;
        RECT 2166.8200 1104.5900 2172.0200 1106.1900 ;
        RECT 2380.6400 1104.5900 2388.6400 1106.1900 ;
        RECT 2387.0400 1104.5900 2392.2400 1106.1900 ;
        RECT 2387.0400 1086.6500 2392.2400 1088.2500 ;
        RECT 2380.6400 1086.6500 2388.6400 1088.2500 ;
        RECT 2440.7800 1104.5900 2448.7800 1106.1900 ;
        RECT 2440.7800 1086.6500 2448.7800 1088.2500 ;
        RECT 6.0000 2560.7200 3364.4200 2563.7200 ;
        RECT 1065.8600 2472.4000 2388.6400 2474.0000 ;
        RECT 1285.9400 2013.1200 2448.7800 2014.7200 ;
        RECT 1285.9400 1553.8400 2448.7800 1555.4400 ;
        RECT 1285.9400 2242.7600 1948.2000 2244.3600 ;
        RECT 1285.9400 1783.4800 1948.2000 1785.0800 ;
        RECT 1285.9400 1324.2000 1948.2000 1325.8000 ;
        RECT 6.0000 2013.3800 1287.6800 2014.9800 ;
        RECT 6.0000 1324.4600 167.1150 1326.0600 ;
        RECT 6.0000 1554.1000 167.1150 1555.7000 ;
        RECT 152.4900 1558.8300 154.5200 1559.3100 ;
        RECT 6.0000 1783.7400 167.1150 1785.3400 ;
        RECT 953.4450 1554.1000 1287.6800 1555.7000 ;
        RECT 953.4450 1324.4600 1067.4600 1326.0600 ;
        RECT 1002.9200 1334.5900 1010.9200 1336.1900 ;
        RECT 1002.9200 1316.4500 1010.9200 1318.0500 ;
        RECT 1059.4600 1334.5900 1067.4600 1336.1900 ;
        RECT 1059.4600 1316.4500 1067.4600 1318.0500 ;
        RECT 1002.9200 1564.2300 1010.9200 1565.8300 ;
        RECT 1002.9200 1546.0900 1010.9200 1547.6900 ;
        RECT 1065.8600 1547.2400 1071.0600 1548.8400 ;
        RECT 1059.4600 1546.0900 1061.3600 1547.6900 ;
        RECT 1059.4600 1564.2300 1067.4600 1565.8300 ;
        RECT 1063.0600 1552.5000 1064.6600 1555.7000 ;
        RECT 1065.8600 1564.1300 1071.0600 1565.7300 ;
        RECT 1285.9400 1334.2300 1291.1400 1335.8300 ;
        RECT 1285.9400 1316.2900 1291.1400 1317.8900 ;
        RECT 1506.1600 1316.2900 1511.3600 1317.8900 ;
        RECT 1499.7600 1334.2300 1507.7600 1335.8300 ;
        RECT 1499.7600 1316.2900 1507.7600 1317.8900 ;
        RECT 1506.1600 1334.2300 1511.3600 1335.8300 ;
        RECT 1279.6800 1547.2400 1287.6800 1548.8400 ;
        RECT 1285.9400 1545.9300 1291.1400 1547.5300 ;
        RECT 1285.9400 1563.8700 1291.1400 1565.4700 ;
        RECT 1279.6800 1564.1300 1287.6800 1565.7300 ;
        RECT 1499.7600 1545.9300 1507.7600 1547.5300 ;
        RECT 1506.1600 1545.9300 1511.3600 1547.5300 ;
        RECT 1506.1600 1563.8700 1511.3600 1565.4700 ;
        RECT 1499.7600 1563.8700 1507.7600 1565.4700 ;
        RECT 953.4450 1783.7400 1067.4600 1785.3400 ;
        RECT 1002.9200 1775.7300 1010.9200 1777.3300 ;
        RECT 1002.9200 1793.8700 1010.9200 1795.4700 ;
        RECT 1059.4600 1775.7300 1067.4600 1777.3300 ;
        RECT 1059.4600 1793.8700 1067.4600 1795.4700 ;
        RECT 1002.9200 2005.3700 1010.9200 2006.9700 ;
        RECT 1002.9200 2023.5100 1010.9200 2025.1100 ;
        RECT 1065.8600 2006.5200 1071.0600 2008.1200 ;
        RECT 1059.4600 2005.3700 1061.3600 2006.9700 ;
        RECT 1063.0600 2011.7800 1064.6600 2014.9800 ;
        RECT 1065.8600 2023.4100 1071.0600 2025.0100 ;
        RECT 1285.9400 1793.5100 1291.1400 1795.1100 ;
        RECT 1285.9400 1775.5700 1291.1400 1777.1700 ;
        RECT 1499.7600 1775.5700 1507.7600 1777.1700 ;
        RECT 1506.1600 1775.5700 1511.3600 1777.1700 ;
        RECT 1506.1600 1793.5100 1511.3600 1795.1100 ;
        RECT 1499.7600 1793.5100 1507.7600 1795.1100 ;
        RECT 1285.9400 2005.2100 1291.1400 2006.8100 ;
        RECT 1279.6800 2006.5200 1287.6800 2008.1200 ;
        RECT 1285.9400 2023.1500 1291.1400 2024.7500 ;
        RECT 1279.6800 2023.4100 1287.6800 2025.0100 ;
        RECT 1506.1600 2005.2100 1511.3600 2006.8100 ;
        RECT 1499.7600 2005.2100 1507.7600 2006.8100 ;
        RECT 1499.7600 2023.1500 1507.7600 2024.7500 ;
        RECT 1506.1600 2023.1500 1511.3600 2024.7500 ;
        RECT 6.0000 2243.0200 1067.4600 2244.6200 ;
        RECT 1002.9200 2235.0100 1010.9200 2236.6100 ;
        RECT 1002.9200 2253.1500 1010.9200 2254.7500 ;
        RECT 1059.4600 2253.1500 1067.4600 2254.7500 ;
        RECT 1059.4600 2235.0100 1067.4600 2236.6100 ;
        RECT 1002.9200 2464.6500 1010.9200 2466.2500 ;
        RECT 1065.8600 2465.8000 1071.0600 2467.4000 ;
        RECT 1059.4600 2464.6500 1061.3600 2466.2500 ;
        RECT 1065.8600 2481.1700 1070.9200 2482.7700 ;
        RECT 1065.8600 2505.5000 1070.9200 2507.1000 ;
        RECT 1285.9400 2252.7900 1291.1400 2254.3900 ;
        RECT 1285.9400 2234.8500 1291.1400 2236.4500 ;
        RECT 1506.1600 2234.8500 1511.3600 2236.4500 ;
        RECT 1506.1600 2252.7900 1511.3600 2254.3900 ;
        RECT 1499.7600 2252.7900 1507.7600 2254.3900 ;
        RECT 1499.7600 2234.8500 1507.7600 2236.4500 ;
        RECT 1300.4600 2458.3800 1302.0600 2458.6200 ;
        RECT 1285.9400 2464.4900 1291.1400 2466.0900 ;
        RECT 1279.6800 2465.8000 1287.6800 2467.4000 ;
        RECT 1285.9400 2481.1700 1291.1400 2482.7700 ;
        RECT 1279.5400 2481.1700 1287.6800 2482.7700 ;
        RECT 1285.9400 2505.5000 1291.1400 2507.1000 ;
        RECT 1279.5400 2505.5000 1287.6800 2507.1000 ;
        RECT 1520.6800 2458.3800 1522.2800 2458.6200 ;
        RECT 1499.7600 2464.4900 1507.7600 2466.0900 ;
        RECT 1506.1600 2464.4900 1511.3600 2466.0900 ;
        RECT 1506.1600 2481.1700 1511.3600 2482.7700 ;
        RECT 1499.7600 2481.1700 1507.7600 2482.7700 ;
        RECT 1506.1600 2505.5000 1511.3600 2507.1000 ;
        RECT 1499.7600 2505.5000 1507.7600 2507.1000 ;
        RECT 1062.9200 2559.1200 1064.5200 2563.7200 ;
        RECT 1063.0600 2559.1200 1064.6600 2563.7200 ;
        RECT 1719.9800 1316.2900 1727.9800 1317.8900 ;
        RECT 1726.3800 1334.2300 1731.5800 1335.8300 ;
        RECT 1726.3800 1316.2900 1731.5800 1317.8900 ;
        RECT 1719.9800 1334.2300 1727.9800 1335.8300 ;
        RECT 1940.2000 1334.2300 1948.2000 1335.8300 ;
        RECT 1940.2000 1316.2900 1948.2000 1317.8900 ;
        RECT 1726.3800 1545.9300 1731.5800 1547.5300 ;
        RECT 1719.9800 1545.9300 1727.9800 1547.5300 ;
        RECT 1719.9800 1563.8700 1727.9800 1565.4700 ;
        RECT 1726.3800 1563.8700 1731.5800 1565.4700 ;
        RECT 1946.6000 1546.9800 1951.8000 1548.5800 ;
        RECT 1940.2000 1545.9300 1942.1000 1547.5300 ;
        RECT 1946.6000 1563.8700 1951.8000 1565.4700 ;
        RECT 1940.2000 1563.8700 1948.2000 1565.4700 ;
        RECT 1943.8000 1552.2400 1945.4000 1555.4400 ;
        RECT 2166.8200 1324.2000 2448.7800 1325.8000 ;
        RECT 2166.8200 1334.2300 2172.0200 1335.8300 ;
        RECT 2166.8200 1316.2900 2172.0200 1317.8900 ;
        RECT 2387.0400 1316.2900 2392.2400 1317.8900 ;
        RECT 2380.6400 1316.2900 2388.6400 1317.8900 ;
        RECT 2380.6400 1334.2300 2388.6400 1335.8300 ;
        RECT 2387.0400 1334.2300 2392.2400 1335.8300 ;
        RECT 2440.7800 1316.2900 2448.7800 1317.8900 ;
        RECT 2440.7800 1334.2300 2448.7800 1335.8300 ;
        RECT 2160.4200 1546.9800 2168.4200 1548.5800 ;
        RECT 2166.8200 1545.9300 2172.0200 1547.5300 ;
        RECT 2166.8200 1563.8700 2172.0200 1565.4700 ;
        RECT 2160.4200 1563.8700 2168.4200 1565.4700 ;
        RECT 2380.6400 1563.8700 2388.6400 1565.4700 ;
        RECT 2387.0400 1563.8700 2392.2400 1565.4700 ;
        RECT 2380.6400 1545.9300 2388.6400 1547.5300 ;
        RECT 2387.0400 1545.9300 2392.2400 1547.5300 ;
        RECT 2440.7800 1563.8700 2448.7800 1565.4700 ;
        RECT 2440.7800 1545.9300 2448.7800 1547.5300 ;
        RECT 1719.9800 1775.5700 1727.9800 1777.1700 ;
        RECT 1726.3800 1793.5100 1731.5800 1795.1100 ;
        RECT 1726.3800 1775.5700 1731.5800 1777.1700 ;
        RECT 1719.9800 1793.5100 1727.9800 1795.1100 ;
        RECT 1940.2000 1793.5100 1948.2000 1795.1100 ;
        RECT 1940.2000 1775.5700 1948.2000 1777.1700 ;
        RECT 1719.9800 2005.2100 1727.9800 2006.8100 ;
        RECT 1726.3800 2005.2100 1731.5800 2006.8100 ;
        RECT 1726.3800 2023.1500 1731.5800 2024.7500 ;
        RECT 1719.9800 2023.1500 1727.9800 2024.7500 ;
        RECT 1946.6000 2006.2600 1951.8000 2007.8600 ;
        RECT 1943.8000 2011.5200 1945.4000 2014.7200 ;
        RECT 1940.2000 2005.2100 1942.1000 2006.8100 ;
        RECT 1940.2000 2023.1500 1948.2000 2024.7500 ;
        RECT 1946.6000 2023.1500 1951.8000 2024.7500 ;
        RECT 2166.8200 1783.4800 2448.7800 1785.0800 ;
        RECT 2166.8200 1793.5100 2172.0200 1795.1100 ;
        RECT 2166.8200 1775.5700 2172.0200 1777.1700 ;
        RECT 2380.6400 1775.5700 2388.6400 1777.1700 ;
        RECT 2387.0400 1775.5700 2392.2400 1777.1700 ;
        RECT 2387.0400 1793.5100 2392.2400 1795.1100 ;
        RECT 2440.7800 1775.5700 2448.7800 1777.1700 ;
        RECT 2440.7800 1793.5100 2448.7800 1795.1100 ;
        RECT 2160.4200 2006.2600 2168.4200 2007.8600 ;
        RECT 2166.8200 2005.2100 2172.0200 2006.8100 ;
        RECT 2166.8200 2023.1500 2172.0200 2024.7500 ;
        RECT 2380.6400 2005.2100 2388.6400 2006.8100 ;
        RECT 2387.0400 2005.2100 2392.2400 2006.8100 ;
        RECT 2440.7800 2005.2100 2448.7800 2006.8100 ;
        RECT 2387.0400 2023.1500 2392.2400 2024.7500 ;
        RECT 2380.6400 2023.1500 2388.6400 2024.7500 ;
        RECT 2440.7800 2023.1500 2448.7800 2024.7500 ;
        RECT 1719.9800 2234.8500 1727.9800 2236.4500 ;
        RECT 1719.9800 2252.7900 1727.9800 2254.3900 ;
        RECT 1726.3800 2252.7900 1731.5800 2254.3900 ;
        RECT 1726.3800 2234.8500 1731.5800 2236.4500 ;
        RECT 1940.2000 2252.7900 1948.2000 2254.3900 ;
        RECT 1940.2000 2234.8500 1948.2000 2236.4500 ;
        RECT 1719.9800 2464.4900 1727.9800 2466.0900 ;
        RECT 1726.3800 2464.4900 1731.5800 2466.0900 ;
        RECT 1726.3800 2481.1700 1731.5800 2482.7700 ;
        RECT 1740.9000 2458.3800 1742.5000 2458.6200 ;
        RECT 1726.3800 2505.5000 1731.5800 2507.1000 ;
        RECT 1719.9800 2505.5000 1727.9800 2507.1000 ;
        RECT 1946.6000 2481.1700 1951.8000 2482.7700 ;
        RECT 1946.6000 2465.5400 1951.8000 2467.1400 ;
        RECT 1940.2000 2464.4900 1942.1000 2466.0900 ;
        RECT 1943.8000 2470.8000 1945.4000 2474.0000 ;
        RECT 1946.6000 2505.5000 1951.8000 2507.1000 ;
        RECT 1940.2000 2505.5000 1948.2000 2507.1000 ;
        RECT 2166.8200 2242.7600 2448.7800 2244.3600 ;
        RECT 2166.8200 2252.7900 2172.0200 2254.3900 ;
        RECT 2166.8200 2234.8500 2172.0200 2236.4500 ;
        RECT 2387.0400 2252.7900 2392.2400 2254.3900 ;
        RECT 2387.0400 2234.8500 2392.2400 2236.4500 ;
        RECT 2380.6400 2234.8500 2388.6400 2236.4500 ;
        RECT 2440.7800 2234.8500 2448.7800 2236.4500 ;
        RECT 2440.7800 2252.7900 2448.7800 2254.3900 ;
        RECT 2166.8200 2464.4900 2172.0200 2466.0900 ;
        RECT 2181.3400 2458.3800 2182.9400 2458.6200 ;
        RECT 2160.4200 2465.5400 2168.4200 2467.1400 ;
        RECT 2166.8200 2481.1700 2172.0200 2482.7700 ;
        RECT 2166.8200 2505.5000 2172.0200 2507.1000 ;
        RECT 2160.4200 2505.5000 2168.4200 2507.1000 ;
        RECT 2387.0400 2464.4900 2392.2400 2466.0900 ;
        RECT 2380.6400 2464.4900 2388.6400 2466.0900 ;
        RECT 2380.6400 2505.5000 2388.6400 2507.1000 ;
        RECT 2440.7800 2464.4900 2448.7800 2466.0900 ;
        RECT 152.2400 1558.8300 152.7400 1559.3100 ;
        RECT 665.7200 442.1000 667.3200 442.5800 ;
        RECT 502.9200 442.1000 504.5200 442.5800 ;
        RECT 6.0000 442.1000 9.0000 442.5800 ;
        RECT 1002.9200 442.1000 1004.5200 442.5800 ;
        RECT 6.0000 12.3400 9.0000 12.8200 ;
        RECT 6.0000 17.7800 9.0000 18.2600 ;
        RECT 6.0000 34.1000 9.0000 34.5800 ;
        RECT 6.0000 23.2200 9.0000 23.7000 ;
        RECT 6.0000 28.6600 9.0000 29.1400 ;
        RECT 6.0000 39.5400 9.0000 40.0200 ;
        RECT 6.0000 44.9800 9.0000 45.4600 ;
        RECT 6.0000 50.4200 9.0000 50.9000 ;
        RECT 6.0000 55.8600 9.0000 56.3400 ;
        RECT 6.0000 61.3000 9.0000 61.7800 ;
        RECT 6.0000 66.7400 9.0000 67.2200 ;
        RECT 6.0000 72.1800 9.0000 72.6600 ;
        RECT 6.0000 77.6200 9.0000 78.1000 ;
        RECT 6.0000 83.0600 9.0000 83.5400 ;
        RECT 6.0000 88.5000 9.0000 88.9800 ;
        RECT 6.0000 93.9400 9.0000 94.4200 ;
        RECT 6.0000 99.3800 9.0000 99.8600 ;
        RECT 6.0000 104.8200 9.0000 105.3000 ;
        RECT 6.0000 110.2600 9.0000 110.7400 ;
        RECT 6.0000 115.7000 9.0000 116.1800 ;
        RECT 6.0000 121.1400 9.0000 121.6200 ;
        RECT 6.0000 126.5800 9.0000 127.0600 ;
        RECT 6.0000 132.0200 9.0000 132.5000 ;
        RECT 6.0000 137.4600 9.0000 137.9400 ;
        RECT 6.0000 142.9000 9.0000 143.3800 ;
        RECT 6.0000 148.3400 9.0000 148.8200 ;
        RECT 6.0000 153.7800 9.0000 154.2600 ;
        RECT 6.0000 159.2200 9.0000 159.7000 ;
        RECT 6.0000 164.6600 9.0000 165.1400 ;
        RECT 6.0000 170.1000 9.0000 170.5800 ;
        RECT 6.0000 175.3700 9.0000 175.8500 ;
        RECT 6.0000 191.8600 9.0000 192.3400 ;
        RECT 6.0000 180.9800 9.0000 181.4600 ;
        RECT 6.0000 186.4200 9.0000 186.9000 ;
        RECT 6.0000 197.3000 9.0000 197.7800 ;
        RECT 6.0000 202.7400 9.0000 203.2200 ;
        RECT 6.0000 208.1800 9.0000 208.6600 ;
        RECT 6.0000 213.6200 9.0000 214.1000 ;
        RECT 6.0000 219.0600 9.0000 219.5400 ;
        RECT 6.0000 224.5000 9.0000 224.9800 ;
        RECT 6.0000 229.9400 9.0000 230.4200 ;
        RECT 6.0000 235.3800 9.0000 235.8600 ;
        RECT 6.0000 240.8200 9.0000 241.3000 ;
        RECT 6.0000 246.2600 9.0000 246.7400 ;
        RECT 6.0000 251.7000 9.0000 252.1800 ;
        RECT 6.0000 257.1400 9.0000 257.6200 ;
        RECT 6.0000 262.5800 9.0000 263.0600 ;
        RECT 6.0000 268.0200 9.0000 268.5000 ;
        RECT 6.0000 273.4600 9.0000 273.9400 ;
        RECT 6.0000 278.9000 9.0000 279.3800 ;
        RECT 6.0000 284.3400 9.0000 284.8200 ;
        RECT 6.0000 289.7800 9.0000 290.2600 ;
        RECT 6.0000 295.2200 9.0000 295.7000 ;
        RECT 6.0000 300.6600 9.0000 301.1400 ;
        RECT 6.0000 306.1000 9.0000 306.5800 ;
        RECT 6.0000 311.5400 9.0000 312.0200 ;
        RECT 6.0000 316.9800 9.0000 317.4600 ;
        RECT 6.0000 322.4200 9.0000 322.9000 ;
        RECT 6.0000 327.8600 9.0000 328.3400 ;
        RECT 6.0000 333.3000 9.0000 333.7800 ;
        RECT 6.0000 349.6200 9.0000 350.1000 ;
        RECT 6.0000 338.7400 9.0000 339.2200 ;
        RECT 6.0000 344.1800 9.0000 344.6600 ;
        RECT 6.0000 355.0600 9.0000 355.5400 ;
        RECT 6.0000 360.5000 9.0000 360.9800 ;
        RECT 6.0000 365.9400 9.0000 366.4200 ;
        RECT 6.0000 371.3800 9.0000 371.8600 ;
        RECT 6.0000 376.8200 9.0000 377.3000 ;
        RECT 6.0000 382.2600 9.0000 382.7400 ;
        RECT 6.0000 387.7000 9.0000 388.1800 ;
        RECT 6.0000 393.1400 9.0000 393.6200 ;
        RECT 6.0000 398.5800 9.0000 399.0600 ;
        RECT 6.0000 404.0200 9.0000 404.5000 ;
        RECT 6.0000 414.9000 9.0000 415.3800 ;
        RECT 6.0000 410.5600 9.0000 411.0400 ;
        RECT 6.0000 420.3400 9.0000 420.8200 ;
        RECT 6.0000 425.7800 9.0000 426.2600 ;
        RECT 6.0000 431.2200 9.0000 431.7000 ;
        RECT 6.0000 436.6600 9.0000 437.1400 ;
        RECT 502.9200 191.8600 504.5200 192.3400 ;
        RECT 502.9200 186.4200 504.5200 186.9000 ;
        RECT 502.9200 180.9800 504.5200 181.4600 ;
        RECT 502.9200 197.3000 504.5200 197.7800 ;
        RECT 502.9200 202.7400 504.5200 203.2200 ;
        RECT 502.9200 208.1800 504.5200 208.6600 ;
        RECT 502.9200 213.6200 504.5200 214.1000 ;
        RECT 502.9200 219.0600 504.5200 219.5400 ;
        RECT 502.9200 224.5000 504.5200 224.9800 ;
        RECT 502.9200 229.9400 504.5200 230.4200 ;
        RECT 665.7200 191.8600 667.3200 192.3400 ;
        RECT 665.7200 186.4200 667.3200 186.9000 ;
        RECT 665.7200 180.9800 667.3200 181.4600 ;
        RECT 665.7200 197.3000 667.3200 197.7800 ;
        RECT 665.7200 202.7400 667.3200 203.2200 ;
        RECT 665.7200 208.1800 667.3200 208.6600 ;
        RECT 665.7200 213.6200 667.3200 214.1000 ;
        RECT 665.7200 219.0600 667.3200 219.5400 ;
        RECT 665.7200 224.5000 667.3200 224.9800 ;
        RECT 665.7200 229.9400 667.3200 230.4200 ;
        RECT 502.9200 235.3800 504.5200 235.8600 ;
        RECT 502.9200 240.8200 504.5200 241.3000 ;
        RECT 502.9200 246.2600 504.5200 246.7400 ;
        RECT 502.9200 251.7000 504.5200 252.1800 ;
        RECT 502.9200 257.1400 504.5200 257.6200 ;
        RECT 502.9200 262.5800 504.5200 263.0600 ;
        RECT 502.9200 268.0200 504.5200 268.5000 ;
        RECT 502.9200 273.4600 504.5200 273.9400 ;
        RECT 502.9200 278.9000 504.5200 279.3800 ;
        RECT 502.9200 284.3400 504.5200 284.8200 ;
        RECT 502.9200 289.7800 504.5200 290.2600 ;
        RECT 502.9200 295.2200 504.5200 295.7000 ;
        RECT 502.9200 300.6600 504.5200 301.1400 ;
        RECT 502.9200 306.1000 504.5200 306.5800 ;
        RECT 502.9200 311.5400 504.5200 312.0200 ;
        RECT 502.9200 316.9800 504.5200 317.4600 ;
        RECT 502.9200 322.4200 504.5200 322.9000 ;
        RECT 502.9200 327.8600 504.5200 328.3400 ;
        RECT 502.9200 333.3000 504.5200 333.7800 ;
        RECT 502.9200 349.6200 504.5200 350.1000 ;
        RECT 502.9200 338.7400 504.5200 339.2200 ;
        RECT 502.9200 344.1800 504.5200 344.6600 ;
        RECT 502.9200 355.0600 504.5200 355.5400 ;
        RECT 502.9200 360.5000 504.5200 360.9800 ;
        RECT 502.9200 365.9400 504.5200 366.4200 ;
        RECT 502.9200 371.3800 504.5200 371.8600 ;
        RECT 502.9200 376.8200 504.5200 377.3000 ;
        RECT 502.9200 382.2600 504.5200 382.7400 ;
        RECT 502.9200 387.7000 504.5200 388.1800 ;
        RECT 502.9200 393.1400 504.5200 393.6200 ;
        RECT 502.9200 398.5800 504.5200 399.0600 ;
        RECT 502.9200 414.9000 504.5200 415.3800 ;
        RECT 502.9200 410.5600 504.5200 411.0400 ;
        RECT 502.9200 404.0200 504.5200 404.5000 ;
        RECT 502.9200 420.3400 504.5200 420.8200 ;
        RECT 502.9200 425.7800 504.5200 426.2600 ;
        RECT 502.9200 431.2200 504.5200 431.7000 ;
        RECT 502.9200 436.6600 504.5200 437.1400 ;
        RECT 665.7200 235.3800 667.3200 235.8600 ;
        RECT 665.7200 240.8200 667.3200 241.3000 ;
        RECT 665.7200 246.2600 667.3200 246.7400 ;
        RECT 665.7200 251.7000 667.3200 252.1800 ;
        RECT 665.7200 257.1400 667.3200 257.6200 ;
        RECT 665.7200 262.5800 667.3200 263.0600 ;
        RECT 665.7200 268.0200 667.3200 268.5000 ;
        RECT 665.7200 273.4600 667.3200 273.9400 ;
        RECT 665.7200 278.9000 667.3200 279.3800 ;
        RECT 665.7200 284.3400 667.3200 284.8200 ;
        RECT 665.7200 289.7800 667.3200 290.2600 ;
        RECT 665.7200 295.2200 667.3200 295.7000 ;
        RECT 665.7200 300.6600 667.3200 301.1400 ;
        RECT 665.7200 306.1000 667.3200 306.5800 ;
        RECT 665.7200 311.5400 667.3200 312.0200 ;
        RECT 665.7200 316.9800 667.3200 317.4600 ;
        RECT 665.7200 322.4200 667.3200 322.9000 ;
        RECT 665.7200 327.8600 667.3200 328.3400 ;
        RECT 665.7200 333.3000 667.3200 333.7800 ;
        RECT 665.7200 349.6200 667.3200 350.1000 ;
        RECT 665.7200 338.7400 667.3200 339.2200 ;
        RECT 665.7200 344.1800 667.3200 344.6600 ;
        RECT 665.7200 355.0600 667.3200 355.5400 ;
        RECT 665.7200 360.5000 667.3200 360.9800 ;
        RECT 665.7200 365.9400 667.3200 366.4200 ;
        RECT 665.7200 371.3800 667.3200 371.8600 ;
        RECT 665.7200 376.8200 667.3200 377.3000 ;
        RECT 665.7200 382.2600 667.3200 382.7400 ;
        RECT 665.7200 387.7000 667.3200 388.1800 ;
        RECT 665.7200 393.1400 667.3200 393.6200 ;
        RECT 665.7200 398.5800 667.3200 399.0600 ;
        RECT 665.7200 404.0200 667.3200 404.5000 ;
        RECT 665.7200 410.5600 667.3200 411.0400 ;
        RECT 665.7200 414.9000 667.3200 415.3800 ;
        RECT 665.7200 420.3400 667.3200 420.8200 ;
        RECT 665.7200 425.7800 667.3200 426.2600 ;
        RECT 665.7200 431.2200 667.3200 431.7000 ;
        RECT 665.7200 436.6600 667.3200 437.1400 ;
        RECT 1065.8600 12.3400 1067.4600 12.8200 ;
        RECT 1065.8600 17.7800 1067.4600 18.2600 ;
        RECT 1285.9400 12.3400 1287.6800 12.8200 ;
        RECT 1285.9400 17.7800 1287.6800 18.2600 ;
        RECT 1506.1600 12.3400 1507.7600 12.8200 ;
        RECT 1506.1600 17.7800 1507.7600 18.2600 ;
        RECT 1002.9200 191.8600 1004.5200 192.3400 ;
        RECT 1002.9200 180.9800 1004.5200 181.4600 ;
        RECT 1002.9200 197.3000 1004.5200 197.7800 ;
        RECT 1002.9200 202.7400 1004.5200 203.2200 ;
        RECT 1002.9200 208.1800 1004.5200 208.6600 ;
        RECT 1002.9200 213.6200 1004.5200 214.1000 ;
        RECT 1002.9200 219.0600 1004.5200 219.5400 ;
        RECT 1002.9200 224.5000 1004.5200 224.9800 ;
        RECT 1002.9200 229.9400 1004.5200 230.4200 ;
        RECT 1065.8600 34.1000 1067.4600 34.5800 ;
        RECT 1065.8600 28.6600 1067.4600 29.1400 ;
        RECT 1065.8600 23.2200 1067.4600 23.7000 ;
        RECT 1065.8600 39.5400 1067.4600 40.0200 ;
        RECT 1065.8600 44.9800 1067.4600 45.4600 ;
        RECT 1065.8600 50.4200 1067.4600 50.9000 ;
        RECT 1065.8600 55.8600 1067.4600 56.3400 ;
        RECT 1065.8600 61.3000 1067.4600 61.7800 ;
        RECT 1065.8600 66.7400 1067.4600 67.2200 ;
        RECT 1065.8600 72.1800 1067.4600 72.6600 ;
        RECT 1065.8600 77.6200 1067.4600 78.1000 ;
        RECT 1065.8600 83.0600 1067.4600 83.5400 ;
        RECT 1065.8600 88.5000 1067.4600 88.9800 ;
        RECT 1065.8600 93.9400 1067.4600 94.4200 ;
        RECT 1065.8600 99.3800 1067.4600 99.8600 ;
        RECT 1065.8600 110.2600 1067.4600 110.7400 ;
        RECT 1065.8600 104.8200 1067.4600 105.3000 ;
        RECT 1065.8600 115.7000 1067.4600 116.1800 ;
        RECT 1065.8600 121.1400 1067.4600 121.6200 ;
        RECT 1065.8600 126.5800 1067.4600 127.0600 ;
        RECT 1065.8600 132.0200 1067.4600 132.5000 ;
        RECT 1065.8600 136.0000 1067.4600 137.9400 ;
        RECT 1065.8600 142.9000 1067.4600 143.3800 ;
        RECT 1065.8600 149.1900 1067.4600 149.6700 ;
        RECT 1065.8600 153.7800 1067.4600 154.2600 ;
        RECT 1065.8600 159.2200 1067.4600 159.7000 ;
        RECT 1065.8600 164.6600 1067.4600 165.1400 ;
        RECT 1073.3200 163.7000 1074.9200 164.1800 ;
        RECT 1065.8600 186.2900 1067.4600 187.9900 ;
        RECT 1002.9200 235.3800 1004.5200 235.8600 ;
        RECT 1002.9200 240.8200 1004.5200 241.3000 ;
        RECT 1002.9200 246.2600 1004.5200 246.7400 ;
        RECT 1002.9200 251.7000 1004.5200 252.1800 ;
        RECT 1002.9200 257.1400 1004.5200 257.6200 ;
        RECT 1002.9200 268.0200 1004.5200 268.5000 ;
        RECT 1002.9200 262.5800 1004.5200 263.0600 ;
        RECT 1002.9200 273.4600 1004.5200 273.9400 ;
        RECT 1002.9200 278.9000 1004.5200 279.3800 ;
        RECT 1002.9200 284.3400 1004.5200 284.8200 ;
        RECT 1002.9200 289.7800 1004.5200 290.2600 ;
        RECT 1002.9200 295.2200 1004.5200 295.7000 ;
        RECT 1002.9200 300.6600 1004.5200 301.1400 ;
        RECT 1002.9200 306.1000 1004.5200 306.5800 ;
        RECT 1002.9200 311.5400 1004.5200 312.0200 ;
        RECT 1002.9200 316.9800 1004.5200 317.4600 ;
        RECT 1002.9200 322.4200 1004.5200 322.9000 ;
        RECT 1002.9200 327.8600 1004.5200 328.3400 ;
        RECT 1002.9200 333.3000 1004.5200 333.7800 ;
        RECT 1002.9200 349.6200 1004.5200 350.1000 ;
        RECT 1002.9200 344.1800 1004.5200 344.6600 ;
        RECT 1002.9200 338.7400 1004.5200 339.2200 ;
        RECT 1002.9200 355.0600 1004.5200 355.5400 ;
        RECT 1002.9200 360.5000 1004.5200 360.9800 ;
        RECT 1002.9200 371.3800 1004.5200 371.8600 ;
        RECT 1002.9200 365.9400 1004.5200 366.4200 ;
        RECT 1002.9200 376.8200 1004.5200 377.3000 ;
        RECT 1002.9200 382.2600 1004.5200 382.7400 ;
        RECT 1002.9200 387.7000 1004.5200 388.1800 ;
        RECT 1002.9200 393.1400 1004.5200 393.6200 ;
        RECT 1013.1800 391.6400 1014.7800 392.1200 ;
        RECT 1002.9200 404.0200 1004.5200 404.5000 ;
        RECT 1002.9200 414.9000 1004.5200 415.3800 ;
        RECT 1002.9200 410.5600 1004.5200 411.0400 ;
        RECT 1002.9200 420.3400 1004.5200 420.8200 ;
        RECT 1002.9200 425.7800 1004.5200 426.2600 ;
        RECT 1002.9200 431.2200 1004.5200 431.7000 ;
        RECT 1002.9200 436.6600 1004.5200 437.1400 ;
        RECT 1285.9400 34.1000 1287.6800 34.5800 ;
        RECT 1285.9400 28.6600 1287.6800 29.1400 ;
        RECT 1285.9400 23.2200 1287.6800 23.7000 ;
        RECT 1285.9400 39.5400 1287.6800 40.0200 ;
        RECT 1285.9400 44.9800 1287.6800 45.4600 ;
        RECT 1285.9400 50.4200 1287.6800 50.9000 ;
        RECT 1285.9400 55.8600 1287.6800 56.3400 ;
        RECT 1285.9400 61.3000 1287.6800 61.7800 ;
        RECT 1285.9400 66.7400 1287.6800 67.2200 ;
        RECT 1285.9400 72.1800 1287.6800 72.6600 ;
        RECT 1285.9400 77.6200 1287.6800 78.1000 ;
        RECT 1285.9400 83.0600 1287.6800 83.5400 ;
        RECT 1285.9400 88.5000 1287.6800 88.9800 ;
        RECT 1285.9400 93.9400 1287.6800 94.4200 ;
        RECT 1285.9400 99.3800 1287.6800 99.8600 ;
        RECT 1285.9400 110.2600 1287.6800 110.7400 ;
        RECT 1285.9400 104.8200 1287.6800 105.3000 ;
        RECT 1285.9400 115.7000 1287.6800 116.1800 ;
        RECT 1285.9400 121.1400 1287.6800 121.6200 ;
        RECT 1285.9400 126.5800 1287.6800 127.0600 ;
        RECT 1285.9400 135.7400 1287.6800 137.6000 ;
        RECT 1285.9400 132.0200 1287.6800 132.5000 ;
        RECT 1285.9400 176.0000 1287.6800 177.8600 ;
        RECT 1285.9400 168.8400 1287.6800 170.7000 ;
        RECT 1293.4000 163.4400 1295.0000 163.9200 ;
        RECT 1285.9400 186.0300 1287.6800 187.8900 ;
        RECT 1506.1600 34.1000 1507.7600 34.5800 ;
        RECT 1506.1600 28.6600 1507.7600 29.1400 ;
        RECT 1506.1600 23.2200 1507.7600 23.7000 ;
        RECT 1506.1600 39.5400 1507.7600 40.0200 ;
        RECT 1506.1600 44.9800 1507.7600 45.4600 ;
        RECT 1506.1600 50.4200 1507.7600 50.9000 ;
        RECT 1506.1600 55.8600 1507.7600 56.3400 ;
        RECT 1506.1600 61.3000 1507.7600 61.7800 ;
        RECT 1506.1600 66.7400 1507.7600 67.2200 ;
        RECT 1506.1600 72.1800 1507.7600 72.6600 ;
        RECT 1506.1600 77.6200 1507.7600 78.1000 ;
        RECT 1506.1600 83.0600 1507.7600 83.5400 ;
        RECT 1506.1600 88.5000 1507.7600 88.9800 ;
        RECT 1506.1600 93.9400 1507.7600 94.4200 ;
        RECT 1506.1600 99.3800 1507.7600 99.8600 ;
        RECT 1506.1600 110.2600 1507.7600 110.7400 ;
        RECT 1506.1600 104.8200 1507.7600 105.3000 ;
        RECT 1506.1600 115.7000 1507.7600 116.1800 ;
        RECT 1506.1600 121.1400 1507.7600 121.6200 ;
        RECT 1506.1600 126.5800 1507.7600 127.0600 ;
        RECT 1506.1600 132.0200 1507.7600 132.5000 ;
        RECT 1513.6200 163.4400 1515.2200 163.9200 ;
        RECT 1293.3000 391.3800 1294.9000 391.8600 ;
        RECT 1513.5200 391.3800 1515.1200 391.8600 ;
        RECT 6.0000 447.5400 9.0000 448.0200 ;
        RECT 6.0000 452.9800 9.0000 453.4600 ;
        RECT 6.0000 458.4200 9.0000 458.9000 ;
        RECT 6.0000 463.8600 9.0000 464.3400 ;
        RECT 6.0000 469.3000 9.0000 469.7800 ;
        RECT 6.0000 474.7400 9.0000 475.2200 ;
        RECT 6.0000 480.1800 9.0000 480.6600 ;
        RECT 6.0000 485.6200 9.0000 486.1000 ;
        RECT 6.0000 491.0600 9.0000 491.5400 ;
        RECT 6.0000 496.5000 9.0000 496.9800 ;
        RECT 6.0000 501.9400 9.0000 502.4200 ;
        RECT 6.0000 507.3800 9.0000 507.8600 ;
        RECT 6.0000 512.8200 9.0000 513.3000 ;
        RECT 6.0000 518.2600 9.0000 518.7400 ;
        RECT 6.0000 523.7000 9.0000 524.1800 ;
        RECT 6.0000 529.1400 9.0000 529.6200 ;
        RECT 6.0000 534.5800 9.0000 535.0600 ;
        RECT 6.0000 540.0200 9.0000 540.5000 ;
        RECT 6.0000 545.4600 9.0000 545.9400 ;
        RECT 6.0000 599.8600 9.0000 600.3400 ;
        RECT 6.0000 550.9000 9.0000 551.3800 ;
        RECT 6.0000 556.3400 9.0000 556.8200 ;
        RECT 6.0000 561.7800 9.0000 562.2600 ;
        RECT 6.0000 567.2200 9.0000 567.7000 ;
        RECT 6.0000 572.6600 9.0000 573.1400 ;
        RECT 6.0000 578.1000 9.0000 578.5800 ;
        RECT 6.0000 583.5400 9.0000 584.0200 ;
        RECT 6.0000 588.9800 9.0000 589.4600 ;
        RECT 6.0000 594.4200 9.0000 594.9000 ;
        RECT 6.0000 605.3000 9.0000 605.7800 ;
        RECT 6.0000 610.7400 9.0000 611.2200 ;
        RECT 6.0000 616.1800 9.0000 616.6600 ;
        RECT 6.0000 621.6200 9.0000 622.1000 ;
        RECT 6.0000 627.0600 9.0000 627.5400 ;
        RECT 6.0000 632.5000 9.0000 632.9800 ;
        RECT 6.0000 635.5400 9.0000 637.5700 ;
        RECT 6.0000 643.3800 9.0000 643.8600 ;
        RECT 6.0000 648.8200 9.0000 649.3000 ;
        RECT 152.9200 643.3800 154.5200 643.8600 ;
        RECT 152.9200 648.8200 154.5200 649.3000 ;
        RECT 6.0000 654.2600 9.0000 654.7400 ;
        RECT 6.0000 659.7000 9.0000 660.1800 ;
        RECT 6.0000 665.1400 9.0000 665.6200 ;
        RECT 6.0000 670.5800 9.0000 671.0600 ;
        RECT 6.0000 676.0200 9.0000 676.5000 ;
        RECT 6.0000 692.3400 9.0000 692.8200 ;
        RECT 6.0000 681.4600 9.0000 681.9400 ;
        RECT 6.0000 686.9000 9.0000 687.3800 ;
        RECT 6.0000 697.7800 9.0000 698.2600 ;
        RECT 6.0000 703.2200 9.0000 703.7000 ;
        RECT 6.0000 708.6600 9.0000 709.1400 ;
        RECT 6.0000 714.1000 9.0000 714.5800 ;
        RECT 6.0000 719.5400 9.0000 720.0200 ;
        RECT 6.0000 724.9800 9.0000 725.4600 ;
        RECT 6.0000 730.4200 9.0000 730.9000 ;
        RECT 6.0000 735.8600 9.0000 736.3400 ;
        RECT 6.0000 741.3000 9.0000 741.7800 ;
        RECT 6.0000 746.7400 9.0000 747.2200 ;
        RECT 6.0000 752.1800 9.0000 752.6600 ;
        RECT 6.0000 757.6200 9.0000 758.1000 ;
        RECT 152.9200 654.2600 154.5200 654.7400 ;
        RECT 152.9200 659.7000 154.5200 660.1800 ;
        RECT 152.9200 665.1400 154.5200 665.6200 ;
        RECT 152.9200 670.5800 154.5200 671.0600 ;
        RECT 152.9200 676.0200 154.5200 676.5000 ;
        RECT 152.9200 692.3400 154.5200 692.8200 ;
        RECT 152.9200 686.9000 154.5200 687.3800 ;
        RECT 152.9200 681.4600 154.5200 681.9400 ;
        RECT 152.9200 697.7800 154.5200 698.2600 ;
        RECT 152.9200 703.2200 154.5200 703.7000 ;
        RECT 152.9200 708.6600 154.5200 709.1400 ;
        RECT 152.9200 714.1000 154.5200 714.5800 ;
        RECT 152.9200 719.5400 154.5200 720.0200 ;
        RECT 152.9200 724.9800 154.5200 725.4600 ;
        RECT 152.9200 730.4200 154.5200 730.9000 ;
        RECT 152.9200 735.8600 154.5200 736.3400 ;
        RECT 152.9200 741.3000 154.5200 741.7800 ;
        RECT 152.9200 746.7400 154.5200 747.2200 ;
        RECT 152.9200 752.1800 154.5200 752.6600 ;
        RECT 152.9200 757.6200 154.5200 758.1000 ;
        RECT 6.0000 763.0600 9.0000 763.5400 ;
        RECT 6.0000 768.5000 9.0000 768.9800 ;
        RECT 6.0000 773.9400 9.0000 774.4200 ;
        RECT 6.0000 779.3800 9.0000 779.8600 ;
        RECT 6.0000 784.8200 9.0000 785.3000 ;
        RECT 6.0000 790.2600 9.0000 790.7400 ;
        RECT 6.0000 795.7000 9.0000 796.1800 ;
        RECT 6.0000 801.1400 9.0000 801.6200 ;
        RECT 6.0000 806.5800 9.0000 807.0600 ;
        RECT 6.0000 812.0200 9.0000 812.5000 ;
        RECT 6.0000 817.4600 9.0000 817.9400 ;
        RECT 6.0000 822.9000 9.0000 823.3800 ;
        RECT 6.0000 828.3400 9.0000 828.8200 ;
        RECT 6.0000 833.7800 9.0000 834.2600 ;
        RECT 6.0000 850.1000 9.0000 850.5800 ;
        RECT 6.0000 839.2200 9.0000 839.7000 ;
        RECT 6.0000 844.6600 9.0000 845.1400 ;
        RECT 6.0000 855.5400 9.0000 856.0200 ;
        RECT 6.0000 860.9800 9.0000 861.4600 ;
        RECT 152.9200 763.0600 154.5200 763.5400 ;
        RECT 152.9200 768.5000 154.5200 768.9800 ;
        RECT 152.9200 773.9400 154.5200 774.4200 ;
        RECT 152.9200 779.3800 154.5200 779.8600 ;
        RECT 152.9200 784.8200 154.5200 785.3000 ;
        RECT 152.9200 790.2600 154.5200 790.7400 ;
        RECT 152.9200 795.7000 154.5200 796.1800 ;
        RECT 152.9200 801.1400 154.5200 801.6200 ;
        RECT 152.9200 806.5800 154.5200 807.0600 ;
        RECT 152.9200 812.0200 154.5200 812.5000 ;
        RECT 152.9200 817.4600 154.5200 817.9400 ;
        RECT 152.9200 822.9000 154.5200 823.3800 ;
        RECT 152.9200 828.3400 154.5200 828.8200 ;
        RECT 152.9200 833.7800 154.5200 834.2600 ;
        RECT 152.9200 850.1000 154.5200 850.5800 ;
        RECT 152.9200 839.2200 154.5200 839.7000 ;
        RECT 152.9200 844.6600 154.5200 845.1400 ;
        RECT 152.9200 855.5400 154.5200 856.0200 ;
        RECT 152.9200 860.9800 154.5200 861.4600 ;
        RECT 502.9200 447.5400 504.5200 448.0200 ;
        RECT 502.9200 452.9800 504.5200 453.4600 ;
        RECT 502.9200 458.4200 504.5200 458.9000 ;
        RECT 502.9200 463.8600 504.5200 464.3400 ;
        RECT 502.9200 469.3000 504.5200 469.7800 ;
        RECT 502.9200 474.7400 504.5200 475.2200 ;
        RECT 502.9200 480.1800 504.5200 480.6600 ;
        RECT 502.9200 485.6200 504.5200 486.1000 ;
        RECT 502.9200 491.0600 504.5200 491.5400 ;
        RECT 502.9200 496.5000 504.5200 496.9800 ;
        RECT 502.9200 501.9400 504.5200 502.4200 ;
        RECT 502.9200 507.3800 504.5200 507.8600 ;
        RECT 502.9200 512.8200 504.5200 513.3000 ;
        RECT 502.9200 518.2600 504.5200 518.7400 ;
        RECT 502.9200 523.7000 504.5200 524.1800 ;
        RECT 502.9200 529.1400 504.5200 529.6200 ;
        RECT 502.9200 534.5800 504.5200 535.0600 ;
        RECT 502.9200 540.0200 504.5200 540.5000 ;
        RECT 502.9200 545.4600 504.5200 545.9400 ;
        RECT 502.9200 599.8600 504.5200 600.3400 ;
        RECT 502.9200 550.9000 504.5200 551.3800 ;
        RECT 502.9200 556.3400 504.5200 556.8200 ;
        RECT 502.9200 561.7800 504.5200 562.2600 ;
        RECT 502.9200 567.2200 504.5200 567.7000 ;
        RECT 502.9200 572.6600 504.5200 573.1400 ;
        RECT 502.9200 583.5400 504.5200 584.0200 ;
        RECT 502.9200 578.1000 504.5200 578.5800 ;
        RECT 502.9200 588.9800 504.5200 589.4600 ;
        RECT 502.9200 594.4200 504.5200 594.9000 ;
        RECT 502.9200 610.7400 504.5200 611.2200 ;
        RECT 502.9200 605.3000 504.5200 605.7800 ;
        RECT 502.9200 616.1800 504.5200 616.6600 ;
        RECT 502.9200 621.6200 504.5200 622.1000 ;
        RECT 502.9200 627.0600 504.5200 627.5400 ;
        RECT 502.9200 632.5000 504.5200 632.9800 ;
        RECT 665.7200 447.5400 667.3200 448.0200 ;
        RECT 665.7200 452.9800 667.3200 453.4600 ;
        RECT 665.7200 463.8600 667.3200 464.3400 ;
        RECT 665.7200 458.4200 667.3200 458.9000 ;
        RECT 665.7200 469.3000 667.3200 469.7800 ;
        RECT 665.7200 474.7400 667.3200 475.2200 ;
        RECT 665.7200 480.1800 667.3200 480.6600 ;
        RECT 665.7200 485.6200 667.3200 486.1000 ;
        RECT 665.7200 491.0600 667.3200 491.5400 ;
        RECT 665.7200 507.3800 667.3200 507.8600 ;
        RECT 665.7200 501.9400 667.3200 502.4200 ;
        RECT 665.7200 496.5000 667.3200 496.9800 ;
        RECT 665.7200 512.8200 667.3200 513.3000 ;
        RECT 665.7200 518.2600 667.3200 518.7400 ;
        RECT 665.7200 523.7000 667.3200 524.1800 ;
        RECT 665.7200 529.1400 667.3200 529.6200 ;
        RECT 665.7200 534.5800 667.3200 535.0600 ;
        RECT 665.7200 540.0200 667.3200 540.5000 ;
        RECT 665.7200 545.4600 667.3200 545.9400 ;
        RECT 665.7200 599.8600 667.3200 600.3400 ;
        RECT 665.7200 550.9000 667.3200 551.3800 ;
        RECT 665.7200 556.3400 667.3200 556.8200 ;
        RECT 665.7200 561.7800 667.3200 562.2600 ;
        RECT 665.7200 567.2200 667.3200 567.7000 ;
        RECT 665.7200 572.6600 667.3200 573.1400 ;
        RECT 665.7200 583.5400 667.3200 584.0200 ;
        RECT 665.7200 578.1000 667.3200 578.5800 ;
        RECT 665.7200 588.9800 667.3200 589.4600 ;
        RECT 665.7200 594.4200 667.3200 594.9000 ;
        RECT 665.7200 610.7400 667.3200 611.2200 ;
        RECT 665.7200 605.3000 667.3200 605.7800 ;
        RECT 665.7200 616.1800 667.3200 616.6600 ;
        RECT 665.7200 621.6200 667.3200 622.1000 ;
        RECT 665.7200 627.0600 667.3200 627.5400 ;
        RECT 665.7200 632.5000 667.3200 632.9800 ;
        RECT 6.0000 871.8600 9.0000 872.3400 ;
        RECT 6.0000 865.1800 9.0000 866.9000 ;
        RECT 6.0000 877.3000 9.0000 877.7800 ;
        RECT 6.0000 882.7400 9.0000 883.2200 ;
        RECT 6.0000 888.1800 9.0000 888.6600 ;
        RECT 6.0000 893.6200 9.0000 894.1000 ;
        RECT 6.0000 899.0600 9.0000 899.5400 ;
        RECT 6.0000 904.5000 9.0000 904.9800 ;
        RECT 6.0000 909.9400 9.0000 910.4200 ;
        RECT 6.0000 915.3800 9.0000 915.8600 ;
        RECT 6.0000 920.8200 9.0000 921.3000 ;
        RECT 6.0000 926.2600 9.0000 926.7400 ;
        RECT 6.0000 931.7000 9.0000 932.1800 ;
        RECT 6.0000 937.1400 9.0000 937.6200 ;
        RECT 6.0000 942.5800 9.0000 943.0600 ;
        RECT 6.0000 948.0200 9.0000 948.5000 ;
        RECT 6.0000 953.4600 9.0000 953.9400 ;
        RECT 6.0000 958.9000 9.0000 959.3800 ;
        RECT 6.0000 964.3400 9.0000 964.8200 ;
        RECT 152.9200 871.8600 154.5200 872.3400 ;
        RECT 152.9200 865.1800 154.5200 866.9000 ;
        RECT 152.9200 877.3000 154.5200 877.7800 ;
        RECT 152.9200 882.7400 154.5200 883.2200 ;
        RECT 152.9200 888.1800 154.5200 888.6600 ;
        RECT 152.9200 893.6200 154.5200 894.1000 ;
        RECT 152.9200 899.0600 154.5200 899.5400 ;
        RECT 152.9200 904.5000 154.5200 904.9800 ;
        RECT 152.9200 909.9400 154.5200 910.4200 ;
        RECT 152.9200 915.3800 154.5200 915.8600 ;
        RECT 152.9200 920.8200 154.5200 921.3000 ;
        RECT 152.9200 926.2600 154.5200 926.7400 ;
        RECT 152.9200 931.7000 154.5200 932.1800 ;
        RECT 152.9200 937.1400 154.5200 937.6200 ;
        RECT 152.9200 942.5800 154.5200 943.0600 ;
        RECT 152.9200 948.0200 154.5200 948.5000 ;
        RECT 152.9200 953.4600 154.5200 953.9400 ;
        RECT 152.9200 958.9000 154.5200 959.3800 ;
        RECT 152.9200 964.3400 154.5200 964.8200 ;
        RECT 6.0000 969.7800 9.0000 970.2600 ;
        RECT 6.0000 975.2200 9.0000 975.7000 ;
        RECT 6.0000 980.6600 9.0000 981.1400 ;
        RECT 6.0000 986.1000 9.0000 986.5800 ;
        RECT 6.0000 991.5400 9.0000 992.0200 ;
        RECT 6.0000 996.9800 9.0000 997.4600 ;
        RECT 6.0000 1002.4200 9.0000 1002.9000 ;
        RECT 6.0000 1007.8600 9.0000 1008.3400 ;
        RECT 6.0000 1013.3000 9.0000 1013.7800 ;
        RECT 6.0000 1018.7400 9.0000 1019.2200 ;
        RECT 6.0000 1024.1800 9.0000 1024.6600 ;
        RECT 6.0000 1029.6200 9.0000 1030.1000 ;
        RECT 6.0000 1035.0600 9.0000 1035.5400 ;
        RECT 6.0000 1040.5000 9.0000 1040.9800 ;
        RECT 6.0000 1045.9400 9.0000 1046.4200 ;
        RECT 6.0000 1051.3800 9.0000 1051.8600 ;
        RECT 6.0000 1056.8200 9.0000 1057.3000 ;
        RECT 6.0000 1062.2600 9.0000 1062.7400 ;
        RECT 6.0000 1067.7000 9.0000 1068.1800 ;
        RECT 6.0000 1073.1400 9.0000 1073.6200 ;
        RECT 152.9200 969.7800 154.5200 970.2600 ;
        RECT 152.9200 975.2200 154.5200 975.7000 ;
        RECT 152.9200 980.6600 154.5200 981.1400 ;
        RECT 152.9200 986.1000 154.5200 986.5800 ;
        RECT 152.9200 991.5400 154.5200 992.0200 ;
        RECT 152.9200 996.9800 154.5200 997.4600 ;
        RECT 152.9200 1002.4200 154.5200 1002.9000 ;
        RECT 152.9200 1007.8600 154.5200 1008.3400 ;
        RECT 152.9200 1013.3000 154.5200 1013.7800 ;
        RECT 152.9200 1018.7400 154.5200 1019.2200 ;
        RECT 152.9200 1024.1800 154.5200 1024.6600 ;
        RECT 152.9200 1029.6200 154.5200 1030.1000 ;
        RECT 152.9200 1035.0600 154.5200 1035.5400 ;
        RECT 152.9200 1040.5000 154.5200 1040.9800 ;
        RECT 152.9200 1045.9400 154.5200 1046.4200 ;
        RECT 152.9200 1051.3800 154.5200 1051.8600 ;
        RECT 152.9200 1056.8200 154.5200 1057.3000 ;
        RECT 152.9200 1062.2600 154.5200 1062.7400 ;
        RECT 152.9200 1067.7000 154.5200 1068.1800 ;
        RECT 152.9200 1073.1400 154.5200 1073.6200 ;
        RECT 6.0000 1100.3400 9.0000 1100.8200 ;
        RECT 6.0000 1078.5800 9.0000 1079.0600 ;
        RECT 6.0000 1084.0200 9.0000 1084.5000 ;
        RECT 6.0000 1089.4600 9.0000 1089.9400 ;
        RECT 6.0000 1105.7800 9.0000 1106.2600 ;
        RECT 6.0000 1111.2200 9.0000 1111.7000 ;
        RECT 6.0000 1116.6600 9.0000 1117.1400 ;
        RECT 6.0000 1122.1000 9.0000 1122.5800 ;
        RECT 6.0000 1127.5400 9.0000 1128.0200 ;
        RECT 6.0000 1132.9800 9.0000 1133.4600 ;
        RECT 6.0000 1138.4200 9.0000 1138.9000 ;
        RECT 6.0000 1143.8600 9.0000 1144.3400 ;
        RECT 6.0000 1149.3000 9.0000 1149.7800 ;
        RECT 6.0000 1154.7400 9.0000 1155.2200 ;
        RECT 6.0000 1160.1800 9.0000 1160.6600 ;
        RECT 6.0000 1165.6200 9.0000 1166.1000 ;
        RECT 6.0000 1171.0600 9.0000 1171.5400 ;
        RECT 6.0000 1176.5000 9.0000 1176.9800 ;
        RECT 152.9200 1100.3400 154.5200 1100.8200 ;
        RECT 152.9200 1078.5800 154.5200 1079.0600 ;
        RECT 152.9200 1084.0200 154.5200 1084.5000 ;
        RECT 152.9200 1089.4600 154.5200 1089.9400 ;
        RECT 152.9200 1105.7800 154.5200 1106.2600 ;
        RECT 152.9200 1111.2200 154.5200 1111.7000 ;
        RECT 152.9200 1116.6600 154.5200 1117.1400 ;
        RECT 152.9200 1122.1000 154.5200 1122.5800 ;
        RECT 152.9200 1127.5400 154.5200 1128.0200 ;
        RECT 152.9200 1132.9800 154.5200 1133.4600 ;
        RECT 152.9200 1138.4200 154.5200 1138.9000 ;
        RECT 152.9200 1143.8600 154.5200 1144.3400 ;
        RECT 152.9200 1149.3000 154.5200 1149.7800 ;
        RECT 152.9200 1154.7400 154.5200 1155.2200 ;
        RECT 152.9200 1160.1800 154.5200 1160.6600 ;
        RECT 152.9200 1165.6200 154.5200 1166.1000 ;
        RECT 152.9200 1171.0600 154.5200 1171.5400 ;
        RECT 152.9200 1176.5000 154.5200 1176.9800 ;
        RECT 6.0000 1181.9400 9.0000 1182.4200 ;
        RECT 6.0000 1187.3800 9.0000 1187.8600 ;
        RECT 6.0000 1192.8200 9.0000 1193.3000 ;
        RECT 6.0000 1198.2600 9.0000 1198.7400 ;
        RECT 6.0000 1203.7000 9.0000 1204.1800 ;
        RECT 6.0000 1209.1400 9.0000 1209.6200 ;
        RECT 6.0000 1214.5800 9.0000 1215.0600 ;
        RECT 6.0000 1220.0200 9.0000 1220.5000 ;
        RECT 6.0000 1225.4600 9.0000 1225.9400 ;
        RECT 6.0000 1230.9000 9.0000 1231.3800 ;
        RECT 6.0000 1258.1000 9.0000 1258.5800 ;
        RECT 6.0000 1236.3400 9.0000 1236.8200 ;
        RECT 6.0000 1241.7800 9.0000 1242.2600 ;
        RECT 6.0000 1247.2200 9.0000 1247.7000 ;
        RECT 6.0000 1252.6600 9.0000 1253.1400 ;
        RECT 6.0000 1263.5400 9.0000 1264.0200 ;
        RECT 6.0000 1268.9800 9.0000 1269.4600 ;
        RECT 6.0000 1274.4200 9.0000 1274.9000 ;
        RECT 6.0000 1279.8600 9.0000 1280.3400 ;
        RECT 152.9200 1181.9400 154.5200 1182.4200 ;
        RECT 152.9200 1187.3800 154.5200 1187.8600 ;
        RECT 152.9200 1192.8200 154.5200 1193.3000 ;
        RECT 152.9200 1198.2600 154.5200 1198.7400 ;
        RECT 152.9200 1203.7000 154.5200 1204.1800 ;
        RECT 152.9200 1209.1400 154.5200 1209.6200 ;
        RECT 152.9200 1214.5800 154.5200 1215.0600 ;
        RECT 152.9200 1220.0200 154.5200 1220.5000 ;
        RECT 152.9200 1225.4600 154.5200 1225.9400 ;
        RECT 152.9200 1230.9000 154.5200 1231.3800 ;
        RECT 152.9200 1258.1000 154.5200 1258.5800 ;
        RECT 152.9200 1236.3400 154.5200 1236.8200 ;
        RECT 152.9200 1241.7800 154.5200 1242.2600 ;
        RECT 152.9200 1247.2200 154.5200 1247.7000 ;
        RECT 152.9200 1252.6600 154.5200 1253.1400 ;
        RECT 152.9200 1263.5400 154.5200 1264.0200 ;
        RECT 152.9200 1268.9800 154.5200 1269.4600 ;
        RECT 152.9200 1274.4200 154.5200 1274.9000 ;
        RECT 152.9200 1279.8600 154.5200 1280.3400 ;
        RECT 1002.9200 452.9800 1004.5200 453.4600 ;
        RECT 1002.9200 447.5400 1004.5200 448.0200 ;
        RECT 1002.9200 458.4200 1004.5200 458.9000 ;
        RECT 1002.9200 463.8600 1004.5200 464.3400 ;
        RECT 1002.9200 469.3000 1004.5200 469.7800 ;
        RECT 1002.9200 474.7400 1004.5200 475.2200 ;
        RECT 1002.9200 480.1800 1004.5200 480.6600 ;
        RECT 1002.9200 485.6200 1004.5200 486.1000 ;
        RECT 1002.9200 491.0600 1004.5200 491.5400 ;
        RECT 1002.9200 501.9400 1004.5200 502.4200 ;
        RECT 1002.9200 496.5000 1004.5200 496.9800 ;
        RECT 1002.9200 507.3800 1004.5200 507.8600 ;
        RECT 1002.9200 512.8200 1004.5200 513.3000 ;
        RECT 1002.9200 518.2600 1004.5200 518.7400 ;
        RECT 1002.9200 529.1400 1004.5200 529.6200 ;
        RECT 1002.9200 523.7000 1004.5200 524.1800 ;
        RECT 1002.9200 534.5800 1004.5200 535.0600 ;
        RECT 1002.9200 540.0200 1004.5200 540.5000 ;
        RECT 1002.9200 545.4600 1004.5200 545.9400 ;
        RECT 1002.9200 599.8600 1004.5200 600.3400 ;
        RECT 1002.9200 550.9000 1004.5200 551.3800 ;
        RECT 1002.9200 556.3400 1004.5200 556.8200 ;
        RECT 1002.9200 561.7800 1004.5200 562.2600 ;
        RECT 1002.9200 567.2200 1004.5200 567.7000 ;
        RECT 1002.9200 572.6600 1004.5200 573.1400 ;
        RECT 1002.9200 583.5400 1004.5200 584.0200 ;
        RECT 1002.9200 578.1000 1004.5200 578.5800 ;
        RECT 1002.9200 588.9800 1004.5200 589.4600 ;
        RECT 1002.9200 594.4200 1004.5200 594.9000 ;
        RECT 965.7200 643.3800 967.3200 643.8600 ;
        RECT 965.7200 648.8200 967.3200 649.3000 ;
        RECT 1002.9200 610.7400 1004.5200 611.2200 ;
        RECT 1002.9200 605.3000 1004.5200 605.7800 ;
        RECT 1002.9200 616.1800 1004.5200 616.6600 ;
        RECT 1002.9200 621.6200 1004.5200 622.1000 ;
        RECT 1002.9200 635.5400 1004.5200 637.5700 ;
        RECT 1002.9200 632.5000 1004.5200 632.9800 ;
        RECT 1002.9200 627.0600 1004.5200 629.1300 ;
        RECT 1002.9200 643.3800 1004.5200 643.8600 ;
        RECT 1002.9200 648.8200 1004.5200 649.3000 ;
        RECT 1055.6000 621.2800 1057.2000 621.7600 ;
        RECT 1073.2200 620.1200 1074.8200 620.6000 ;
        RECT 1060.5600 627.5300 1062.1600 629.1300 ;
        RECT 1065.8600 645.5700 1067.4600 647.2700 ;
        RECT 965.7200 654.2600 967.3200 654.7400 ;
        RECT 965.7200 659.7000 967.3200 660.1800 ;
        RECT 965.7200 665.1400 967.3200 665.6200 ;
        RECT 965.7200 670.5800 967.3200 671.0600 ;
        RECT 965.7200 676.0200 967.3200 676.5000 ;
        RECT 965.7200 692.3400 967.3200 692.8200 ;
        RECT 965.7200 686.9000 967.3200 687.3800 ;
        RECT 965.7200 681.4600 967.3200 681.9400 ;
        RECT 965.7200 697.7800 967.3200 698.2600 ;
        RECT 965.7200 703.2200 967.3200 703.7000 ;
        RECT 1002.9200 654.2600 1004.5200 654.7400 ;
        RECT 1002.9200 659.7000 1004.5200 660.1800 ;
        RECT 1002.9200 665.1400 1004.5200 665.6200 ;
        RECT 1002.9200 670.5800 1004.5200 671.0600 ;
        RECT 1002.9200 676.0200 1004.5200 676.5000 ;
        RECT 1002.9200 692.3400 1004.5200 692.8200 ;
        RECT 1002.9200 686.9000 1004.5200 687.3800 ;
        RECT 1002.9200 681.4600 1004.5200 681.9400 ;
        RECT 1002.9200 697.7800 1004.5200 698.2600 ;
        RECT 1002.9200 703.2200 1004.5200 703.7000 ;
        RECT 965.7200 708.6600 967.3200 709.1400 ;
        RECT 965.7200 714.1000 967.3200 714.5800 ;
        RECT 965.7200 719.5400 967.3200 720.0200 ;
        RECT 965.7200 724.9800 967.3200 725.4600 ;
        RECT 965.7200 730.4200 967.3200 730.9000 ;
        RECT 965.7200 735.8600 967.3200 736.3400 ;
        RECT 965.7200 741.3000 967.3200 741.7800 ;
        RECT 965.7200 746.7400 967.3200 747.2200 ;
        RECT 1002.9200 708.6600 1004.5200 709.1400 ;
        RECT 1002.9200 714.1000 1004.5200 714.5800 ;
        RECT 1002.9200 719.5400 1004.5200 720.0200 ;
        RECT 1002.9200 724.9800 1004.5200 725.4600 ;
        RECT 1002.9200 730.4200 1004.5200 730.9000 ;
        RECT 1002.9200 735.8600 1004.5200 736.3400 ;
        RECT 1002.9200 741.3000 1004.5200 741.7800 ;
        RECT 1002.9200 746.7400 1004.5200 747.2200 ;
        RECT 1013.1800 850.9200 1014.7800 851.4000 ;
        RECT 1293.3000 621.0200 1294.9000 621.5000 ;
        RECT 1285.9400 635.2800 1287.6800 637.1400 ;
        RECT 1285.9400 627.3700 1287.6800 630.2800 ;
        RECT 1285.9400 645.3100 1287.6800 647.1700 ;
        RECT 1513.5200 621.0200 1515.1200 621.5000 ;
        RECT 1293.3000 850.6600 1294.9000 851.1400 ;
        RECT 1513.5200 850.6600 1515.1200 851.1400 ;
        RECT 1073.2200 1079.4000 1074.8200 1079.8800 ;
        RECT 1055.6000 1080.5600 1057.2000 1081.0400 ;
        RECT 1060.5600 1086.8100 1062.1600 1088.4100 ;
        RECT 1065.8600 1104.8500 1067.4600 1106.5500 ;
        RECT 1285.9400 1094.5600 1287.6800 1096.4200 ;
        RECT 1285.9400 1086.6500 1287.6800 1089.5600 ;
        RECT 1293.3000 1080.3000 1294.9000 1080.7800 ;
        RECT 1285.9400 1104.5900 1287.6800 1106.4500 ;
        RECT 1513.5200 1080.3000 1515.1200 1080.7800 ;
        RECT 3361.4200 442.1000 3364.4200 442.5800 ;
        RECT 2447.1800 442.1000 2448.7800 442.5800 ;
        RECT 2492.9200 442.1000 2494.5200 442.5800 ;
        RECT 3305.7200 442.1000 3307.3200 442.5800 ;
        RECT 1726.3800 12.3400 1727.9800 12.8200 ;
        RECT 1726.3800 17.7800 1727.9800 18.2600 ;
        RECT 1946.6000 12.3400 1948.2000 12.8200 ;
        RECT 1946.6000 17.7800 1948.2000 18.2600 ;
        RECT 2166.8200 12.3400 2168.4200 12.8200 ;
        RECT 2166.8200 17.7800 2168.4200 18.2600 ;
        RECT 2387.0400 12.3400 2388.6400 12.8200 ;
        RECT 2387.0400 17.7800 2388.6400 18.2600 ;
        RECT 2447.1800 12.3400 2448.7800 12.8200 ;
        RECT 2447.1800 17.7800 2448.7800 18.2600 ;
        RECT 2492.9200 12.3400 2494.5200 12.8200 ;
        RECT 2492.9200 17.7800 2494.5200 18.2600 ;
        RECT 1726.3800 34.1000 1727.9800 34.5800 ;
        RECT 1726.3800 28.6600 1727.9800 29.1400 ;
        RECT 1726.3800 23.2200 1727.9800 23.7000 ;
        RECT 1726.3800 39.5400 1727.9800 40.0200 ;
        RECT 1726.3800 44.9800 1727.9800 45.4600 ;
        RECT 1726.3800 50.4200 1727.9800 50.9000 ;
        RECT 1726.3800 55.8600 1727.9800 56.3400 ;
        RECT 1726.3800 61.3000 1727.9800 61.7800 ;
        RECT 1726.3800 66.7400 1727.9800 67.2200 ;
        RECT 1726.3800 72.1800 1727.9800 72.6600 ;
        RECT 1726.3800 77.6200 1727.9800 78.1000 ;
        RECT 1726.3800 83.0600 1727.9800 83.5400 ;
        RECT 1726.3800 88.5000 1727.9800 88.9800 ;
        RECT 1726.3800 93.9400 1727.9800 94.4200 ;
        RECT 1726.3800 99.3800 1727.9800 99.8600 ;
        RECT 1726.3800 110.2600 1727.9800 110.7400 ;
        RECT 1726.3800 104.8200 1727.9800 105.3000 ;
        RECT 1726.3800 115.7000 1727.9800 116.1800 ;
        RECT 1726.3800 121.1400 1727.9800 121.6200 ;
        RECT 1726.3800 126.5800 1727.9800 127.0600 ;
        RECT 1726.3800 132.0200 1727.9800 132.5000 ;
        RECT 1733.8400 163.4400 1735.4400 163.9200 ;
        RECT 1946.6000 34.1000 1948.2000 34.5800 ;
        RECT 1946.6000 28.6600 1948.2000 29.1400 ;
        RECT 1946.6000 23.2200 1948.2000 23.7000 ;
        RECT 1946.6000 39.5400 1948.2000 40.0200 ;
        RECT 1946.6000 44.9800 1948.2000 45.4600 ;
        RECT 1946.6000 50.4200 1948.2000 50.9000 ;
        RECT 1946.6000 55.8600 1948.2000 56.3400 ;
        RECT 1946.6000 61.3000 1948.2000 61.7800 ;
        RECT 1946.6000 66.7400 1948.2000 67.2200 ;
        RECT 1946.6000 72.1800 1948.2000 72.6600 ;
        RECT 1946.6000 77.6200 1948.2000 78.1000 ;
        RECT 1946.6000 83.0600 1948.2000 83.5400 ;
        RECT 1946.6000 88.5000 1948.2000 88.9800 ;
        RECT 1946.6000 93.9400 1948.2000 94.4200 ;
        RECT 1946.6000 99.3800 1948.2000 99.8600 ;
        RECT 1946.6000 110.2600 1948.2000 110.7400 ;
        RECT 1946.6000 104.8200 1948.2000 105.3000 ;
        RECT 1946.6000 115.7000 1948.2000 116.1800 ;
        RECT 1946.6000 121.1400 1948.2000 121.6200 ;
        RECT 1946.6000 126.5800 1948.2000 127.0600 ;
        RECT 1946.6000 132.0200 1948.2000 132.5000 ;
        RECT 1954.0600 163.4400 1955.6600 163.9200 ;
        RECT 1733.7400 391.3800 1735.3400 391.8600 ;
        RECT 2166.8200 34.1000 2168.4200 34.5800 ;
        RECT 2166.8200 28.6600 2168.4200 29.1400 ;
        RECT 2166.8200 23.2200 2168.4200 23.7000 ;
        RECT 2166.8200 39.5400 2168.4200 40.0200 ;
        RECT 2166.8200 44.9800 2168.4200 45.4600 ;
        RECT 2166.8200 50.4200 2168.4200 50.9000 ;
        RECT 2166.8200 55.8600 2168.4200 56.3400 ;
        RECT 2166.8200 61.3000 2168.4200 61.7800 ;
        RECT 2166.8200 66.7400 2168.4200 67.2200 ;
        RECT 2166.8200 72.1800 2168.4200 72.6600 ;
        RECT 2166.8200 77.6200 2168.4200 78.1000 ;
        RECT 2166.8200 83.0600 2168.4200 83.5400 ;
        RECT 2166.8200 88.5000 2168.4200 88.9800 ;
        RECT 2166.8200 93.9400 2168.4200 94.4200 ;
        RECT 2166.8200 99.3800 2168.4200 99.8600 ;
        RECT 2166.8200 110.2600 2168.4200 110.7400 ;
        RECT 2166.8200 104.8200 2168.4200 105.3000 ;
        RECT 2166.8200 115.7000 2168.4200 116.1800 ;
        RECT 2166.8200 121.1400 2168.4200 121.6200 ;
        RECT 2166.8200 126.5800 2168.4200 127.0600 ;
        RECT 2166.8200 132.0200 2168.4200 132.5000 ;
        RECT 2174.2800 163.4400 2175.8800 163.9200 ;
        RECT 2387.0400 34.1000 2388.6400 34.5800 ;
        RECT 2387.0400 28.6600 2388.6400 29.1400 ;
        RECT 2387.0400 23.2200 2388.6400 23.7000 ;
        RECT 2387.0400 39.5400 2388.6400 40.0200 ;
        RECT 2387.0400 44.9800 2388.6400 45.4600 ;
        RECT 2387.0400 50.4200 2388.6400 50.9000 ;
        RECT 2387.0400 55.8600 2388.6400 56.3400 ;
        RECT 2387.0400 61.3000 2388.6400 61.7800 ;
        RECT 2387.0400 66.7400 2388.6400 67.2200 ;
        RECT 2387.0400 72.1800 2388.6400 72.6600 ;
        RECT 2387.0400 77.6200 2388.6400 78.1000 ;
        RECT 2387.0400 83.0600 2388.6400 83.5400 ;
        RECT 2387.0400 88.5000 2388.6400 88.9800 ;
        RECT 2387.0400 93.9400 2388.6400 94.4200 ;
        RECT 2387.0400 99.3800 2388.6400 99.8600 ;
        RECT 2387.0400 110.2600 2388.6400 110.7400 ;
        RECT 2387.0400 104.8200 2388.6400 105.3000 ;
        RECT 2387.0400 115.7000 2388.6400 116.1800 ;
        RECT 2387.0400 121.1400 2388.6400 121.6200 ;
        RECT 2447.1800 34.1000 2448.7800 34.5800 ;
        RECT 2447.1800 28.6600 2448.7800 29.1400 ;
        RECT 2447.1800 23.2200 2448.7800 23.7000 ;
        RECT 2447.1800 39.5400 2448.7800 40.0200 ;
        RECT 2447.1800 44.9800 2448.7800 45.4600 ;
        RECT 2447.1800 50.4200 2448.7800 50.9000 ;
        RECT 2447.1800 55.8600 2448.7800 56.3400 ;
        RECT 2447.1800 61.3000 2448.7800 61.7800 ;
        RECT 2447.1800 66.7400 2448.7800 67.2200 ;
        RECT 2447.1800 72.1800 2448.7800 72.6600 ;
        RECT 2492.9200 34.1000 2494.5200 34.5800 ;
        RECT 2492.9200 28.6600 2494.5200 29.1400 ;
        RECT 2492.9200 23.2200 2494.5200 23.7000 ;
        RECT 2492.9200 39.5400 2494.5200 40.0200 ;
        RECT 2492.9200 44.9800 2494.5200 45.4600 ;
        RECT 2492.9200 50.4200 2494.5200 50.9000 ;
        RECT 2492.9200 55.8600 2494.5200 56.3400 ;
        RECT 2492.9200 61.3000 2494.5200 61.7800 ;
        RECT 2492.9200 66.7400 2494.5200 67.2200 ;
        RECT 2492.9200 72.1800 2494.5200 72.6600 ;
        RECT 2447.1800 77.6200 2448.7800 78.1000 ;
        RECT 2447.1800 83.0600 2448.7800 83.5400 ;
        RECT 2447.1800 88.5000 2448.7800 88.9800 ;
        RECT 2447.1800 93.9400 2448.7800 94.4200 ;
        RECT 2447.1800 99.3800 2448.7800 99.8600 ;
        RECT 2447.1800 110.2600 2448.7800 110.7400 ;
        RECT 2447.1800 104.8200 2448.7800 105.3000 ;
        RECT 2447.1800 115.7000 2448.7800 116.1800 ;
        RECT 2447.1800 121.1400 2448.7800 121.6200 ;
        RECT 2492.9200 77.6200 2494.5200 78.1000 ;
        RECT 2492.9200 83.0600 2494.5200 83.5400 ;
        RECT 2492.9200 88.5000 2494.5200 88.9800 ;
        RECT 2492.9200 93.9400 2494.5200 94.4200 ;
        RECT 2492.9200 99.3800 2494.5200 99.8600 ;
        RECT 2492.9200 110.2600 2494.5200 110.7400 ;
        RECT 2492.9200 104.8200 2494.5200 105.3000 ;
        RECT 2492.9200 115.7000 2494.5200 116.1800 ;
        RECT 2492.9200 121.1400 2494.5200 121.6200 ;
        RECT 2387.0400 126.5800 2388.6400 127.0600 ;
        RECT 2387.0400 132.0200 2388.6400 132.5000 ;
        RECT 2389.5000 137.4600 2390.0000 137.9400 ;
        RECT 2387.0400 142.9000 2388.6400 143.3800 ;
        RECT 2387.0400 148.3400 2388.6400 148.8200 ;
        RECT 2387.0400 153.7800 2388.6400 154.2600 ;
        RECT 2387.0400 159.2200 2388.6400 159.7000 ;
        RECT 2387.0400 164.6600 2388.6400 165.1400 ;
        RECT 2387.0400 168.8400 2388.6400 170.5800 ;
        RECT 2447.1800 126.5800 2448.7800 127.0600 ;
        RECT 2447.1800 132.0200 2448.7800 132.5000 ;
        RECT 2447.1800 137.4600 2448.7800 137.9400 ;
        RECT 2447.1800 142.9000 2448.7800 143.3800 ;
        RECT 2447.1800 148.3400 2448.7800 148.8200 ;
        RECT 2447.1800 153.7800 2448.7800 154.2600 ;
        RECT 2447.1800 159.2200 2448.7800 159.7000 ;
        RECT 2447.1800 164.6600 2448.7800 165.1400 ;
        RECT 2447.1800 170.1000 2448.7800 170.5800 ;
        RECT 2447.1800 175.5400 2448.7800 177.6000 ;
        RECT 2492.9200 126.5800 2494.5200 127.0600 ;
        RECT 2492.9200 132.0200 2494.5200 132.5000 ;
        RECT 2492.9200 137.4600 2494.5200 137.9400 ;
        RECT 2492.9200 142.9000 2494.5200 143.3800 ;
        RECT 2492.9200 148.3400 2494.5200 148.8200 ;
        RECT 2492.9200 153.7800 2494.5200 154.2600 ;
        RECT 2492.9200 159.2200 2494.5200 159.7000 ;
        RECT 2492.9200 164.6600 2494.5200 165.1400 ;
        RECT 2492.9200 170.1000 2494.5200 170.5800 ;
        RECT 2492.9200 175.5400 2494.5200 176.0200 ;
        RECT 2447.1800 191.8600 2448.7800 192.3400 ;
        RECT 2447.1800 180.9800 2448.7800 181.4600 ;
        RECT 2447.1800 186.4200 2448.7800 186.9000 ;
        RECT 2447.1800 197.3000 2448.7800 197.7800 ;
        RECT 2447.1800 202.7400 2448.7800 203.2200 ;
        RECT 2447.1800 208.1800 2448.7800 208.6600 ;
        RECT 2447.1800 213.6200 2448.7800 214.1000 ;
        RECT 2447.1800 219.0600 2448.7800 219.5400 ;
        RECT 2447.1800 224.5000 2448.7800 224.9800 ;
        RECT 2447.1800 229.9400 2448.7800 230.4200 ;
        RECT 2492.9200 191.8600 2494.5200 192.3400 ;
        RECT 2492.9200 186.4200 2494.5200 186.9000 ;
        RECT 2492.9200 180.9800 2494.5200 181.4600 ;
        RECT 2492.9200 197.3000 2494.5200 197.7800 ;
        RECT 2492.9200 202.7400 2494.5200 203.2200 ;
        RECT 2492.9200 208.1800 2494.5200 208.6600 ;
        RECT 2492.9200 213.6200 2494.5200 214.1000 ;
        RECT 2492.9200 219.0600 2494.5200 219.5400 ;
        RECT 2492.9200 224.5000 2494.5200 224.9800 ;
        RECT 2492.9200 229.9400 2494.5200 230.4200 ;
        RECT 2174.1800 391.3800 2175.7800 391.8600 ;
        RECT 2447.1800 235.3800 2448.7800 235.8600 ;
        RECT 2447.1800 240.8200 2448.7800 241.3000 ;
        RECT 2447.1800 246.2600 2448.7800 246.7400 ;
        RECT 2447.1800 251.7000 2448.7800 252.1800 ;
        RECT 2447.1800 257.1400 2448.7800 257.6200 ;
        RECT 2447.1800 262.5800 2448.7800 263.0600 ;
        RECT 2447.1800 268.0200 2448.7800 268.5000 ;
        RECT 2447.1800 273.4600 2448.7800 273.9400 ;
        RECT 2447.1800 278.9000 2448.7800 279.3800 ;
        RECT 2492.9200 235.3800 2494.5200 235.8600 ;
        RECT 2492.9200 240.8200 2494.5200 241.3000 ;
        RECT 2492.9200 246.2600 2494.5200 246.7400 ;
        RECT 2492.9200 251.7000 2494.5200 252.1800 ;
        RECT 2492.9200 257.1400 2494.5200 257.6200 ;
        RECT 2492.9200 268.0200 2494.5200 268.5000 ;
        RECT 2492.9200 262.5800 2494.5200 263.0600 ;
        RECT 2492.9200 273.4600 2494.5200 273.9400 ;
        RECT 2492.9200 278.9000 2494.5200 279.3800 ;
        RECT 2447.1800 284.3400 2448.7800 284.8200 ;
        RECT 2447.1800 289.7800 2448.7800 290.2600 ;
        RECT 2447.1800 295.2200 2448.7800 295.7000 ;
        RECT 2447.1800 300.6600 2448.7800 301.1400 ;
        RECT 2447.1800 306.1000 2448.7800 306.5800 ;
        RECT 2447.1800 311.5400 2448.7800 312.0200 ;
        RECT 2447.1800 316.9800 2448.7800 317.4600 ;
        RECT 2447.1800 322.4200 2448.7800 322.9000 ;
        RECT 2447.1800 327.8600 2448.7800 328.3400 ;
        RECT 2447.1800 333.3000 2448.7800 333.7800 ;
        RECT 2492.9200 284.3400 2494.5200 284.8200 ;
        RECT 2492.9200 289.7800 2494.5200 290.2600 ;
        RECT 2492.9200 295.2200 2494.5200 295.7000 ;
        RECT 2492.9200 300.6600 2494.5200 301.1400 ;
        RECT 2492.9200 306.1000 2494.5200 306.5800 ;
        RECT 2492.9200 311.5400 2494.5200 312.0200 ;
        RECT 2492.9200 316.9800 2494.5200 317.4600 ;
        RECT 2492.9200 322.4200 2494.5200 322.9000 ;
        RECT 2492.9200 327.8600 2494.5200 328.3400 ;
        RECT 2492.9200 333.3000 2494.5200 333.7800 ;
        RECT 2394.4000 391.3800 2396.0000 391.8600 ;
        RECT 2447.1800 349.6200 2448.7800 350.1000 ;
        RECT 2447.1800 338.7400 2448.7800 339.2200 ;
        RECT 2447.1800 344.1800 2448.7800 344.6600 ;
        RECT 2447.1800 355.0600 2448.7800 355.5400 ;
        RECT 2447.1800 360.5000 2448.7800 360.9800 ;
        RECT 2447.1800 365.9400 2448.7800 366.4200 ;
        RECT 2447.1800 371.3800 2448.7800 371.8600 ;
        RECT 2447.1800 376.8200 2448.7800 377.3000 ;
        RECT 2447.1800 382.2600 2448.7800 382.7400 ;
        RECT 2447.1800 387.7000 2448.7800 388.1800 ;
        RECT 2492.9200 349.6200 2494.5200 350.1000 ;
        RECT 2492.9200 344.1800 2494.5200 344.6600 ;
        RECT 2492.9200 338.7400 2494.5200 339.2200 ;
        RECT 2492.9200 355.0600 2494.5200 355.5400 ;
        RECT 2492.9200 360.5000 2494.5200 360.9800 ;
        RECT 2492.9200 371.3800 2494.5200 371.8600 ;
        RECT 2492.9200 365.9400 2494.5200 366.4200 ;
        RECT 2492.9200 376.8200 2494.5200 377.3000 ;
        RECT 2492.9200 382.2600 2494.5200 382.7400 ;
        RECT 2492.9200 387.7000 2494.5200 388.1800 ;
        RECT 2447.1800 393.1400 2448.7800 393.6200 ;
        RECT 2447.1800 404.0200 2448.7800 404.5000 ;
        RECT 2447.1800 409.4600 2448.7800 409.9400 ;
        RECT 2449.6400 414.9000 2450.1400 415.3800 ;
        RECT 2447.1800 425.7800 2448.7800 426.2600 ;
        RECT 2447.1800 420.3400 2448.7800 420.8200 ;
        RECT 2447.1800 431.2200 2448.7800 431.7000 ;
        RECT 2447.1800 436.6600 2448.7800 437.1400 ;
        RECT 2492.9200 393.1400 2494.5200 393.6200 ;
        RECT 2492.9200 398.5800 2494.5200 399.0600 ;
        RECT 2492.9200 404.0200 2494.5200 404.5000 ;
        RECT 2492.9200 409.4600 2494.5200 409.9400 ;
        RECT 2492.9200 414.9000 2494.5200 415.3800 ;
        RECT 2492.9200 425.7800 2494.5200 426.2600 ;
        RECT 2492.9200 420.3400 2494.5200 420.8200 ;
        RECT 2492.9200 431.2200 2494.5200 431.7000 ;
        RECT 2492.9200 436.6600 2494.5200 437.1400 ;
        RECT 3305.7200 12.3400 3307.3200 12.8200 ;
        RECT 3305.7200 17.7800 3307.3200 18.2600 ;
        RECT 3361.4200 17.7800 3364.4200 18.2600 ;
        RECT 3361.4200 12.3400 3364.4200 12.8200 ;
        RECT 3305.7200 34.1000 3307.3200 34.5800 ;
        RECT 3305.7200 28.6600 3307.3200 29.1400 ;
        RECT 3305.7200 23.2200 3307.3200 23.7000 ;
        RECT 3305.7200 39.5400 3307.3200 40.0200 ;
        RECT 3305.7200 44.9800 3307.3200 45.4600 ;
        RECT 3305.7200 50.4200 3307.3200 50.9000 ;
        RECT 3305.7200 55.8600 3307.3200 56.3400 ;
        RECT 3305.7200 61.3000 3307.3200 61.7800 ;
        RECT 3305.7200 66.7400 3307.3200 67.2200 ;
        RECT 3305.7200 72.1800 3307.3200 72.6600 ;
        RECT 3361.4200 34.1000 3364.4200 34.5800 ;
        RECT 3361.4200 23.2200 3364.4200 23.7000 ;
        RECT 3361.4200 28.6600 3364.4200 29.1400 ;
        RECT 3361.4200 39.5400 3364.4200 40.0200 ;
        RECT 3361.4200 44.9800 3364.4200 45.4600 ;
        RECT 3361.4200 50.4200 3364.4200 50.9000 ;
        RECT 3361.4200 55.8600 3364.4200 56.3400 ;
        RECT 3361.4200 61.3000 3364.4200 61.7800 ;
        RECT 3361.4200 66.7400 3364.4200 67.2200 ;
        RECT 3361.4200 72.1800 3364.4200 72.6600 ;
        RECT 3305.7200 77.6200 3307.3200 78.1000 ;
        RECT 3305.7200 83.0600 3307.3200 83.5400 ;
        RECT 3305.7200 88.5000 3307.3200 88.9800 ;
        RECT 3305.7200 93.9400 3307.3200 94.4200 ;
        RECT 3305.7200 99.3800 3307.3200 99.8600 ;
        RECT 3305.7200 110.2600 3307.3200 110.7400 ;
        RECT 3305.7200 104.8200 3307.3200 105.3000 ;
        RECT 3305.7200 115.7000 3307.3200 116.1800 ;
        RECT 3305.7200 121.1400 3307.3200 121.6200 ;
        RECT 3361.4200 77.6200 3364.4200 78.1000 ;
        RECT 3361.4200 83.0600 3364.4200 83.5400 ;
        RECT 3361.4200 88.5000 3364.4200 88.9800 ;
        RECT 3361.4200 93.9400 3364.4200 94.4200 ;
        RECT 3361.4200 99.3800 3364.4200 99.8600 ;
        RECT 3361.4200 104.8200 3364.4200 105.3000 ;
        RECT 3361.4200 110.2600 3364.4200 110.7400 ;
        RECT 3361.4200 115.7000 3364.4200 116.1800 ;
        RECT 3361.4200 121.1400 3364.4200 121.6200 ;
        RECT 3305.7200 126.5800 3307.3200 127.0600 ;
        RECT 3305.7200 132.0200 3307.3200 132.5000 ;
        RECT 3305.7200 137.4600 3307.3200 137.9400 ;
        RECT 3305.7200 142.9000 3307.3200 143.3800 ;
        RECT 3305.7200 148.3400 3307.3200 148.8200 ;
        RECT 3305.7200 153.7800 3307.3200 154.2600 ;
        RECT 3305.7200 159.2200 3307.3200 159.7000 ;
        RECT 3305.7200 164.6600 3307.3200 165.1400 ;
        RECT 3305.7200 170.1000 3307.3200 170.5800 ;
        RECT 3305.7200 175.5400 3307.3200 176.0200 ;
        RECT 3361.4200 126.5800 3364.4200 127.0600 ;
        RECT 3361.4200 132.0200 3364.4200 132.5000 ;
        RECT 3361.4200 137.4600 3364.4200 137.9400 ;
        RECT 3361.4200 142.9000 3364.4200 143.3800 ;
        RECT 3361.4200 148.3400 3364.4200 148.8200 ;
        RECT 3361.4200 153.7800 3364.4200 154.2600 ;
        RECT 3361.4200 159.2200 3364.4200 159.7000 ;
        RECT 3361.4200 164.6600 3364.4200 165.1400 ;
        RECT 3361.4200 170.1000 3364.4200 170.5800 ;
        RECT 3361.4200 175.5400 3364.4200 176.0200 ;
        RECT 3305.7200 191.8600 3307.3200 192.3400 ;
        RECT 3305.7200 186.4200 3307.3200 186.9000 ;
        RECT 3305.7200 180.9800 3307.3200 181.4600 ;
        RECT 3305.7200 197.3000 3307.3200 197.7800 ;
        RECT 3305.7200 202.7400 3307.3200 203.2200 ;
        RECT 3305.7200 208.1800 3307.3200 208.6600 ;
        RECT 3305.7200 213.6200 3307.3200 214.1000 ;
        RECT 3305.7200 219.0600 3307.3200 219.5400 ;
        RECT 3305.7200 224.5000 3307.3200 224.9800 ;
        RECT 3305.7200 229.9400 3307.3200 230.4200 ;
        RECT 3361.4200 191.8600 3364.4200 192.3400 ;
        RECT 3361.4200 180.9800 3364.4200 181.4600 ;
        RECT 3361.4200 186.4200 3364.4200 186.9000 ;
        RECT 3361.4200 197.3000 3364.4200 197.7800 ;
        RECT 3361.4200 202.7400 3364.4200 203.2200 ;
        RECT 3361.4200 208.1800 3364.4200 208.6600 ;
        RECT 3361.4200 213.6200 3364.4200 214.1000 ;
        RECT 3361.4200 219.0600 3364.4200 219.5400 ;
        RECT 3361.4200 224.5000 3364.4200 224.9800 ;
        RECT 3361.4200 229.9400 3364.4200 230.4200 ;
        RECT 3305.7200 235.3800 3307.3200 235.8600 ;
        RECT 3305.7200 240.8200 3307.3200 241.3000 ;
        RECT 3305.7200 246.2600 3307.3200 246.7400 ;
        RECT 3305.7200 251.7000 3307.3200 252.1800 ;
        RECT 3305.7200 257.1400 3307.3200 257.6200 ;
        RECT 3305.7200 268.0200 3307.3200 268.5000 ;
        RECT 3305.7200 262.5800 3307.3200 263.0600 ;
        RECT 3305.7200 273.4600 3307.3200 273.9400 ;
        RECT 3305.7200 278.9000 3307.3200 279.3800 ;
        RECT 3361.4200 235.3800 3364.4200 235.8600 ;
        RECT 3361.4200 240.8200 3364.4200 241.3000 ;
        RECT 3361.4200 246.2600 3364.4200 246.7400 ;
        RECT 3361.4200 251.7000 3364.4200 252.1800 ;
        RECT 3361.4200 257.1400 3364.4200 257.6200 ;
        RECT 3361.4200 262.5800 3364.4200 263.0600 ;
        RECT 3361.4200 268.0200 3364.4200 268.5000 ;
        RECT 3361.4200 273.4600 3364.4200 273.9400 ;
        RECT 3361.4200 278.9000 3364.4200 279.3800 ;
        RECT 3305.7200 284.3400 3307.3200 284.8200 ;
        RECT 3305.7200 289.7800 3307.3200 290.2600 ;
        RECT 3305.7200 295.2200 3307.3200 295.7000 ;
        RECT 3305.7200 300.6600 3307.3200 301.1400 ;
        RECT 3305.7200 306.1000 3307.3200 306.5800 ;
        RECT 3305.7200 311.5400 3307.3200 312.0200 ;
        RECT 3305.7200 316.9800 3307.3200 317.4600 ;
        RECT 3305.7200 322.4200 3307.3200 322.9000 ;
        RECT 3305.7200 327.8600 3307.3200 328.3400 ;
        RECT 3305.7200 333.3000 3307.3200 333.7800 ;
        RECT 3361.4200 284.3400 3364.4200 284.8200 ;
        RECT 3361.4200 289.7800 3364.4200 290.2600 ;
        RECT 3361.4200 295.2200 3364.4200 295.7000 ;
        RECT 3361.4200 300.6600 3364.4200 301.1400 ;
        RECT 3361.4200 306.1000 3364.4200 306.5800 ;
        RECT 3361.4200 311.5400 3364.4200 312.0200 ;
        RECT 3361.4200 316.9800 3364.4200 317.4600 ;
        RECT 3361.4200 322.4200 3364.4200 322.9000 ;
        RECT 3361.4200 327.8600 3364.4200 328.3400 ;
        RECT 3361.4200 333.3000 3364.4200 333.7800 ;
        RECT 3305.7200 349.6200 3307.3200 350.1000 ;
        RECT 3305.7200 344.1800 3307.3200 344.6600 ;
        RECT 3305.7200 338.7400 3307.3200 339.2200 ;
        RECT 3305.7200 355.0600 3307.3200 355.5400 ;
        RECT 3305.7200 360.5000 3307.3200 360.9800 ;
        RECT 3305.7200 371.3800 3307.3200 371.8600 ;
        RECT 3305.7200 365.9400 3307.3200 366.4200 ;
        RECT 3305.7200 376.8200 3307.3200 377.3000 ;
        RECT 3305.7200 382.2600 3307.3200 382.7400 ;
        RECT 3305.7200 387.7000 3307.3200 388.1800 ;
        RECT 3361.4200 349.6200 3364.4200 350.1000 ;
        RECT 3361.4200 338.7400 3364.4200 339.2200 ;
        RECT 3361.4200 344.1800 3364.4200 344.6600 ;
        RECT 3361.4200 355.0600 3364.4200 355.5400 ;
        RECT 3361.4200 360.5000 3364.4200 360.9800 ;
        RECT 3361.4200 365.9400 3364.4200 366.4200 ;
        RECT 3361.4200 371.3800 3364.4200 371.8600 ;
        RECT 3361.4200 376.8200 3364.4200 377.3000 ;
        RECT 3361.4200 382.2600 3364.4200 382.7400 ;
        RECT 3361.4200 387.7000 3364.4200 388.1800 ;
        RECT 3305.7200 393.1400 3307.3200 393.6200 ;
        RECT 3305.7200 398.5800 3307.3200 399.0600 ;
        RECT 3305.7200 404.0200 3307.3200 404.5000 ;
        RECT 3305.7200 409.4600 3307.3200 409.9400 ;
        RECT 3305.7200 414.9000 3307.3200 415.3800 ;
        RECT 3305.7200 425.7800 3307.3200 426.2600 ;
        RECT 3305.7200 420.3400 3307.3200 420.8200 ;
        RECT 3305.7200 431.2200 3307.3200 431.7000 ;
        RECT 3305.7200 436.6600 3307.3200 437.1400 ;
        RECT 3361.4200 393.1400 3364.4200 393.6200 ;
        RECT 3361.4200 398.5800 3364.4200 399.0600 ;
        RECT 3361.4200 404.0200 3364.4200 404.5000 ;
        RECT 3361.4200 409.4600 3364.4200 409.9400 ;
        RECT 3361.4200 414.9000 3364.4200 415.3800 ;
        RECT 3361.4200 420.3400 3364.4200 420.8200 ;
        RECT 3361.4200 425.7800 3364.4200 426.2600 ;
        RECT 3361.4200 431.2200 3364.4200 431.7000 ;
        RECT 3361.4200 436.6600 3364.4200 437.1400 ;
        RECT 1733.7400 621.0200 1735.3400 621.5000 ;
        RECT 1941.3000 627.3700 1942.9000 628.9700 ;
        RECT 1953.9600 619.8600 1955.5600 620.3400 ;
        RECT 1733.7400 850.6600 1735.3400 851.1400 ;
        RECT 2174.1800 621.0200 2175.7800 621.5000 ;
        RECT 2166.8200 627.3700 2168.4200 630.0200 ;
        RECT 2447.1800 447.5400 2448.7800 448.0200 ;
        RECT 2447.1800 452.9800 2448.7800 453.4600 ;
        RECT 2447.1800 458.4200 2448.7800 458.9000 ;
        RECT 2447.1800 463.8600 2448.7800 464.3400 ;
        RECT 2447.1800 469.3000 2448.7800 469.7800 ;
        RECT 2447.1800 474.7400 2448.7800 475.2200 ;
        RECT 2447.1800 480.1800 2448.7800 480.6600 ;
        RECT 2447.1800 485.6200 2448.7800 486.1000 ;
        RECT 2447.1800 491.0600 2448.7800 491.5400 ;
        RECT 2492.9200 452.9800 2494.5200 453.4600 ;
        RECT 2492.9200 447.5400 2494.5200 448.0200 ;
        RECT 2492.9200 458.4200 2494.5200 458.9000 ;
        RECT 2492.9200 463.8600 2494.5200 464.3400 ;
        RECT 2492.9200 469.3000 2494.5200 469.7800 ;
        RECT 2492.9200 474.7400 2494.5200 475.2200 ;
        RECT 2492.9200 480.1800 2494.5200 480.6600 ;
        RECT 2492.9200 485.6200 2494.5200 486.1000 ;
        RECT 2492.9200 491.0600 2494.5200 491.5400 ;
        RECT 2447.1800 496.5000 2448.7800 496.9800 ;
        RECT 2447.1800 501.9400 2448.7800 502.4200 ;
        RECT 2447.1800 507.3800 2448.7800 507.8600 ;
        RECT 2447.1800 512.8200 2448.7800 513.3000 ;
        RECT 2447.1800 518.2600 2448.7800 518.7400 ;
        RECT 2447.1800 523.7000 2448.7800 524.1800 ;
        RECT 2447.1800 529.1400 2448.7800 529.6200 ;
        RECT 2447.1800 534.5800 2448.7800 535.0600 ;
        RECT 2447.1800 540.0200 2448.7800 540.5000 ;
        RECT 2447.1800 545.4600 2448.7800 545.9400 ;
        RECT 2492.9200 501.9400 2494.5200 502.4200 ;
        RECT 2492.9200 496.5000 2494.5200 496.9800 ;
        RECT 2492.9200 507.3800 2494.5200 507.8600 ;
        RECT 2492.9200 512.8200 2494.5200 513.3000 ;
        RECT 2492.9200 518.2600 2494.5200 518.7400 ;
        RECT 2492.9200 529.1400 2494.5200 529.6200 ;
        RECT 2492.9200 523.7000 2494.5200 524.1800 ;
        RECT 2492.9200 534.5800 2494.5200 535.0600 ;
        RECT 2492.9200 540.0200 2494.5200 540.5000 ;
        RECT 2492.9200 545.4600 2494.5200 545.9400 ;
        RECT 2394.4000 621.0200 2396.0000 621.5000 ;
        RECT 2447.1800 599.8600 2448.7800 600.3400 ;
        RECT 2492.9200 599.8600 2494.5200 600.3400 ;
        RECT 2447.1800 550.9000 2448.7800 551.3800 ;
        RECT 2447.1800 556.3400 2448.7800 556.8200 ;
        RECT 2447.1800 561.7800 2448.7800 562.2600 ;
        RECT 2447.1800 567.2200 2448.7800 567.7000 ;
        RECT 2447.1800 572.6600 2448.7800 573.1400 ;
        RECT 2447.1800 578.1000 2448.7800 578.5800 ;
        RECT 2447.1800 583.5400 2448.7800 584.0200 ;
        RECT 2447.1800 588.9800 2448.7800 589.4600 ;
        RECT 2447.1800 594.4200 2448.7800 594.9000 ;
        RECT 2492.9200 550.9000 2494.5200 551.3800 ;
        RECT 2492.9200 556.3400 2494.5200 556.8200 ;
        RECT 2492.9200 561.7800 2494.5200 562.2600 ;
        RECT 2492.9200 567.2200 2494.5200 567.7000 ;
        RECT 2492.9200 572.6600 2494.5200 573.1400 ;
        RECT 2492.9200 583.5400 2494.5200 584.0200 ;
        RECT 2492.9200 578.1000 2494.5200 578.5800 ;
        RECT 2492.9200 588.9800 2494.5200 589.4600 ;
        RECT 2492.9200 594.4200 2494.5200 594.9000 ;
        RECT 2447.1800 605.3000 2448.7800 605.7800 ;
        RECT 2447.1800 610.7400 2448.7800 611.2200 ;
        RECT 2447.1800 616.1800 2448.7800 616.6600 ;
        RECT 2447.1800 621.6200 2448.7800 622.1000 ;
        RECT 2447.1800 627.0600 2448.7800 628.9700 ;
        RECT 2447.1800 632.5000 2448.7800 632.9800 ;
        RECT 2447.1800 637.9400 2448.7800 638.4200 ;
        RECT 2447.1800 643.3800 2448.7800 643.8600 ;
        RECT 2447.1800 648.8200 2448.7800 649.3000 ;
        RECT 2492.9200 610.7400 2494.5200 611.2200 ;
        RECT 2492.9200 605.3000 2494.5200 605.7800 ;
        RECT 2492.9200 616.1800 2494.5200 616.6600 ;
        RECT 2492.9200 621.6200 2494.5200 622.1000 ;
        RECT 2492.9200 627.0600 2494.5200 627.5400 ;
        RECT 2492.9200 632.5000 2494.5200 632.9800 ;
        RECT 2492.9200 637.9400 2494.5200 638.4200 ;
        RECT 2492.9200 643.3800 2494.5200 643.8600 ;
        RECT 2492.9200 648.8200 2494.5200 649.3000 ;
        RECT 2174.1800 850.6600 2175.7800 851.1400 ;
        RECT 2447.1800 654.2600 2448.7800 654.7400 ;
        RECT 2447.1800 659.7000 2448.7800 660.1800 ;
        RECT 2447.1800 665.1400 2448.7800 665.6200 ;
        RECT 2447.1800 670.5800 2448.7800 671.0600 ;
        RECT 2447.1800 676.0200 2448.7800 676.5000 ;
        RECT 2447.1800 692.3400 2448.7800 692.8200 ;
        RECT 2447.1800 681.4600 2448.7800 681.9400 ;
        RECT 2447.1800 686.9000 2448.7800 687.3800 ;
        RECT 2447.1800 697.7800 2448.7800 698.2600 ;
        RECT 2447.1800 703.2200 2448.7800 703.7000 ;
        RECT 2492.9200 654.2600 2494.5200 654.7400 ;
        RECT 2492.9200 659.7000 2494.5200 660.1800 ;
        RECT 2492.9200 665.1400 2494.5200 665.6200 ;
        RECT 2492.9200 670.5800 2494.5200 671.0600 ;
        RECT 2492.9200 676.0200 2494.5200 676.5000 ;
        RECT 2492.9200 692.3400 2494.5200 692.8200 ;
        RECT 2492.9200 686.9000 2494.5200 687.3800 ;
        RECT 2492.9200 681.4600 2494.5200 681.9400 ;
        RECT 2492.9200 697.7800 2494.5200 698.2600 ;
        RECT 2492.9200 703.2200 2494.5200 703.7000 ;
        RECT 2447.1800 708.6600 2448.7800 709.1400 ;
        RECT 2447.1800 714.1000 2448.7800 714.5800 ;
        RECT 2447.1800 719.5400 2448.7800 720.0200 ;
        RECT 2447.1800 724.9800 2448.7800 725.4600 ;
        RECT 2447.1800 730.4200 2448.7800 730.9000 ;
        RECT 2447.1800 741.3000 2448.7800 741.7800 ;
        RECT 2447.1800 735.8600 2448.7800 736.3400 ;
        RECT 2447.1800 746.7400 2448.7800 747.2200 ;
        RECT 2492.9200 708.6600 2494.5200 709.1400 ;
        RECT 2492.9200 714.1000 2494.5200 714.5800 ;
        RECT 2492.9200 719.5400 2494.5200 720.0200 ;
        RECT 2492.9200 724.9800 2494.5200 725.4600 ;
        RECT 2492.9200 730.4200 2494.5200 730.9000 ;
        RECT 2492.9200 735.8600 2494.5200 736.3400 ;
        RECT 2492.9200 741.3000 2494.5200 741.7800 ;
        RECT 2492.9200 746.7400 2494.5200 747.2200 ;
        RECT 2394.4000 850.6600 2396.0000 851.1400 ;
        RECT 1733.7400 1080.3000 1735.3400 1080.7800 ;
        RECT 1941.3000 1086.6500 1942.9000 1088.2500 ;
        RECT 1953.9600 1079.1400 1955.5600 1079.6200 ;
        RECT 2166.8200 1086.6500 2168.4200 1089.3000 ;
        RECT 2174.1800 1080.3000 2175.7800 1080.7800 ;
        RECT 2394.4000 1080.3000 2396.0000 1080.7800 ;
        RECT 3305.7200 452.9800 3307.3200 453.4600 ;
        RECT 3305.7200 447.5400 3307.3200 448.0200 ;
        RECT 3305.7200 458.4200 3307.3200 458.9000 ;
        RECT 3305.7200 463.8600 3307.3200 464.3400 ;
        RECT 3305.7200 469.3000 3307.3200 469.7800 ;
        RECT 3305.7200 474.7400 3307.3200 475.2200 ;
        RECT 3305.7200 480.1800 3307.3200 480.6600 ;
        RECT 3305.7200 485.6200 3307.3200 486.1000 ;
        RECT 3305.7200 491.0600 3307.3200 491.5400 ;
        RECT 3361.4200 447.5400 3364.4200 448.0200 ;
        RECT 3361.4200 452.9800 3364.4200 453.4600 ;
        RECT 3361.4200 458.4200 3364.4200 458.9000 ;
        RECT 3361.4200 463.8600 3364.4200 464.3400 ;
        RECT 3361.4200 469.3000 3364.4200 469.7800 ;
        RECT 3361.4200 474.7400 3364.4200 475.2200 ;
        RECT 3361.4200 480.1800 3364.4200 480.6600 ;
        RECT 3361.4200 485.6200 3364.4200 486.1000 ;
        RECT 3361.4200 491.0600 3364.4200 491.5400 ;
        RECT 3305.7200 501.9400 3307.3200 502.4200 ;
        RECT 3305.7200 496.5000 3307.3200 496.9800 ;
        RECT 3305.7200 507.3800 3307.3200 507.8600 ;
        RECT 3305.7200 512.8200 3307.3200 513.3000 ;
        RECT 3305.7200 518.2600 3307.3200 518.7400 ;
        RECT 3305.7200 529.1400 3307.3200 529.6200 ;
        RECT 3305.7200 523.7000 3307.3200 524.1800 ;
        RECT 3305.7200 534.5800 3307.3200 535.0600 ;
        RECT 3305.7200 540.0200 3307.3200 540.5000 ;
        RECT 3305.7200 545.4600 3307.3200 545.9400 ;
        RECT 3361.4200 496.5000 3364.4200 496.9800 ;
        RECT 3361.4200 501.9400 3364.4200 502.4200 ;
        RECT 3361.4200 507.3800 3364.4200 507.8600 ;
        RECT 3361.4200 512.8200 3364.4200 513.3000 ;
        RECT 3361.4200 518.2600 3364.4200 518.7400 ;
        RECT 3361.4200 523.7000 3364.4200 524.1800 ;
        RECT 3361.4200 529.1400 3364.4200 529.6200 ;
        RECT 3361.4200 534.5800 3364.4200 535.0600 ;
        RECT 3361.4200 540.0200 3364.4200 540.5000 ;
        RECT 3361.4200 545.4600 3364.4200 545.9400 ;
        RECT 3361.4200 599.8600 3364.4200 600.3400 ;
        RECT 3305.7200 599.8600 3307.3200 600.3400 ;
        RECT 3305.7200 550.9000 3307.3200 551.3800 ;
        RECT 3305.7200 556.3400 3307.3200 556.8200 ;
        RECT 3305.7200 561.7800 3307.3200 562.2600 ;
        RECT 3305.7200 567.2200 3307.3200 567.7000 ;
        RECT 3305.7200 572.6600 3307.3200 573.1400 ;
        RECT 3305.7200 583.5400 3307.3200 584.0200 ;
        RECT 3305.7200 578.1000 3307.3200 578.5800 ;
        RECT 3305.7200 588.9800 3307.3200 589.4600 ;
        RECT 3305.7200 594.4200 3307.3200 594.9000 ;
        RECT 3361.4200 550.9000 3364.4200 551.3800 ;
        RECT 3361.4200 556.3400 3364.4200 556.8200 ;
        RECT 3361.4200 561.7800 3364.4200 562.2600 ;
        RECT 3361.4200 567.2200 3364.4200 567.7000 ;
        RECT 3361.4200 572.6600 3364.4200 573.1400 ;
        RECT 3361.4200 578.1000 3364.4200 578.5800 ;
        RECT 3361.4200 583.5400 3364.4200 584.0200 ;
        RECT 3361.4200 588.9800 3364.4200 589.4600 ;
        RECT 3361.4200 594.4200 3364.4200 594.9000 ;
        RECT 3305.7200 610.7400 3307.3200 611.2200 ;
        RECT 3305.7200 605.3000 3307.3200 605.7800 ;
        RECT 3305.7200 616.1800 3307.3200 616.6600 ;
        RECT 3305.7200 621.6200 3307.3200 622.1000 ;
        RECT 3305.7200 627.0600 3307.3200 627.5400 ;
        RECT 3305.7200 632.5000 3307.3200 632.9800 ;
        RECT 3305.7200 637.9400 3307.3200 638.4200 ;
        RECT 3305.7200 643.3800 3307.3200 643.8600 ;
        RECT 3305.7200 648.8200 3307.3200 649.3000 ;
        RECT 3361.4200 605.3000 3364.4200 605.7800 ;
        RECT 3361.4200 610.7400 3364.4200 611.2200 ;
        RECT 3361.4200 616.1800 3364.4200 616.6600 ;
        RECT 3361.4200 621.6200 3364.4200 622.1000 ;
        RECT 3361.4200 627.0600 3364.4200 627.5400 ;
        RECT 3361.4200 632.5000 3364.4200 632.9800 ;
        RECT 3361.4200 637.9400 3364.4200 638.4200 ;
        RECT 3361.4200 643.3800 3364.4200 643.8600 ;
        RECT 3361.4200 648.8200 3364.4200 649.3000 ;
        RECT 3305.7200 654.2600 3307.3200 654.7400 ;
        RECT 3305.7200 659.7000 3307.3200 660.1800 ;
        RECT 3305.7200 665.1400 3307.3200 665.6200 ;
        RECT 3305.7200 670.5800 3307.3200 671.0600 ;
        RECT 3305.7200 676.0200 3307.3200 676.5000 ;
        RECT 3305.7200 692.3400 3307.3200 692.8200 ;
        RECT 3305.7200 686.9000 3307.3200 687.3800 ;
        RECT 3305.7200 681.4600 3307.3200 681.9400 ;
        RECT 3305.7200 697.7800 3307.3200 698.2600 ;
        RECT 3305.7200 703.2200 3307.3200 703.7000 ;
        RECT 3361.4200 654.2600 3364.4200 654.7400 ;
        RECT 3361.4200 659.7000 3364.4200 660.1800 ;
        RECT 3361.4200 665.1400 3364.4200 665.6200 ;
        RECT 3361.4200 670.5800 3364.4200 671.0600 ;
        RECT 3361.4200 676.0200 3364.4200 676.5000 ;
        RECT 3361.4200 692.3400 3364.4200 692.8200 ;
        RECT 3361.4200 681.4600 3364.4200 681.9400 ;
        RECT 3361.4200 686.9000 3364.4200 687.3800 ;
        RECT 3361.4200 697.7800 3364.4200 698.2600 ;
        RECT 3361.4200 703.2200 3364.4200 703.7000 ;
        RECT 3305.7200 708.6600 3307.3200 709.1400 ;
        RECT 3305.7200 714.1000 3307.3200 714.5800 ;
        RECT 3305.7200 719.5400 3307.3200 720.0200 ;
        RECT 3305.7200 724.9800 3307.3200 725.4600 ;
        RECT 3305.7200 730.4200 3307.3200 730.9000 ;
        RECT 3305.7200 735.8600 3307.3200 736.3400 ;
        RECT 3305.7200 741.3000 3307.3200 741.7800 ;
        RECT 3305.7200 746.7400 3307.3200 747.2200 ;
        RECT 3305.7200 752.1800 3307.3200 752.6600 ;
        RECT 3305.7200 757.6200 3307.3200 758.1000 ;
        RECT 3361.4200 708.6600 3364.4200 709.1400 ;
        RECT 3361.4200 714.1000 3364.4200 714.5800 ;
        RECT 3361.4200 719.5400 3364.4200 720.0200 ;
        RECT 3361.4200 724.9800 3364.4200 725.4600 ;
        RECT 3361.4200 730.4200 3364.4200 730.9000 ;
        RECT 3361.4200 735.8600 3364.4200 736.3400 ;
        RECT 3361.4200 741.3000 3364.4200 741.7800 ;
        RECT 3361.4200 746.7400 3364.4200 747.2200 ;
        RECT 3361.4200 752.1800 3364.4200 752.6600 ;
        RECT 3361.4200 757.6200 3364.4200 758.1000 ;
        RECT 3305.7200 763.0600 3307.3200 763.5400 ;
        RECT 3305.7200 768.5000 3307.3200 768.9800 ;
        RECT 3305.7200 773.9400 3307.3200 774.4200 ;
        RECT 3305.7200 779.3800 3307.3200 779.8600 ;
        RECT 3305.7200 784.8200 3307.3200 785.3000 ;
        RECT 3305.7200 790.2600 3307.3200 790.7400 ;
        RECT 3305.7200 795.7000 3307.3200 796.1800 ;
        RECT 3305.7200 801.1400 3307.3200 801.6200 ;
        RECT 3305.7200 806.5800 3307.3200 807.0600 ;
        RECT 3361.4200 763.0600 3364.4200 763.5400 ;
        RECT 3361.4200 768.5000 3364.4200 768.9800 ;
        RECT 3361.4200 773.9400 3364.4200 774.4200 ;
        RECT 3361.4200 779.3800 3364.4200 779.8600 ;
        RECT 3361.4200 784.8200 3364.4200 785.3000 ;
        RECT 3361.4200 790.2600 3364.4200 790.7400 ;
        RECT 3361.4200 795.7000 3364.4200 796.1800 ;
        RECT 3361.4200 801.1400 3364.4200 801.6200 ;
        RECT 3361.4200 806.5800 3364.4200 807.0600 ;
        RECT 3305.7200 812.0200 3307.3200 812.5000 ;
        RECT 3305.7200 817.4600 3307.3200 817.9400 ;
        RECT 3305.7200 822.9000 3307.3200 823.3800 ;
        RECT 3305.7200 828.3400 3307.3200 828.8200 ;
        RECT 3305.7200 833.7800 3307.3200 834.2600 ;
        RECT 3305.7200 850.1000 3307.3200 850.5800 ;
        RECT 3305.7200 839.2200 3307.3200 839.7000 ;
        RECT 3305.7200 844.6600 3307.3200 845.1400 ;
        RECT 3305.7200 855.5400 3307.3200 856.0200 ;
        RECT 3305.7200 860.9800 3307.3200 861.4600 ;
        RECT 3361.4200 812.0200 3364.4200 812.5000 ;
        RECT 3361.4200 817.4600 3364.4200 817.9400 ;
        RECT 3361.4200 822.9000 3364.4200 823.3800 ;
        RECT 3361.4200 828.3400 3364.4200 828.8200 ;
        RECT 3361.4200 833.7800 3364.4200 834.2600 ;
        RECT 3361.4200 850.1000 3364.4200 850.5800 ;
        RECT 3361.4200 839.2200 3364.4200 839.7000 ;
        RECT 3361.4200 844.6600 3364.4200 845.1400 ;
        RECT 3361.4200 855.5400 3364.4200 856.0200 ;
        RECT 3361.4200 860.9800 3364.4200 861.4600 ;
        RECT 3305.7200 866.4200 3307.3200 866.9000 ;
        RECT 3305.7200 871.8600 3307.3200 872.3400 ;
        RECT 3305.7200 877.3000 3307.3200 877.7800 ;
        RECT 3305.7200 882.7400 3307.3200 883.2200 ;
        RECT 3305.7200 888.1800 3307.3200 888.6600 ;
        RECT 3305.7200 893.6200 3307.3200 894.1000 ;
        RECT 3305.7200 899.0600 3307.3200 899.5400 ;
        RECT 3305.7200 904.5000 3307.3200 904.9800 ;
        RECT 3305.7200 909.9400 3307.3200 910.4200 ;
        RECT 3305.7200 915.3800 3307.3200 915.8600 ;
        RECT 3361.4200 866.4200 3364.4200 866.9000 ;
        RECT 3361.4200 871.8600 3364.4200 872.3400 ;
        RECT 3361.4200 877.3000 3364.4200 877.7800 ;
        RECT 3361.4200 882.7400 3364.4200 883.2200 ;
        RECT 3361.4200 888.1800 3364.4200 888.6600 ;
        RECT 3361.4200 893.6200 3364.4200 894.1000 ;
        RECT 3361.4200 899.0600 3364.4200 899.5400 ;
        RECT 3361.4200 904.5000 3364.4200 904.9800 ;
        RECT 3361.4200 909.9400 3364.4200 910.4200 ;
        RECT 3361.4200 915.3800 3364.4200 915.8600 ;
        RECT 3305.7200 920.8200 3307.3200 921.3000 ;
        RECT 3305.7200 926.2600 3307.3200 926.7400 ;
        RECT 3305.7200 931.7000 3307.3200 932.1800 ;
        RECT 3305.7200 937.1400 3307.3200 937.6200 ;
        RECT 3305.7200 942.5800 3307.3200 943.0600 ;
        RECT 3305.7200 948.0200 3307.3200 948.5000 ;
        RECT 3305.7200 953.4600 3307.3200 953.9400 ;
        RECT 3305.7200 958.9000 3307.3200 959.3800 ;
        RECT 3305.7200 964.3400 3307.3200 964.8200 ;
        RECT 3361.4200 920.8200 3364.4200 921.3000 ;
        RECT 3361.4200 926.2600 3364.4200 926.7400 ;
        RECT 3361.4200 931.7000 3364.4200 932.1800 ;
        RECT 3361.4200 937.1400 3364.4200 937.6200 ;
        RECT 3361.4200 942.5800 3364.4200 943.0600 ;
        RECT 3361.4200 948.0200 3364.4200 948.5000 ;
        RECT 3361.4200 953.4600 3364.4200 953.9400 ;
        RECT 3361.4200 958.9000 3364.4200 959.3800 ;
        RECT 3361.4200 964.3400 3364.4200 964.8200 ;
        RECT 3305.7200 969.7800 3307.3200 970.2600 ;
        RECT 3305.7200 975.2200 3307.3200 975.7000 ;
        RECT 3305.7200 980.6600 3307.3200 981.1400 ;
        RECT 3305.7200 986.1000 3307.3200 986.5800 ;
        RECT 3305.7200 991.5400 3307.3200 992.0200 ;
        RECT 3305.7200 996.9800 3307.3200 997.4600 ;
        RECT 3305.7200 1002.4200 3307.3200 1002.9000 ;
        RECT 3305.7200 1007.8600 3307.3200 1008.3400 ;
        RECT 3305.7200 1013.3000 3307.3200 1013.7800 ;
        RECT 3305.7200 1018.7400 3307.3200 1019.2200 ;
        RECT 3361.4200 969.7800 3364.4200 970.2600 ;
        RECT 3361.4200 975.2200 3364.4200 975.7000 ;
        RECT 3361.4200 980.6600 3364.4200 981.1400 ;
        RECT 3361.4200 986.1000 3364.4200 986.5800 ;
        RECT 3361.4200 991.5400 3364.4200 992.0200 ;
        RECT 3361.4200 996.9800 3364.4200 997.4600 ;
        RECT 3361.4200 1002.4200 3364.4200 1002.9000 ;
        RECT 3361.4200 1007.8600 3364.4200 1008.3400 ;
        RECT 3361.4200 1013.3000 3364.4200 1013.7800 ;
        RECT 3361.4200 1018.7400 3364.4200 1019.2200 ;
        RECT 3305.7200 1024.1800 3307.3200 1024.6600 ;
        RECT 3305.7200 1029.6200 3307.3200 1030.1000 ;
        RECT 3305.7200 1035.0600 3307.3200 1035.5400 ;
        RECT 3305.7200 1040.5000 3307.3200 1040.9800 ;
        RECT 3305.7200 1045.9400 3307.3200 1046.4200 ;
        RECT 3305.7200 1051.3800 3307.3200 1051.8600 ;
        RECT 3305.7200 1056.8200 3307.3200 1057.3000 ;
        RECT 3305.7200 1062.2600 3307.3200 1062.7400 ;
        RECT 3305.7200 1067.7000 3307.3200 1068.1800 ;
        RECT 3305.7200 1073.1400 3307.3200 1073.6200 ;
        RECT 3361.4200 1024.1800 3364.4200 1024.6600 ;
        RECT 3361.4200 1029.6200 3364.4200 1030.1000 ;
        RECT 3361.4200 1035.0600 3364.4200 1035.5400 ;
        RECT 3361.4200 1040.5000 3364.4200 1040.9800 ;
        RECT 3361.4200 1045.9400 3364.4200 1046.4200 ;
        RECT 3361.4200 1051.3800 3364.4200 1051.8600 ;
        RECT 3361.4200 1056.8200 3364.4200 1057.3000 ;
        RECT 3361.4200 1062.2600 3364.4200 1062.7400 ;
        RECT 3361.4200 1067.7000 3364.4200 1068.1800 ;
        RECT 3361.4200 1073.1400 3364.4200 1073.6200 ;
        RECT 3305.7200 1100.3400 3307.3200 1100.8200 ;
        RECT 3305.7200 1078.5800 3307.3200 1079.0600 ;
        RECT 3305.7200 1084.0200 3307.3200 1084.5000 ;
        RECT 3305.7200 1089.4600 3307.3200 1089.9400 ;
        RECT 3305.7200 1094.9000 3307.3200 1095.3800 ;
        RECT 3305.7200 1105.7800 3307.3200 1106.2600 ;
        RECT 3305.7200 1111.2200 3307.3200 1111.7000 ;
        RECT 3305.7200 1116.6600 3307.3200 1117.1400 ;
        RECT 3305.7200 1122.1000 3307.3200 1122.5800 ;
        RECT 3361.4200 1100.3400 3364.4200 1100.8200 ;
        RECT 3361.4200 1078.5800 3364.4200 1079.0600 ;
        RECT 3361.4200 1084.0200 3364.4200 1084.5000 ;
        RECT 3361.4200 1089.4600 3364.4200 1089.9400 ;
        RECT 3361.4200 1094.9000 3364.4200 1095.3800 ;
        RECT 3361.4200 1105.7800 3364.4200 1106.2600 ;
        RECT 3361.4200 1111.2200 3364.4200 1111.7000 ;
        RECT 3361.4200 1116.6600 3364.4200 1117.1400 ;
        RECT 3361.4200 1122.1000 3364.4200 1122.5800 ;
        RECT 3305.7200 1127.5400 3307.3200 1128.0200 ;
        RECT 3305.7200 1132.9800 3307.3200 1133.4600 ;
        RECT 3305.7200 1138.4200 3307.3200 1138.9000 ;
        RECT 3305.7200 1143.8600 3307.3200 1144.3400 ;
        RECT 3305.7200 1149.3000 3307.3200 1149.7800 ;
        RECT 3305.7200 1154.7400 3307.3200 1155.2200 ;
        RECT 3305.7200 1160.1800 3307.3200 1160.6600 ;
        RECT 3305.7200 1165.6200 3307.3200 1166.1000 ;
        RECT 3305.7200 1171.0600 3307.3200 1171.5400 ;
        RECT 3305.7200 1176.5000 3307.3200 1176.9800 ;
        RECT 3361.4200 1127.5400 3364.4200 1128.0200 ;
        RECT 3361.4200 1132.9800 3364.4200 1133.4600 ;
        RECT 3361.4200 1138.4200 3364.4200 1138.9000 ;
        RECT 3361.4200 1143.8600 3364.4200 1144.3400 ;
        RECT 3361.4200 1149.3000 3364.4200 1149.7800 ;
        RECT 3361.4200 1154.7400 3364.4200 1155.2200 ;
        RECT 3361.4200 1160.1800 3364.4200 1160.6600 ;
        RECT 3361.4200 1165.6200 3364.4200 1166.1000 ;
        RECT 3361.4200 1171.0600 3364.4200 1171.5400 ;
        RECT 3361.4200 1176.5000 3364.4200 1176.9800 ;
        RECT 3305.7200 1181.9400 3307.3200 1182.4200 ;
        RECT 3305.7200 1187.3800 3307.3200 1187.8600 ;
        RECT 3305.7200 1192.8200 3307.3200 1193.3000 ;
        RECT 3305.7200 1198.2600 3307.3200 1198.7400 ;
        RECT 3305.7200 1203.7000 3307.3200 1204.1800 ;
        RECT 3305.7200 1209.1400 3307.3200 1209.6200 ;
        RECT 3305.7200 1214.5800 3307.3200 1215.0600 ;
        RECT 3305.7200 1220.0200 3307.3200 1220.5000 ;
        RECT 3305.7200 1225.4600 3307.3200 1225.9400 ;
        RECT 3305.7200 1230.9000 3307.3200 1231.3800 ;
        RECT 3361.4200 1181.9400 3364.4200 1182.4200 ;
        RECT 3361.4200 1187.3800 3364.4200 1187.8600 ;
        RECT 3361.4200 1192.8200 3364.4200 1193.3000 ;
        RECT 3361.4200 1198.2600 3364.4200 1198.7400 ;
        RECT 3361.4200 1203.7000 3364.4200 1204.1800 ;
        RECT 3361.4200 1209.1400 3364.4200 1209.6200 ;
        RECT 3361.4200 1214.5800 3364.4200 1215.0600 ;
        RECT 3361.4200 1220.0200 3364.4200 1220.5000 ;
        RECT 3361.4200 1225.4600 3364.4200 1225.9400 ;
        RECT 3361.4200 1230.9000 3364.4200 1231.3800 ;
        RECT 3305.7200 1258.1000 3307.3200 1258.5800 ;
        RECT 3305.7200 1236.3400 3307.3200 1236.8200 ;
        RECT 3305.7200 1241.7800 3307.3200 1242.2600 ;
        RECT 3305.7200 1247.2200 3307.3200 1247.7000 ;
        RECT 3305.7200 1252.6600 3307.3200 1253.1400 ;
        RECT 3305.7200 1263.5400 3307.3200 1264.0200 ;
        RECT 3305.7200 1268.9800 3307.3200 1269.4600 ;
        RECT 3305.7200 1274.4200 3307.3200 1274.9000 ;
        RECT 3305.7200 1279.8600 3307.3200 1280.3400 ;
        RECT 3361.4200 1258.1000 3364.4200 1258.5800 ;
        RECT 3361.4200 1236.3400 3364.4200 1236.8200 ;
        RECT 3361.4200 1241.7800 3364.4200 1242.2600 ;
        RECT 3361.4200 1247.2200 3364.4200 1247.7000 ;
        RECT 3361.4200 1252.6600 3364.4200 1253.1400 ;
        RECT 3361.4200 1263.5400 3364.4200 1264.0200 ;
        RECT 3361.4200 1268.9800 3364.4200 1269.4600 ;
        RECT 3361.4200 1274.4200 3364.4200 1274.9000 ;
        RECT 3361.4200 1279.8600 3364.4200 1280.3400 ;
        RECT 6.0000 1285.3000 9.0000 1285.7800 ;
        RECT 6.0000 1290.7400 9.0000 1291.2200 ;
        RECT 6.0000 1296.1800 9.0000 1296.6600 ;
        RECT 6.0000 1301.6200 9.0000 1302.1000 ;
        RECT 6.0000 1307.0600 9.0000 1307.5400 ;
        RECT 6.0000 1312.5000 9.0000 1312.9800 ;
        RECT 6.0000 1317.9400 9.0000 1318.4200 ;
        RECT 6.0000 1323.3800 9.0000 1323.8600 ;
        RECT 6.0000 1328.9900 9.0000 1329.4700 ;
        RECT 6.0000 1334.2600 9.0000 1334.7400 ;
        RECT 6.0000 1350.5800 9.0000 1351.0600 ;
        RECT 6.0000 1339.7000 9.0000 1340.1800 ;
        RECT 6.0000 1345.1400 9.0000 1345.6200 ;
        RECT 6.0000 1356.0200 9.0000 1356.5000 ;
        RECT 6.0000 1361.4600 9.0000 1361.9400 ;
        RECT 6.0000 1366.9000 9.0000 1367.3800 ;
        RECT 6.0000 1372.3400 9.0000 1372.8200 ;
        RECT 6.0000 1377.7800 9.0000 1378.2600 ;
        RECT 6.0000 1383.2200 9.0000 1383.7000 ;
        RECT 6.0000 1388.6600 9.0000 1389.1400 ;
        RECT 152.9200 1285.3000 154.5200 1285.7800 ;
        RECT 152.9200 1290.7400 154.5200 1291.2200 ;
        RECT 152.9200 1296.1800 154.5200 1296.6600 ;
        RECT 152.9200 1301.6200 154.5200 1302.1000 ;
        RECT 152.9200 1307.0600 154.5200 1307.5400 ;
        RECT 152.9200 1312.5000 154.5200 1312.9800 ;
        RECT 152.9200 1317.9400 154.5200 1318.4200 ;
        RECT 152.9200 1323.3800 154.5200 1323.8600 ;
        RECT 152.9200 1328.9900 154.5200 1329.4700 ;
        RECT 152.9200 1334.2600 154.5200 1334.7400 ;
        RECT 152.9200 1350.5800 154.5200 1351.0600 ;
        RECT 152.9200 1339.7000 154.5200 1340.1800 ;
        RECT 152.9200 1345.1400 154.5200 1345.6200 ;
        RECT 152.9200 1356.0200 154.5200 1356.5000 ;
        RECT 152.9200 1361.4600 154.5200 1361.9400 ;
        RECT 152.9200 1366.9000 154.5200 1367.3800 ;
        RECT 152.9200 1372.3400 154.5200 1372.8200 ;
        RECT 152.9200 1377.7800 154.5200 1378.2600 ;
        RECT 152.9200 1383.2200 154.5200 1383.7000 ;
        RECT 152.9200 1388.6600 154.5200 1389.1400 ;
        RECT 6.0000 1394.1000 9.0000 1394.5800 ;
        RECT 6.0000 1399.5400 9.0000 1400.0200 ;
        RECT 6.0000 1404.9800 9.0000 1405.4600 ;
        RECT 6.0000 1410.4200 9.0000 1410.9000 ;
        RECT 6.0000 1415.8600 9.0000 1416.3400 ;
        RECT 6.0000 1421.3000 9.0000 1421.7800 ;
        RECT 6.0000 1426.7400 9.0000 1427.2200 ;
        RECT 6.0000 1432.1800 9.0000 1432.6600 ;
        RECT 6.0000 1437.6200 9.0000 1438.1000 ;
        RECT 6.0000 1443.0600 9.0000 1443.5400 ;
        RECT 6.0000 1448.5000 9.0000 1448.9800 ;
        RECT 6.0000 1453.9400 9.0000 1454.4200 ;
        RECT 6.0000 1459.3800 9.0000 1459.8600 ;
        RECT 6.0000 1464.8200 9.0000 1465.3000 ;
        RECT 6.0000 1470.2600 9.0000 1470.7400 ;
        RECT 6.0000 1475.7000 9.0000 1476.1800 ;
        RECT 6.0000 1481.1400 9.0000 1481.6200 ;
        RECT 6.0000 1486.5800 9.0000 1487.0600 ;
        RECT 6.0000 1492.0200 9.0000 1492.5000 ;
        RECT 152.9200 1394.1000 154.5200 1394.5800 ;
        RECT 152.9200 1399.5400 154.5200 1400.0200 ;
        RECT 152.9200 1404.9800 154.5200 1405.4600 ;
        RECT 152.9200 1410.4200 154.5200 1410.9000 ;
        RECT 152.9200 1415.8600 154.5200 1416.3400 ;
        RECT 152.9200 1421.3000 154.5200 1421.7800 ;
        RECT 152.9200 1426.7400 154.5200 1427.2200 ;
        RECT 152.9200 1432.1800 154.5200 1432.6600 ;
        RECT 152.9200 1437.6200 154.5200 1438.1000 ;
        RECT 152.9200 1443.0600 154.5200 1443.5400 ;
        RECT 152.9200 1448.5000 154.5200 1448.9800 ;
        RECT 152.9200 1453.9400 154.5200 1454.4200 ;
        RECT 152.9200 1459.3800 154.5200 1459.8600 ;
        RECT 152.9200 1464.8200 154.5200 1465.3000 ;
        RECT 152.9200 1470.2600 154.5200 1470.7400 ;
        RECT 152.9200 1475.7000 154.5200 1476.1800 ;
        RECT 152.9200 1481.1400 154.5200 1481.6200 ;
        RECT 152.9200 1486.5800 154.5200 1487.0600 ;
        RECT 152.9200 1492.0200 154.5200 1492.5000 ;
        RECT 6.0000 1600.8200 9.0000 1601.3000 ;
        RECT 152.9200 1600.8200 154.5200 1601.3000 ;
        RECT 6.0000 1508.3400 9.0000 1508.8200 ;
        RECT 6.0000 1497.4600 9.0000 1497.9400 ;
        RECT 6.0000 1502.9000 9.0000 1503.3800 ;
        RECT 6.0000 1513.7800 9.0000 1514.2600 ;
        RECT 6.0000 1519.2200 9.0000 1519.7000 ;
        RECT 6.0000 1524.6600 9.0000 1525.1400 ;
        RECT 6.0000 1530.1000 9.0000 1530.5800 ;
        RECT 6.0000 1535.5400 9.0000 1536.0200 ;
        RECT 6.0000 1540.9800 9.0000 1541.4600 ;
        RECT 6.0000 1546.4200 9.0000 1546.9000 ;
        RECT 6.0000 1551.8600 9.0000 1552.3400 ;
        RECT 6.0000 1558.8300 9.0000 1559.3100 ;
        RECT 6.0000 1562.7400 9.0000 1563.2200 ;
        RECT 6.0000 1568.1800 9.0000 1568.6600 ;
        RECT 6.0000 1573.6200 9.0000 1574.1000 ;
        RECT 6.0000 1579.0600 9.0000 1579.5400 ;
        RECT 6.0000 1584.5000 9.0000 1584.9800 ;
        RECT 6.0000 1589.9400 9.0000 1590.4200 ;
        RECT 6.0000 1595.3800 9.0000 1595.8600 ;
        RECT 152.9200 1508.3400 154.5200 1508.8200 ;
        RECT 152.9200 1497.4600 154.5200 1497.9400 ;
        RECT 152.9200 1502.9000 154.5200 1503.3800 ;
        RECT 152.9200 1513.7800 154.5200 1514.2600 ;
        RECT 152.9200 1519.2200 154.5200 1519.7000 ;
        RECT 152.9200 1524.6600 154.5200 1525.1400 ;
        RECT 152.9200 1530.1000 154.5200 1530.5800 ;
        RECT 152.9200 1535.5400 154.5200 1536.0200 ;
        RECT 152.9200 1540.9800 154.5200 1541.4600 ;
        RECT 152.9200 1546.4200 154.5200 1546.9000 ;
        RECT 152.9200 1551.8600 154.5200 1552.3400 ;
        RECT 152.9200 1562.7400 154.5200 1563.2200 ;
        RECT 152.9200 1568.1800 154.5200 1568.6600 ;
        RECT 152.9200 1573.6200 154.5200 1574.1000 ;
        RECT 152.9200 1579.0600 154.5200 1579.5400 ;
        RECT 152.9200 1584.5000 154.5200 1584.9800 ;
        RECT 152.9200 1589.9400 154.5200 1590.4200 ;
        RECT 152.9200 1595.3800 154.5200 1595.8600 ;
        RECT 6.0000 1606.2600 9.0000 1606.7400 ;
        RECT 6.0000 1611.7000 9.0000 1612.1800 ;
        RECT 6.0000 1617.1400 9.0000 1617.6200 ;
        RECT 6.0000 1622.5800 9.0000 1623.0600 ;
        RECT 6.0000 1628.0200 9.0000 1628.5000 ;
        RECT 6.0000 1633.4600 9.0000 1633.9400 ;
        RECT 6.0000 1638.9000 9.0000 1639.3800 ;
        RECT 6.0000 1644.3400 9.0000 1644.8200 ;
        RECT 6.0000 1649.7800 9.0000 1650.2600 ;
        RECT 6.0000 1655.2200 9.0000 1655.7000 ;
        RECT 6.0000 1660.6600 9.0000 1661.1400 ;
        RECT 6.0000 1666.1000 9.0000 1666.5800 ;
        RECT 6.0000 1671.5400 9.0000 1672.0200 ;
        RECT 6.0000 1676.9800 9.0000 1677.4600 ;
        RECT 6.0000 1682.4200 9.0000 1682.9000 ;
        RECT 6.0000 1687.8600 9.0000 1688.3400 ;
        RECT 6.0000 1693.3000 9.0000 1693.7800 ;
        RECT 6.0000 1698.7400 9.0000 1699.2200 ;
        RECT 6.0000 1704.1800 9.0000 1704.6600 ;
        RECT 152.9200 1606.2600 154.5200 1606.7400 ;
        RECT 152.9200 1611.7000 154.5200 1612.1800 ;
        RECT 152.9200 1617.1400 154.5200 1617.6200 ;
        RECT 152.9200 1622.5800 154.5200 1623.0600 ;
        RECT 152.9200 1628.0200 154.5200 1628.5000 ;
        RECT 152.9200 1633.4600 154.5200 1633.9400 ;
        RECT 152.9200 1638.9000 154.5200 1639.3800 ;
        RECT 152.9200 1644.3400 154.5200 1644.8200 ;
        RECT 152.9200 1649.7800 154.5200 1650.2600 ;
        RECT 152.9200 1655.2200 154.5200 1655.7000 ;
        RECT 152.9200 1660.6600 154.5200 1661.1400 ;
        RECT 152.9200 1666.1000 154.5200 1666.5800 ;
        RECT 152.9200 1671.5400 154.5200 1672.0200 ;
        RECT 152.9200 1676.9800 154.5200 1677.4600 ;
        RECT 152.9200 1682.4200 154.5200 1682.9000 ;
        RECT 152.9200 1687.8600 154.5200 1688.3400 ;
        RECT 152.9200 1693.3000 154.5200 1693.7800 ;
        RECT 152.9200 1698.7400 154.5200 1699.2200 ;
        RECT 152.9200 1704.1800 154.5200 1704.6600 ;
        RECT 6.0000 1916.3400 9.0000 1916.8200 ;
        RECT 152.9200 1916.3400 154.5200 1916.8200 ;
        RECT 6.0000 1758.5800 9.0000 1759.0600 ;
        RECT 6.0000 1709.6200 9.0000 1710.1000 ;
        RECT 6.0000 1715.0600 9.0000 1715.5400 ;
        RECT 6.0000 1720.5000 9.0000 1720.9800 ;
        RECT 6.0000 1725.9400 9.0000 1726.4200 ;
        RECT 6.0000 1731.3800 9.0000 1731.8600 ;
        RECT 6.0000 1736.8200 9.0000 1737.3000 ;
        RECT 6.0000 1742.2600 9.0000 1742.7400 ;
        RECT 6.0000 1747.7000 9.0000 1748.1800 ;
        RECT 6.0000 1753.1400 9.0000 1753.6200 ;
        RECT 6.0000 1783.7400 9.0000 1785.7500 ;
        RECT 6.0000 1764.0200 9.0000 1764.5000 ;
        RECT 6.0000 1769.4600 9.0000 1769.9400 ;
        RECT 6.0000 1774.9000 9.0000 1775.3800 ;
        RECT 6.0000 1780.3400 9.0000 1780.8200 ;
        RECT 6.0000 1791.2200 9.0000 1791.7000 ;
        RECT 6.0000 1796.6600 9.0000 1797.1400 ;
        RECT 6.0000 1802.1000 9.0000 1802.5800 ;
        RECT 6.0000 1807.5400 9.0000 1808.0200 ;
        RECT 152.9200 1758.5800 154.5200 1759.0600 ;
        RECT 152.9200 1709.6200 154.5200 1710.1000 ;
        RECT 152.9200 1715.0600 154.5200 1715.5400 ;
        RECT 152.9200 1720.5000 154.5200 1720.9800 ;
        RECT 152.9200 1725.9400 154.5200 1726.4200 ;
        RECT 152.9200 1731.3800 154.5200 1731.8600 ;
        RECT 152.9200 1736.8200 154.5200 1737.3000 ;
        RECT 152.9200 1742.2600 154.5200 1742.7400 ;
        RECT 152.9200 1747.7000 154.5200 1748.1800 ;
        RECT 152.9200 1753.1400 154.5200 1753.6200 ;
        RECT 152.9200 1783.7400 154.5200 1785.7500 ;
        RECT 152.9200 1764.0200 154.5200 1764.5000 ;
        RECT 152.9200 1769.4600 154.5200 1769.9400 ;
        RECT 152.9200 1774.9000 154.5200 1775.3800 ;
        RECT 152.9200 1780.3400 154.5200 1780.8200 ;
        RECT 152.9200 1791.2200 154.5200 1791.7000 ;
        RECT 152.9200 1796.6600 154.5200 1797.1400 ;
        RECT 152.9200 1802.1000 154.5200 1802.5800 ;
        RECT 152.9200 1807.5400 154.5200 1808.0200 ;
        RECT 6.0000 1812.9800 9.0000 1813.4600 ;
        RECT 6.0000 1818.4200 9.0000 1818.9000 ;
        RECT 6.0000 1823.8600 9.0000 1824.3400 ;
        RECT 6.0000 1829.3000 9.0000 1829.7800 ;
        RECT 6.0000 1834.7400 9.0000 1835.2200 ;
        RECT 6.0000 1840.1800 9.0000 1840.6600 ;
        RECT 6.0000 1845.6200 9.0000 1846.1000 ;
        RECT 6.0000 1851.0600 9.0000 1851.5400 ;
        RECT 6.0000 1856.5000 9.0000 1856.9800 ;
        RECT 6.0000 1861.9400 9.0000 1862.4200 ;
        RECT 6.0000 1867.3800 9.0000 1867.8600 ;
        RECT 6.0000 1872.8200 9.0000 1873.3000 ;
        RECT 6.0000 1878.2600 9.0000 1878.7400 ;
        RECT 6.0000 1883.7000 9.0000 1884.1800 ;
        RECT 6.0000 1889.1400 9.0000 1889.6200 ;
        RECT 6.0000 1894.5800 9.0000 1895.0600 ;
        RECT 6.0000 1900.0200 9.0000 1900.5000 ;
        RECT 6.0000 1905.4600 9.0000 1905.9400 ;
        RECT 6.0000 1910.9000 9.0000 1911.3800 ;
        RECT 152.9200 1812.9800 154.5200 1813.4600 ;
        RECT 152.9200 1818.4200 154.5200 1818.9000 ;
        RECT 152.9200 1823.8600 154.5200 1824.3400 ;
        RECT 152.9200 1829.3000 154.5200 1829.7800 ;
        RECT 152.9200 1834.7400 154.5200 1835.2200 ;
        RECT 152.9200 1840.1800 154.5200 1840.6600 ;
        RECT 152.9200 1845.6200 154.5200 1846.1000 ;
        RECT 152.9200 1851.0600 154.5200 1851.5400 ;
        RECT 152.9200 1856.5000 154.5200 1856.9800 ;
        RECT 152.9200 1861.9400 154.5200 1862.4200 ;
        RECT 152.9200 1867.3800 154.5200 1867.8600 ;
        RECT 152.9200 1872.8200 154.5200 1873.3000 ;
        RECT 152.9200 1878.2600 154.5200 1878.7400 ;
        RECT 152.9200 1883.7000 154.5200 1884.1800 ;
        RECT 152.9200 1889.1400 154.5200 1889.6200 ;
        RECT 152.9200 1894.5800 154.5200 1895.0600 ;
        RECT 152.9200 1900.0200 154.5200 1900.5000 ;
        RECT 152.9200 1905.4600 154.5200 1905.9400 ;
        RECT 152.9200 1910.9000 154.5200 1911.3800 ;
        RECT 6.0000 1921.7800 9.0000 1922.2600 ;
        RECT 6.0000 1927.2200 9.0000 1927.7000 ;
        RECT 6.0000 1932.6600 9.0000 1933.1400 ;
        RECT 6.0000 1938.1000 9.0000 1938.5800 ;
        RECT 6.0000 1943.5400 9.0000 1944.0200 ;
        RECT 6.0000 1948.9800 9.0000 1949.4600 ;
        RECT 6.0000 1954.4200 9.0000 1954.9000 ;
        RECT 6.0000 1959.8600 9.0000 1960.3400 ;
        RECT 6.0000 1965.3000 9.0000 1965.7800 ;
        RECT 6.0000 1970.7400 9.0000 1971.2200 ;
        RECT 6.0000 1976.1800 9.0000 1976.6600 ;
        RECT 6.0000 1981.6200 9.0000 1982.1000 ;
        RECT 6.0000 1987.0600 9.0000 1987.5400 ;
        RECT 6.0000 1992.5000 9.0000 1992.9800 ;
        RECT 6.0000 2008.8200 9.0000 2009.3000 ;
        RECT 6.0000 1997.9400 9.0000 1998.4200 ;
        RECT 6.0000 2003.3800 9.0000 2003.8600 ;
        RECT 6.0000 2019.7000 9.0000 2020.1800 ;
        RECT 152.9200 1921.7800 154.5200 1922.2600 ;
        RECT 152.9200 1927.2200 154.5200 1927.7000 ;
        RECT 152.9200 1932.6600 154.5200 1933.1400 ;
        RECT 152.9200 1938.1000 154.5200 1938.5800 ;
        RECT 152.9200 1943.5400 154.5200 1944.0200 ;
        RECT 152.9200 1948.9800 154.5200 1949.4600 ;
        RECT 152.9200 1954.4200 154.5200 1954.9000 ;
        RECT 152.9200 1959.8600 154.5200 1960.3400 ;
        RECT 152.9200 1965.3000 154.5200 1965.7800 ;
        RECT 152.9200 1970.7400 154.5200 1971.2200 ;
        RECT 152.9200 1976.1800 154.5200 1976.6600 ;
        RECT 152.9200 1981.6200 154.5200 1982.1000 ;
        RECT 152.9200 1987.0600 154.5200 1987.5400 ;
        RECT 152.9200 1992.5000 154.5200 1992.9800 ;
        RECT 152.9200 2008.8200 154.5200 2009.3000 ;
        RECT 152.9200 1997.9400 154.5200 1998.4200 ;
        RECT 152.9200 2003.3800 154.5200 2003.8600 ;
        RECT 6.0000 2025.1400 9.0000 2025.6200 ;
        RECT 6.0000 2030.5800 9.0000 2031.0600 ;
        RECT 6.0000 2036.0200 9.0000 2036.5000 ;
        RECT 6.0000 2041.4600 9.0000 2041.9400 ;
        RECT 6.0000 2046.9000 9.0000 2047.3800 ;
        RECT 6.0000 2052.3400 9.0000 2052.8200 ;
        RECT 6.0000 2057.7800 9.0000 2058.2600 ;
        RECT 6.0000 2063.2200 9.0000 2063.7000 ;
        RECT 6.0000 2068.6600 9.0000 2069.1400 ;
        RECT 6.0000 2074.1000 9.0000 2074.5800 ;
        RECT 6.0000 2079.5400 9.0000 2080.0200 ;
        RECT 6.0000 2084.9800 9.0000 2085.4600 ;
        RECT 6.0000 2090.4200 9.0000 2090.9000 ;
        RECT 6.0000 2095.8600 9.0000 2096.3400 ;
        RECT 6.0000 2101.3000 9.0000 2101.7800 ;
        RECT 6.0000 2106.7400 9.0000 2107.2200 ;
        RECT 6.0000 2112.1800 9.0000 2112.6600 ;
        RECT 6.0000 2117.6200 9.0000 2118.1000 ;
        RECT 6.0000 2123.0600 9.0000 2123.5400 ;
        RECT 1013.1800 1310.2000 1014.7800 1310.6800 ;
        RECT 1060.5600 1546.0900 1062.1600 1547.6900 ;
        RECT 1055.6000 1539.8400 1057.2000 1540.3200 ;
        RECT 1073.2200 1538.6800 1074.8200 1539.1600 ;
        RECT 1065.8600 1564.1300 1067.4600 1565.8300 ;
        RECT 1293.3000 1309.9400 1294.9000 1310.4200 ;
        RECT 1513.5200 1309.9400 1515.1200 1310.4200 ;
        RECT 1285.9400 1545.9300 1287.6800 1548.8400 ;
        RECT 1293.3000 1539.5800 1294.9000 1540.0600 ;
        RECT 1285.9400 1553.8400 1287.6800 1555.7000 ;
        RECT 1285.9400 1563.8700 1287.6800 1565.7300 ;
        RECT 1513.5200 1539.5800 1515.1200 1540.0600 ;
        RECT 1013.1800 1769.4800 1014.7800 1769.9600 ;
        RECT 965.7200 1970.7400 967.3200 1971.2200 ;
        RECT 965.7200 1976.1800 967.3200 1976.6600 ;
        RECT 965.7200 1981.6200 967.3200 1982.1000 ;
        RECT 965.7200 1987.0600 967.3200 1987.5400 ;
        RECT 965.7200 1992.5000 967.3200 1992.9800 ;
        RECT 965.7200 2008.8200 967.3200 2009.3000 ;
        RECT 965.7200 1997.9400 967.3200 1998.4200 ;
        RECT 965.7200 2003.3800 967.3200 2003.8600 ;
        RECT 1002.9200 1970.7400 1004.5200 1971.2200 ;
        RECT 1002.9200 1976.1800 1004.5200 1976.6600 ;
        RECT 1002.9200 1981.6200 1004.5200 1982.1000 ;
        RECT 1002.9200 1987.0600 1004.5200 1987.5400 ;
        RECT 1002.9200 1992.5000 1004.5200 1992.9800 ;
        RECT 1002.9200 2008.8200 1004.5200 2009.3000 ;
        RECT 1002.9200 1997.9400 1004.5200 1998.4200 ;
        RECT 1002.9200 2003.3800 1004.5200 2003.8600 ;
        RECT 1002.9200 2019.7000 1004.5200 2020.1800 ;
        RECT 1002.9200 2030.5800 1004.5200 2031.0600 ;
        RECT 1001.3300 2025.1400 1001.8300 2025.6200 ;
        RECT 1002.9200 2036.0200 1004.5200 2036.5000 ;
        RECT 1002.9200 2041.4600 1004.5200 2041.9400 ;
        RECT 1002.9200 2046.9000 1004.5200 2047.3800 ;
        RECT 1002.9200 2052.3400 1004.5200 2052.8200 ;
        RECT 1002.9200 2057.7800 1004.5200 2058.2600 ;
        RECT 1002.9200 2063.2200 1004.5200 2063.7000 ;
        RECT 1002.9200 2068.6600 1004.5200 2069.1400 ;
        RECT 1002.9200 2074.1000 1004.5200 2074.5800 ;
        RECT 1002.9200 2084.9800 1004.5200 2085.4600 ;
        RECT 1002.9200 2079.5400 1004.5200 2080.0200 ;
        RECT 1002.9200 2090.4200 1004.5200 2090.9000 ;
        RECT 1002.9200 2095.8600 1004.5200 2096.3400 ;
        RECT 1002.9200 2101.3000 1004.5200 2101.7800 ;
        RECT 1002.9200 2106.7400 1004.5200 2107.2200 ;
        RECT 1002.9200 2112.1800 1004.5200 2112.6600 ;
        RECT 1002.9200 2117.6200 1004.5200 2118.1000 ;
        RECT 1002.9200 2123.0600 1004.5200 2123.5400 ;
        RECT 1073.2200 1997.9600 1074.8200 1998.4400 ;
        RECT 1060.5600 2005.3700 1062.1600 2006.9700 ;
        RECT 1055.6000 1999.1200 1057.2000 1999.6000 ;
        RECT 1293.3000 1769.2200 1294.9000 1769.7000 ;
        RECT 1513.5200 1769.2200 1515.1200 1769.7000 ;
        RECT 1285.9400 2013.1200 1287.6800 2014.9800 ;
        RECT 1285.9400 2005.2100 1287.6800 2008.1200 ;
        RECT 1293.3000 1998.8600 1294.9000 1999.3400 ;
        RECT 1285.9400 2023.1500 1287.6800 2025.0100 ;
        RECT 1513.5200 1998.8600 1515.1200 1999.3400 ;
        RECT 6.0000 2128.5000 9.0000 2128.9800 ;
        RECT 6.0000 2133.9400 9.0000 2134.4200 ;
        RECT 6.0000 2139.3800 9.0000 2139.8600 ;
        RECT 6.0000 2144.8200 9.0000 2145.3000 ;
        RECT 6.0000 2150.2600 9.0000 2150.7400 ;
        RECT 6.0000 2166.5800 9.0000 2167.0600 ;
        RECT 6.0000 2155.7000 9.0000 2156.1800 ;
        RECT 6.0000 2161.1400 9.0000 2161.6200 ;
        RECT 6.0000 2172.0200 9.0000 2172.5000 ;
        RECT 6.0000 2177.4600 9.0000 2177.9400 ;
        RECT 6.0000 2182.9000 9.0000 2183.3800 ;
        RECT 6.0000 2188.3400 9.0000 2188.8200 ;
        RECT 6.0000 2193.7800 9.0000 2194.2600 ;
        RECT 6.0000 2199.2200 9.0000 2199.7000 ;
        RECT 6.0000 2204.6600 9.0000 2205.1400 ;
        RECT 6.0000 2210.1000 9.0000 2210.5800 ;
        RECT 6.0000 2215.5400 9.0000 2216.0200 ;
        RECT 6.0000 2220.9800 9.0000 2221.4600 ;
        RECT 6.0000 2226.4200 9.0000 2226.9000 ;
        RECT 6.0000 2231.8600 9.0000 2232.3400 ;
        RECT 6.0000 2259.0600 9.0000 2259.5400 ;
        RECT 6.0000 2237.3000 9.0000 2237.7800 ;
        RECT 6.0000 2242.7400 9.0000 2244.6200 ;
        RECT 6.0000 2248.1800 9.0000 2248.6600 ;
        RECT 6.0000 2253.6200 9.0000 2254.1000 ;
        RECT 6.0000 2264.5000 9.0000 2264.9800 ;
        RECT 6.0000 2269.9400 9.0000 2270.4200 ;
        RECT 6.0000 2275.3800 9.0000 2275.8600 ;
        RECT 6.0000 2280.8200 9.0000 2281.3000 ;
        RECT 6.0000 2286.2600 9.0000 2286.7400 ;
        RECT 6.0000 2291.7000 9.0000 2292.1800 ;
        RECT 6.0000 2297.1400 9.0000 2297.6200 ;
        RECT 6.0000 2302.5800 9.0000 2303.0600 ;
        RECT 6.0000 2308.0200 9.0000 2308.5000 ;
        RECT 6.0000 2313.4600 9.0000 2313.9400 ;
        RECT 6.0000 2318.9000 9.0000 2319.3800 ;
        RECT 6.0000 2324.3400 9.0000 2324.8200 ;
        RECT 6.0000 2329.7800 9.0000 2330.2600 ;
        RECT 6.0000 2335.2200 9.0000 2335.7000 ;
        RECT 6.0000 2340.6600 9.0000 2341.1400 ;
        RECT 6.0000 2346.1000 9.0000 2346.5800 ;
        RECT 6.0000 2351.5400 9.0000 2352.0200 ;
        RECT 6.0000 2356.9800 9.0000 2357.4600 ;
        RECT 6.0000 2362.4200 9.0000 2362.9000 ;
        RECT 6.0000 2367.8600 9.0000 2368.3400 ;
        RECT 6.0000 2373.3000 9.0000 2373.7800 ;
        RECT 6.0000 2378.7400 9.0000 2379.2200 ;
        RECT 6.0000 2384.1800 9.0000 2384.6600 ;
        RECT 6.0000 2389.6200 9.0000 2390.1000 ;
        RECT 6.0000 2416.8200 9.0000 2417.3000 ;
        RECT 6.0000 2395.0600 9.0000 2395.5400 ;
        RECT 6.0000 2400.5000 9.0000 2400.9800 ;
        RECT 6.0000 2405.9400 9.0000 2406.4200 ;
        RECT 6.0000 2411.3800 9.0000 2411.8600 ;
        RECT 6.0000 2422.2600 9.0000 2422.7400 ;
        RECT 6.0000 2427.7000 9.0000 2428.1800 ;
        RECT 6.0000 2433.1400 9.0000 2433.6200 ;
        RECT 6.0000 2438.5800 9.0000 2439.0600 ;
        RECT 6.0000 2444.0200 9.0000 2444.5000 ;
        RECT 6.0000 2449.4600 9.0000 2449.9400 ;
        RECT 6.0000 2454.9000 9.0000 2455.3800 ;
        RECT 6.0000 2460.3400 9.0000 2460.8200 ;
        RECT 6.0000 2465.7800 9.0000 2466.2600 ;
        RECT 6.0000 2471.2200 9.0000 2471.7000 ;
        RECT 6.0000 2476.6600 9.0000 2477.1400 ;
        RECT 6.0000 2482.1000 9.0000 2482.5800 ;
        RECT 6.0000 2487.5400 9.0000 2488.0200 ;
        RECT 6.0000 2492.9800 9.0000 2493.4600 ;
        RECT 6.0000 2498.4200 9.0000 2498.9000 ;
        RECT 6.0000 2503.8600 9.0000 2504.3400 ;
        RECT 6.0000 2509.3000 9.0000 2509.7800 ;
        RECT 6.0000 2514.7400 9.0000 2515.2200 ;
        RECT 6.0000 2520.1800 9.0000 2520.6600 ;
        RECT 6.0000 2525.6200 9.0000 2526.1000 ;
        RECT 6.0000 2531.0600 9.0000 2531.5400 ;
        RECT 6.0000 2536.5000 9.0000 2536.9800 ;
        RECT 6.0000 2541.9400 9.0000 2542.4200 ;
        RECT 6.0000 2547.3800 9.0000 2547.8600 ;
        RECT 6.0000 2552.8200 9.0000 2553.3000 ;
        RECT 6.0000 2558.2600 9.0000 2558.7400 ;
        RECT 1002.9200 2128.5000 1004.5200 2128.9800 ;
        RECT 1002.9200 2133.9400 1004.5200 2134.4200 ;
        RECT 1002.9200 2139.3800 1004.5200 2139.8600 ;
        RECT 1002.9200 2144.8200 1004.5200 2145.3000 ;
        RECT 1002.9200 2150.2600 1004.5200 2150.7400 ;
        RECT 1002.9200 2166.5800 1004.5200 2167.0600 ;
        RECT 1002.9200 2161.1400 1004.5200 2161.6200 ;
        RECT 1002.9200 2155.7000 1004.5200 2156.1800 ;
        RECT 1002.9200 2172.0200 1004.5200 2172.5000 ;
        RECT 1002.9200 2177.4600 1004.5200 2177.9400 ;
        RECT 1002.9200 2182.9000 1004.5200 2183.3800 ;
        RECT 1002.9200 2188.3400 1004.5200 2188.8200 ;
        RECT 1002.9200 2193.7800 1004.5200 2194.2600 ;
        RECT 1002.9200 2199.2200 1004.5200 2199.7000 ;
        RECT 1002.9200 2204.6600 1004.5200 2205.1400 ;
        RECT 1002.9200 2210.1000 1004.5200 2210.5800 ;
        RECT 1002.9200 2215.5400 1004.5200 2216.0200 ;
        RECT 1002.9200 2220.9800 1004.5200 2221.4600 ;
        RECT 1002.9200 2226.4200 1004.5200 2226.9000 ;
        RECT 1002.9200 2231.8600 1004.5200 2232.3400 ;
        RECT 1002.9200 2259.0600 1004.5200 2259.5400 ;
        RECT 1002.9200 2237.3000 1004.5200 2237.7800 ;
        RECT 1002.9200 2242.7400 1004.5200 2244.6200 ;
        RECT 1002.9200 2248.1800 1004.5200 2248.6600 ;
        RECT 1002.9200 2264.5000 1004.5200 2264.9800 ;
        RECT 1002.9200 2269.9400 1004.5200 2270.4200 ;
        RECT 1002.9200 2275.3800 1004.5200 2275.8600 ;
        RECT 1002.9200 2280.8200 1004.5200 2281.3000 ;
        RECT 1002.9200 2286.2600 1004.5200 2286.7400 ;
        RECT 1002.9200 2291.7000 1004.5200 2292.1800 ;
        RECT 1002.9200 2297.1400 1004.5200 2297.6200 ;
        RECT 1002.9200 2302.5800 1004.5200 2303.0600 ;
        RECT 1002.9200 2308.0200 1004.5200 2308.5000 ;
        RECT 1002.9200 2318.9000 1004.5200 2319.3800 ;
        RECT 1002.9200 2313.4600 1004.5200 2313.9400 ;
        RECT 1002.9200 2324.3400 1004.5200 2324.8200 ;
        RECT 1002.9200 2329.7800 1004.5200 2330.2600 ;
        RECT 1002.9200 2335.2200 1004.5200 2335.7000 ;
        RECT 1055.6000 2228.7600 1057.2000 2229.2400 ;
        RECT 1055.6000 2262.5600 1057.2000 2263.0400 ;
        RECT 1002.9200 2346.1000 1004.5200 2346.5800 ;
        RECT 1002.9200 2340.6600 1004.5200 2341.1400 ;
        RECT 1002.9200 2351.5400 1004.5200 2352.0200 ;
        RECT 1002.9200 2356.9800 1004.5200 2357.4600 ;
        RECT 1002.9200 2362.4200 1004.5200 2362.9000 ;
        RECT 1002.9200 2367.8600 1004.5200 2368.3400 ;
        RECT 1002.9200 2373.3000 1004.5200 2373.7800 ;
        RECT 1002.9200 2378.7400 1004.5200 2379.2200 ;
        RECT 1002.9200 2384.1800 1004.5200 2384.6600 ;
        RECT 1002.9200 2389.6200 1004.5200 2390.1000 ;
        RECT 1002.9200 2416.8200 1004.5200 2417.3000 ;
        RECT 1002.9200 2400.5000 1004.5200 2400.9800 ;
        RECT 1002.9200 2395.0600 1004.5200 2395.5400 ;
        RECT 1002.9200 2405.9400 1004.5200 2406.4200 ;
        RECT 1002.9200 2411.3800 1004.5200 2411.8600 ;
        RECT 1002.9200 2427.7000 1004.5200 2428.1800 ;
        RECT 1002.9200 2422.2600 1004.5200 2422.7400 ;
        RECT 1002.9200 2433.1400 1004.5200 2433.6200 ;
        RECT 1002.9200 2438.5800 1004.5200 2439.0600 ;
        RECT 1002.9200 2444.0200 1004.5200 2444.5000 ;
        RECT 1002.9200 2449.4600 1004.5200 2449.9400 ;
        RECT 1002.9200 2454.9000 1004.5200 2455.3800 ;
        RECT 1002.9200 2460.3400 1004.5200 2460.8200 ;
        RECT 1002.9200 2464.6500 1004.5200 2466.2600 ;
        RECT 1013.1800 2482.1000 1014.7800 2482.5800 ;
        RECT 1002.9200 2482.1000 1004.5200 2482.5800 ;
        RECT 1002.9200 2476.6600 1004.5200 2477.1400 ;
        RECT 1002.9200 2471.2200 1004.5200 2471.7000 ;
        RECT 1013.1800 2487.5400 1014.7800 2488.0200 ;
        RECT 1013.1800 2492.9800 1014.7800 2493.4600 ;
        RECT 1002.9200 2492.9800 1004.5200 2493.4600 ;
        RECT 1002.9200 2487.5400 1004.5200 2488.0200 ;
        RECT 1013.1800 2498.4200 1014.7800 2498.9000 ;
        RECT 1013.1800 2503.8600 1014.7800 2504.3400 ;
        RECT 1002.9200 2503.8600 1004.5200 2504.3400 ;
        RECT 1002.9200 2498.4200 1004.5200 2498.9000 ;
        RECT 1013.1800 2509.3000 1014.7800 2509.7800 ;
        RECT 1013.1800 2514.7400 1014.7800 2515.2200 ;
        RECT 1013.1800 2520.1800 1014.7800 2520.6600 ;
        RECT 1002.9200 2509.3000 1004.5200 2509.7800 ;
        RECT 1002.9200 2514.7400 1004.5200 2515.2200 ;
        RECT 1002.9200 2520.1800 1004.5200 2520.6600 ;
        RECT 1013.1800 2525.6200 1014.7800 2526.1000 ;
        RECT 1013.1800 2531.0600 1014.7800 2531.5400 ;
        RECT 1002.9200 2525.6200 1004.5200 2526.1000 ;
        RECT 1002.9200 2531.0600 1004.5200 2531.5400 ;
        RECT 1013.1800 2536.5000 1014.7800 2536.9800 ;
        RECT 1013.1800 2541.9400 1014.7800 2542.4200 ;
        RECT 1013.1800 2547.3800 1014.7800 2547.8600 ;
        RECT 1002.9200 2536.5000 1004.5200 2536.9800 ;
        RECT 1002.9200 2541.9400 1004.5200 2542.4200 ;
        RECT 1002.9200 2547.3800 1004.5200 2547.8600 ;
        RECT 1060.5600 2464.6500 1062.1600 2466.2500 ;
        RECT 1073.2200 2457.2400 1074.8200 2457.7200 ;
        RECT 1055.6000 2482.1000 1057.2000 2482.5800 ;
        RECT 1065.8600 2487.5400 1067.4600 2488.0200 ;
        RECT 1065.8600 2492.9800 1067.4600 2493.4600 ;
        RECT 1055.6000 2492.9800 1057.2000 2493.4600 ;
        RECT 1055.6000 2487.5400 1057.2000 2488.0200 ;
        RECT 1073.1800 2489.2200 1074.7800 2489.7000 ;
        RECT 1065.8600 2498.4200 1067.4600 2498.9000 ;
        RECT 1065.8600 2505.0500 1067.4600 2507.1000 ;
        RECT 1055.6000 2498.4200 1057.2000 2498.9000 ;
        RECT 1055.6000 2503.8600 1057.2000 2504.3400 ;
        RECT 1065.8600 2509.3000 1067.4600 2509.7800 ;
        RECT 1065.8600 2514.7400 1067.4600 2515.2200 ;
        RECT 1065.8600 2520.1800 1067.4600 2520.6600 ;
        RECT 1055.6000 2509.3000 1057.2000 2509.7800 ;
        RECT 1055.6000 2514.7400 1057.2000 2515.2200 ;
        RECT 1055.6000 2520.1800 1057.2000 2520.6600 ;
        RECT 1073.1800 2520.1800 1074.7800 2520.6600 ;
        RECT 1065.8600 2525.6200 1067.4600 2526.1000 ;
        RECT 1065.8600 2531.0600 1067.4600 2531.5400 ;
        RECT 1055.6000 2525.6200 1057.2000 2526.1000 ;
        RECT 1055.6000 2531.0600 1057.2000 2531.5400 ;
        RECT 1073.1800 2525.6200 1074.7800 2526.1000 ;
        RECT 1073.1800 2531.0600 1074.7800 2531.5400 ;
        RECT 1065.8600 2536.5000 1067.4600 2536.9800 ;
        RECT 1065.8600 2541.9400 1067.4600 2542.4200 ;
        RECT 1065.8600 2547.3800 1067.4600 2547.8600 ;
        RECT 1055.6000 2536.5000 1057.2000 2536.9800 ;
        RECT 1055.6000 2541.9400 1057.2000 2542.4200 ;
        RECT 1055.6000 2547.3800 1057.2000 2547.8600 ;
        RECT 1073.1800 2536.5000 1074.7800 2536.9800 ;
        RECT 1073.1800 2541.9400 1074.7800 2542.4200 ;
        RECT 1073.1800 2547.3800 1074.7800 2547.8600 ;
        RECT 1293.3000 2228.5000 1294.9000 2228.9800 ;
        RECT 1513.5200 2228.5000 1515.1200 2228.9800 ;
        RECT 1285.9400 2464.4900 1287.6800 2467.4000 ;
        RECT 1300.4600 2458.1400 1302.0600 2458.6200 ;
        RECT 1293.4000 2489.2200 1295.0000 2489.7000 ;
        RECT 1275.6800 2520.1800 1277.2800 2520.6600 ;
        RECT 1285.9400 2520.1800 1287.6800 2520.6600 ;
        RECT 1293.4000 2520.1800 1295.0000 2520.6600 ;
        RECT 1275.6800 2525.6200 1277.2800 2526.1000 ;
        RECT 1275.6800 2531.0600 1277.2800 2531.5400 ;
        RECT 1285.9400 2525.6200 1287.6800 2526.1000 ;
        RECT 1285.9400 2531.0600 1287.6800 2531.5400 ;
        RECT 1275.6800 2536.5000 1277.2800 2536.9800 ;
        RECT 1275.6800 2541.9400 1277.2800 2542.4200 ;
        RECT 1275.6800 2547.3800 1277.2800 2547.8600 ;
        RECT 1285.9400 2536.5000 1287.6800 2536.9800 ;
        RECT 1285.9400 2541.9400 1287.6800 2542.4200 ;
        RECT 1285.9400 2547.3800 1287.6800 2547.8600 ;
        RECT 1293.4000 2525.6200 1295.0000 2526.1000 ;
        RECT 1293.4000 2531.0600 1295.0000 2531.5400 ;
        RECT 1293.4000 2536.5000 1295.0000 2536.9800 ;
        RECT 1293.4000 2541.9400 1295.0000 2542.4200 ;
        RECT 1293.4000 2547.3800 1295.0000 2547.8600 ;
        RECT 1520.6800 2458.1400 1522.2800 2458.6200 ;
        RECT 1513.6200 2489.2200 1515.2200 2489.7000 ;
        RECT 1495.9000 2520.1800 1497.5000 2520.6600 ;
        RECT 1506.1600 2520.1800 1507.7600 2520.6600 ;
        RECT 1513.6200 2520.1800 1515.2200 2520.6600 ;
        RECT 1495.9000 2525.6200 1497.5000 2526.1000 ;
        RECT 1495.9000 2531.0600 1497.5000 2531.5400 ;
        RECT 1495.9000 2536.5000 1497.5000 2536.9800 ;
        RECT 1495.9000 2541.9400 1497.5000 2542.4200 ;
        RECT 1495.9000 2547.3800 1497.5000 2547.8600 ;
        RECT 1513.6200 2525.6200 1515.2200 2526.1000 ;
        RECT 1513.6200 2531.0600 1515.2200 2531.5400 ;
        RECT 1506.1600 2525.6200 1507.7600 2526.1000 ;
        RECT 1506.1600 2531.0600 1507.7600 2531.5400 ;
        RECT 1513.6200 2536.5000 1515.2200 2536.9800 ;
        RECT 1513.6200 2541.9400 1515.2200 2542.4200 ;
        RECT 1513.6200 2547.3800 1515.2200 2547.8600 ;
        RECT 1506.1600 2536.5000 1507.7600 2536.9800 ;
        RECT 1506.1600 2541.9400 1507.7600 2542.4200 ;
        RECT 1506.1600 2547.3800 1507.7600 2547.8600 ;
        RECT 1013.1800 2552.8200 1014.7800 2553.3000 ;
        RECT 1013.1800 2558.2600 1014.7800 2558.7400 ;
        RECT 1002.9200 2552.8200 1004.5200 2553.3000 ;
        RECT 1002.9200 2558.2600 1004.5200 2558.7400 ;
        RECT 1065.8600 2552.8200 1067.4600 2553.3000 ;
        RECT 1065.8600 2558.2600 1067.4600 2558.7400 ;
        RECT 1055.6000 2552.8200 1057.2000 2553.3000 ;
        RECT 1055.6000 2558.2600 1057.2000 2558.7400 ;
        RECT 1073.1800 2552.8200 1074.7800 2553.3000 ;
        RECT 1073.1800 2558.2600 1074.7800 2558.7400 ;
        RECT 1275.6800 2552.8200 1277.2800 2553.3000 ;
        RECT 1275.6800 2558.2600 1277.2800 2558.7400 ;
        RECT 1285.9400 2552.8200 1287.6800 2553.3000 ;
        RECT 1285.9400 2558.2600 1287.6800 2558.7400 ;
        RECT 1293.4000 2552.8200 1295.0000 2553.3000 ;
        RECT 1293.4000 2558.2600 1295.0000 2558.7400 ;
        RECT 1495.9000 2552.8200 1497.5000 2553.3000 ;
        RECT 1495.9000 2558.2600 1497.5000 2558.7400 ;
        RECT 1513.6200 2552.8200 1515.2200 2553.3000 ;
        RECT 1513.6200 2558.2600 1515.2200 2558.7400 ;
        RECT 1506.1600 2558.2600 1507.7600 2558.7400 ;
        RECT 1506.1600 2552.8200 1507.7600 2553.3000 ;
        RECT 1733.7400 1309.9400 1735.3400 1310.4200 ;
        RECT 1733.7400 1539.5800 1735.3400 1540.0600 ;
        RECT 1941.3000 1545.9300 1942.9000 1547.5300 ;
        RECT 1953.9600 1538.4200 1955.5600 1538.9000 ;
        RECT 2174.1800 1309.9400 2175.7800 1310.4200 ;
        RECT 2394.4000 1309.9400 2396.0000 1310.4200 ;
        RECT 2166.8200 1545.9300 2168.4200 1548.5800 ;
        RECT 2174.1800 1539.5800 2175.7800 1540.0600 ;
        RECT 2394.4000 1539.5800 2396.0000 1540.0600 ;
        RECT 1733.7400 1769.2200 1735.3400 1769.7000 ;
        RECT 1733.7400 1998.8600 1735.3400 1999.3400 ;
        RECT 1941.3000 2005.2100 1942.9000 2006.8100 ;
        RECT 1953.9600 1997.7000 1955.5600 1998.1800 ;
        RECT 2174.1800 1769.2200 2175.7800 1769.7000 ;
        RECT 2394.4000 1769.2200 2396.0000 1769.7000 ;
        RECT 2166.8200 2005.2100 2168.4200 2007.8600 ;
        RECT 2174.1800 1998.8600 2175.7800 1999.3400 ;
        RECT 2394.4000 1998.8600 2396.0000 1999.3400 ;
        RECT 2447.1800 1970.7400 2448.7800 1971.2200 ;
        RECT 2447.1800 1976.1800 2448.7800 1976.6600 ;
        RECT 2447.1800 1981.6200 2448.7800 1982.1000 ;
        RECT 2447.1800 1987.0600 2448.7800 1987.5400 ;
        RECT 2447.1800 1992.5000 2448.7800 1992.9800 ;
        RECT 2447.1800 2008.8200 2448.7800 2009.3000 ;
        RECT 2447.1800 1997.9400 2448.7800 1998.4200 ;
        RECT 2447.1800 2003.3800 2448.7800 2003.8600 ;
        RECT 2447.1800 2013.1200 2448.7800 2014.7400 ;
        RECT 2447.1800 2019.7000 2448.7800 2020.1800 ;
        RECT 2492.9200 1970.7400 2494.5200 1971.2200 ;
        RECT 2492.9200 1976.1800 2494.5200 1976.6600 ;
        RECT 2492.9200 1981.6200 2494.5200 1982.1000 ;
        RECT 2492.9200 1987.0600 2494.5200 1987.5400 ;
        RECT 2492.9200 1992.5000 2494.5200 1992.9800 ;
        RECT 2492.9200 2008.8200 2494.5200 2009.3000 ;
        RECT 2492.9200 2003.3800 2494.5200 2003.8600 ;
        RECT 2492.9200 1997.9400 2494.5200 1998.4200 ;
        RECT 2492.9200 2014.2600 2494.5200 2014.7400 ;
        RECT 2492.9200 2019.7000 2494.5200 2020.1800 ;
        RECT 2447.1800 2025.1400 2448.7800 2025.6200 ;
        RECT 2447.1800 2030.5800 2448.7800 2031.0600 ;
        RECT 2447.1800 2036.0200 2448.7800 2036.5000 ;
        RECT 2447.1800 2041.4600 2448.7800 2041.9400 ;
        RECT 2447.1800 2046.9000 2448.7800 2047.3800 ;
        RECT 2447.1800 2052.3400 2448.7800 2052.8200 ;
        RECT 2447.1800 2057.7800 2448.7800 2058.2600 ;
        RECT 2447.1800 2063.2200 2448.7800 2063.7000 ;
        RECT 2447.1800 2068.6600 2448.7800 2069.1400 ;
        RECT 2447.1800 2074.1000 2448.7800 2074.5800 ;
        RECT 2492.9200 2025.1400 2494.5200 2025.6200 ;
        RECT 2492.9200 2030.5800 2494.5200 2031.0600 ;
        RECT 2492.9200 2036.0200 2494.5200 2036.5000 ;
        RECT 2492.9200 2041.4600 2494.5200 2041.9400 ;
        RECT 2492.9200 2046.9000 2494.5200 2047.3800 ;
        RECT 2492.9200 2052.3400 2494.5200 2052.8200 ;
        RECT 2492.9200 2057.7800 2494.5200 2058.2600 ;
        RECT 2492.9200 2063.2200 2494.5200 2063.7000 ;
        RECT 2492.9200 2068.6600 2494.5200 2069.1400 ;
        RECT 2492.9200 2074.1000 2494.5200 2074.5800 ;
        RECT 2447.1800 2079.5400 2448.7800 2080.0200 ;
        RECT 2447.1800 2084.9800 2448.7800 2085.4600 ;
        RECT 2447.1800 2090.4200 2448.7800 2090.9000 ;
        RECT 2447.1800 2095.8600 2448.7800 2096.3400 ;
        RECT 2447.1800 2101.3000 2448.7800 2101.7800 ;
        RECT 2447.1800 2106.7400 2448.7800 2107.2200 ;
        RECT 2447.1800 2112.1800 2448.7800 2112.6600 ;
        RECT 2447.1800 2117.6200 2448.7800 2118.1000 ;
        RECT 2447.1800 2123.0600 2448.7800 2123.5400 ;
        RECT 2492.9200 2084.9800 2494.5200 2085.4600 ;
        RECT 2492.9200 2079.5400 2494.5200 2080.0200 ;
        RECT 2492.9200 2090.4200 2494.5200 2090.9000 ;
        RECT 2492.9200 2095.8600 2494.5200 2096.3400 ;
        RECT 2492.9200 2101.3000 2494.5200 2101.7800 ;
        RECT 2492.9200 2106.7400 2494.5200 2107.2200 ;
        RECT 2492.9200 2112.1800 2494.5200 2112.6600 ;
        RECT 2492.9200 2117.6200 2494.5200 2118.1000 ;
        RECT 2492.9200 2123.0600 2494.5200 2123.5400 ;
        RECT 3305.7200 1285.3000 3307.3200 1285.7800 ;
        RECT 3305.7200 1290.7400 3307.3200 1291.2200 ;
        RECT 3305.7200 1296.1800 3307.3200 1296.6600 ;
        RECT 3305.7200 1301.6200 3307.3200 1302.1000 ;
        RECT 3305.7200 1307.0600 3307.3200 1307.5400 ;
        RECT 3305.7200 1312.5000 3307.3200 1312.9800 ;
        RECT 3305.7200 1317.9400 3307.3200 1318.4200 ;
        RECT 3305.7200 1323.3800 3307.3200 1323.8600 ;
        RECT 3305.7200 1328.8200 3307.3200 1329.3000 ;
        RECT 3305.7200 1334.2600 3307.3200 1334.7400 ;
        RECT 3361.4200 1285.3000 3364.4200 1285.7800 ;
        RECT 3361.4200 1290.7400 3364.4200 1291.2200 ;
        RECT 3361.4200 1296.1800 3364.4200 1296.6600 ;
        RECT 3361.4200 1301.6200 3364.4200 1302.1000 ;
        RECT 3361.4200 1307.0600 3364.4200 1307.5400 ;
        RECT 3361.4200 1312.5000 3364.4200 1312.9800 ;
        RECT 3361.4200 1317.9400 3364.4200 1318.4200 ;
        RECT 3361.4200 1323.3800 3364.4200 1323.8600 ;
        RECT 3361.4200 1328.8200 3364.4200 1329.3000 ;
        RECT 3361.4200 1334.2600 3364.4200 1334.7400 ;
        RECT 3305.7200 1350.5800 3307.3200 1351.0600 ;
        RECT 3305.7200 1339.7000 3307.3200 1340.1800 ;
        RECT 3305.7200 1345.1400 3307.3200 1345.6200 ;
        RECT 3305.7200 1356.0200 3307.3200 1356.5000 ;
        RECT 3305.7200 1361.4600 3307.3200 1361.9400 ;
        RECT 3305.7200 1366.9000 3307.3200 1367.3800 ;
        RECT 3305.7200 1372.3400 3307.3200 1372.8200 ;
        RECT 3305.7200 1377.7800 3307.3200 1378.2600 ;
        RECT 3305.7200 1383.2200 3307.3200 1383.7000 ;
        RECT 3305.7200 1388.6600 3307.3200 1389.1400 ;
        RECT 3361.4200 1350.5800 3364.4200 1351.0600 ;
        RECT 3361.4200 1339.7000 3364.4200 1340.1800 ;
        RECT 3361.4200 1345.1400 3364.4200 1345.6200 ;
        RECT 3361.4200 1356.0200 3364.4200 1356.5000 ;
        RECT 3361.4200 1361.4600 3364.4200 1361.9400 ;
        RECT 3361.4200 1366.9000 3364.4200 1367.3800 ;
        RECT 3361.4200 1372.3400 3364.4200 1372.8200 ;
        RECT 3361.4200 1377.7800 3364.4200 1378.2600 ;
        RECT 3361.4200 1383.2200 3364.4200 1383.7000 ;
        RECT 3361.4200 1388.6600 3364.4200 1389.1400 ;
        RECT 3305.7200 1394.1000 3307.3200 1394.5800 ;
        RECT 3305.7200 1399.5400 3307.3200 1400.0200 ;
        RECT 3305.7200 1404.9800 3307.3200 1405.4600 ;
        RECT 3305.7200 1410.4200 3307.3200 1410.9000 ;
        RECT 3305.7200 1415.8600 3307.3200 1416.3400 ;
        RECT 3305.7200 1421.3000 3307.3200 1421.7800 ;
        RECT 3305.7200 1426.7400 3307.3200 1427.2200 ;
        RECT 3305.7200 1432.1800 3307.3200 1432.6600 ;
        RECT 3305.7200 1437.6200 3307.3200 1438.1000 ;
        RECT 3361.4200 1394.1000 3364.4200 1394.5800 ;
        RECT 3361.4200 1399.5400 3364.4200 1400.0200 ;
        RECT 3361.4200 1404.9800 3364.4200 1405.4600 ;
        RECT 3361.4200 1410.4200 3364.4200 1410.9000 ;
        RECT 3361.4200 1415.8600 3364.4200 1416.3400 ;
        RECT 3361.4200 1421.3000 3364.4200 1421.7800 ;
        RECT 3361.4200 1426.7400 3364.4200 1427.2200 ;
        RECT 3361.4200 1432.1800 3364.4200 1432.6600 ;
        RECT 3361.4200 1437.6200 3364.4200 1438.1000 ;
        RECT 3305.7200 1443.0600 3307.3200 1443.5400 ;
        RECT 3305.7200 1448.5000 3307.3200 1448.9800 ;
        RECT 3305.7200 1453.9400 3307.3200 1454.4200 ;
        RECT 3305.7200 1459.3800 3307.3200 1459.8600 ;
        RECT 3305.7200 1464.8200 3307.3200 1465.3000 ;
        RECT 3305.7200 1470.2600 3307.3200 1470.7400 ;
        RECT 3305.7200 1475.7000 3307.3200 1476.1800 ;
        RECT 3305.7200 1481.1400 3307.3200 1481.6200 ;
        RECT 3305.7200 1486.5800 3307.3200 1487.0600 ;
        RECT 3305.7200 1492.0200 3307.3200 1492.5000 ;
        RECT 3361.4200 1443.0600 3364.4200 1443.5400 ;
        RECT 3361.4200 1448.5000 3364.4200 1448.9800 ;
        RECT 3361.4200 1453.9400 3364.4200 1454.4200 ;
        RECT 3361.4200 1459.3800 3364.4200 1459.8600 ;
        RECT 3361.4200 1464.8200 3364.4200 1465.3000 ;
        RECT 3361.4200 1470.2600 3364.4200 1470.7400 ;
        RECT 3361.4200 1475.7000 3364.4200 1476.1800 ;
        RECT 3361.4200 1481.1400 3364.4200 1481.6200 ;
        RECT 3361.4200 1486.5800 3364.4200 1487.0600 ;
        RECT 3361.4200 1492.0200 3364.4200 1492.5000 ;
        RECT 3361.4200 1600.8200 3364.4200 1601.3000 ;
        RECT 3305.7200 1600.8200 3307.3200 1601.3000 ;
        RECT 3305.7200 1508.3400 3307.3200 1508.8200 ;
        RECT 3305.7200 1497.4600 3307.3200 1497.9400 ;
        RECT 3305.7200 1502.9000 3307.3200 1503.3800 ;
        RECT 3305.7200 1513.7800 3307.3200 1514.2600 ;
        RECT 3305.7200 1519.2200 3307.3200 1519.7000 ;
        RECT 3305.7200 1524.6600 3307.3200 1525.1400 ;
        RECT 3305.7200 1530.1000 3307.3200 1530.5800 ;
        RECT 3305.7200 1535.5400 3307.3200 1536.0200 ;
        RECT 3305.7200 1540.9800 3307.3200 1541.4600 ;
        RECT 3305.7200 1546.4200 3307.3200 1546.9000 ;
        RECT 3361.4200 1508.3400 3364.4200 1508.8200 ;
        RECT 3361.4200 1497.4600 3364.4200 1497.9400 ;
        RECT 3361.4200 1502.9000 3364.4200 1503.3800 ;
        RECT 3361.4200 1513.7800 3364.4200 1514.2600 ;
        RECT 3361.4200 1519.2200 3364.4200 1519.7000 ;
        RECT 3361.4200 1524.6600 3364.4200 1525.1400 ;
        RECT 3361.4200 1530.1000 3364.4200 1530.5800 ;
        RECT 3361.4200 1535.5400 3364.4200 1536.0200 ;
        RECT 3361.4200 1540.9800 3364.4200 1541.4600 ;
        RECT 3361.4200 1546.4200 3364.4200 1546.9000 ;
        RECT 3305.7200 1551.8600 3307.3200 1552.3400 ;
        RECT 3305.7200 1557.3000 3307.3200 1557.7800 ;
        RECT 3305.7200 1562.7400 3307.3200 1563.2200 ;
        RECT 3305.7200 1568.1800 3307.3200 1568.6600 ;
        RECT 3305.7200 1573.6200 3307.3200 1574.1000 ;
        RECT 3305.7200 1579.0600 3307.3200 1579.5400 ;
        RECT 3305.7200 1584.5000 3307.3200 1584.9800 ;
        RECT 3305.7200 1589.9400 3307.3200 1590.4200 ;
        RECT 3305.7200 1595.3800 3307.3200 1595.8600 ;
        RECT 3361.4200 1551.8600 3364.4200 1552.3400 ;
        RECT 3361.4200 1557.3000 3364.4200 1557.7800 ;
        RECT 3361.4200 1562.7400 3364.4200 1563.2200 ;
        RECT 3361.4200 1568.1800 3364.4200 1568.6600 ;
        RECT 3361.4200 1573.6200 3364.4200 1574.1000 ;
        RECT 3361.4200 1579.0600 3364.4200 1579.5400 ;
        RECT 3361.4200 1584.5000 3364.4200 1584.9800 ;
        RECT 3361.4200 1589.9400 3364.4200 1590.4200 ;
        RECT 3361.4200 1595.3800 3364.4200 1595.8600 ;
        RECT 3305.7200 1606.2600 3307.3200 1606.7400 ;
        RECT 3305.7200 1611.7000 3307.3200 1612.1800 ;
        RECT 3305.7200 1617.1400 3307.3200 1617.6200 ;
        RECT 3305.7200 1622.5800 3307.3200 1623.0600 ;
        RECT 3305.7200 1628.0200 3307.3200 1628.5000 ;
        RECT 3305.7200 1633.4600 3307.3200 1633.9400 ;
        RECT 3305.7200 1638.9000 3307.3200 1639.3800 ;
        RECT 3305.7200 1644.3400 3307.3200 1644.8200 ;
        RECT 3305.7200 1649.7800 3307.3200 1650.2600 ;
        RECT 3361.4200 1606.2600 3364.4200 1606.7400 ;
        RECT 3361.4200 1611.7000 3364.4200 1612.1800 ;
        RECT 3361.4200 1617.1400 3364.4200 1617.6200 ;
        RECT 3361.4200 1622.5800 3364.4200 1623.0600 ;
        RECT 3361.4200 1628.0200 3364.4200 1628.5000 ;
        RECT 3361.4200 1633.4600 3364.4200 1633.9400 ;
        RECT 3361.4200 1638.9000 3364.4200 1639.3800 ;
        RECT 3361.4200 1644.3400 3364.4200 1644.8200 ;
        RECT 3361.4200 1649.7800 3364.4200 1650.2600 ;
        RECT 3305.7200 1655.2200 3307.3200 1655.7000 ;
        RECT 3305.7200 1660.6600 3307.3200 1661.1400 ;
        RECT 3305.7200 1666.1000 3307.3200 1666.5800 ;
        RECT 3305.7200 1671.5400 3307.3200 1672.0200 ;
        RECT 3305.7200 1676.9800 3307.3200 1677.4600 ;
        RECT 3305.7200 1682.4200 3307.3200 1682.9000 ;
        RECT 3305.7200 1687.8600 3307.3200 1688.3400 ;
        RECT 3305.7200 1693.3000 3307.3200 1693.7800 ;
        RECT 3305.7200 1698.7400 3307.3200 1699.2200 ;
        RECT 3305.7200 1704.1800 3307.3200 1704.6600 ;
        RECT 3361.4200 1655.2200 3364.4200 1655.7000 ;
        RECT 3361.4200 1660.6600 3364.4200 1661.1400 ;
        RECT 3361.4200 1666.1000 3364.4200 1666.5800 ;
        RECT 3361.4200 1671.5400 3364.4200 1672.0200 ;
        RECT 3361.4200 1676.9800 3364.4200 1677.4600 ;
        RECT 3361.4200 1682.4200 3364.4200 1682.9000 ;
        RECT 3361.4200 1687.8600 3364.4200 1688.3400 ;
        RECT 3361.4200 1693.3000 3364.4200 1693.7800 ;
        RECT 3361.4200 1698.7400 3364.4200 1699.2200 ;
        RECT 3361.4200 1704.1800 3364.4200 1704.6600 ;
        RECT 3361.4200 1916.3400 3364.4200 1916.8200 ;
        RECT 3305.7200 1916.3400 3307.3200 1916.8200 ;
        RECT 3361.4200 1758.5800 3364.4200 1759.0600 ;
        RECT 3305.7200 1758.5800 3307.3200 1759.0600 ;
        RECT 3305.7200 1709.6200 3307.3200 1710.1000 ;
        RECT 3305.7200 1715.0600 3307.3200 1715.5400 ;
        RECT 3305.7200 1720.5000 3307.3200 1720.9800 ;
        RECT 3305.7200 1725.9400 3307.3200 1726.4200 ;
        RECT 3305.7200 1731.3800 3307.3200 1731.8600 ;
        RECT 3305.7200 1736.8200 3307.3200 1737.3000 ;
        RECT 3305.7200 1742.2600 3307.3200 1742.7400 ;
        RECT 3305.7200 1747.7000 3307.3200 1748.1800 ;
        RECT 3305.7200 1753.1400 3307.3200 1753.6200 ;
        RECT 3361.4200 1709.6200 3364.4200 1710.1000 ;
        RECT 3361.4200 1715.0600 3364.4200 1715.5400 ;
        RECT 3361.4200 1720.5000 3364.4200 1720.9800 ;
        RECT 3361.4200 1725.9400 3364.4200 1726.4200 ;
        RECT 3361.4200 1731.3800 3364.4200 1731.8600 ;
        RECT 3361.4200 1736.8200 3364.4200 1737.3000 ;
        RECT 3361.4200 1742.2600 3364.4200 1742.7400 ;
        RECT 3361.4200 1747.7000 3364.4200 1748.1800 ;
        RECT 3361.4200 1753.1400 3364.4200 1753.6200 ;
        RECT 3305.7200 1764.0200 3307.3200 1764.5000 ;
        RECT 3305.7200 1769.4600 3307.3200 1769.9400 ;
        RECT 3305.7200 1774.9000 3307.3200 1775.3800 ;
        RECT 3305.7200 1780.3400 3307.3200 1780.8200 ;
        RECT 3305.7200 1785.7800 3307.3200 1786.2600 ;
        RECT 3305.7200 1791.2200 3307.3200 1791.7000 ;
        RECT 3305.7200 1796.6600 3307.3200 1797.1400 ;
        RECT 3305.7200 1802.1000 3307.3200 1802.5800 ;
        RECT 3305.7200 1807.5400 3307.3200 1808.0200 ;
        RECT 3361.4200 1764.0200 3364.4200 1764.5000 ;
        RECT 3361.4200 1769.4600 3364.4200 1769.9400 ;
        RECT 3361.4200 1774.9000 3364.4200 1775.3800 ;
        RECT 3361.4200 1780.3400 3364.4200 1780.8200 ;
        RECT 3361.4200 1785.7800 3364.4200 1786.2600 ;
        RECT 3361.4200 1791.2200 3364.4200 1791.7000 ;
        RECT 3361.4200 1796.6600 3364.4200 1797.1400 ;
        RECT 3361.4200 1802.1000 3364.4200 1802.5800 ;
        RECT 3361.4200 1807.5400 3364.4200 1808.0200 ;
        RECT 3305.7200 1812.9800 3307.3200 1813.4600 ;
        RECT 3305.7200 1818.4200 3307.3200 1818.9000 ;
        RECT 3305.7200 1823.8600 3307.3200 1824.3400 ;
        RECT 3305.7200 1829.3000 3307.3200 1829.7800 ;
        RECT 3305.7200 1834.7400 3307.3200 1835.2200 ;
        RECT 3305.7200 1840.1800 3307.3200 1840.6600 ;
        RECT 3305.7200 1845.6200 3307.3200 1846.1000 ;
        RECT 3305.7200 1851.0600 3307.3200 1851.5400 ;
        RECT 3305.7200 1856.5000 3307.3200 1856.9800 ;
        RECT 3305.7200 1861.9400 3307.3200 1862.4200 ;
        RECT 3361.4200 1812.9800 3364.4200 1813.4600 ;
        RECT 3361.4200 1818.4200 3364.4200 1818.9000 ;
        RECT 3361.4200 1823.8600 3364.4200 1824.3400 ;
        RECT 3361.4200 1829.3000 3364.4200 1829.7800 ;
        RECT 3361.4200 1834.7400 3364.4200 1835.2200 ;
        RECT 3361.4200 1840.1800 3364.4200 1840.6600 ;
        RECT 3361.4200 1845.6200 3364.4200 1846.1000 ;
        RECT 3361.4200 1851.0600 3364.4200 1851.5400 ;
        RECT 3361.4200 1856.5000 3364.4200 1856.9800 ;
        RECT 3361.4200 1861.9400 3364.4200 1862.4200 ;
        RECT 3305.7200 1867.3800 3307.3200 1867.8600 ;
        RECT 3305.7200 1872.8200 3307.3200 1873.3000 ;
        RECT 3305.7200 1878.2600 3307.3200 1878.7400 ;
        RECT 3305.7200 1883.7000 3307.3200 1884.1800 ;
        RECT 3305.7200 1889.1400 3307.3200 1889.6200 ;
        RECT 3305.7200 1894.5800 3307.3200 1895.0600 ;
        RECT 3305.7200 1900.0200 3307.3200 1900.5000 ;
        RECT 3305.7200 1905.4600 3307.3200 1905.9400 ;
        RECT 3305.7200 1910.9000 3307.3200 1911.3800 ;
        RECT 3361.4200 1867.3800 3364.4200 1867.8600 ;
        RECT 3361.4200 1872.8200 3364.4200 1873.3000 ;
        RECT 3361.4200 1878.2600 3364.4200 1878.7400 ;
        RECT 3361.4200 1883.7000 3364.4200 1884.1800 ;
        RECT 3361.4200 1889.1400 3364.4200 1889.6200 ;
        RECT 3361.4200 1894.5800 3364.4200 1895.0600 ;
        RECT 3361.4200 1900.0200 3364.4200 1900.5000 ;
        RECT 3361.4200 1905.4600 3364.4200 1905.9400 ;
        RECT 3361.4200 1910.9000 3364.4200 1911.3800 ;
        RECT 3305.7200 1921.7800 3307.3200 1922.2600 ;
        RECT 3305.7200 1927.2200 3307.3200 1927.7000 ;
        RECT 3305.7200 1932.6600 3307.3200 1933.1400 ;
        RECT 3305.7200 1938.1000 3307.3200 1938.5800 ;
        RECT 3305.7200 1943.5400 3307.3200 1944.0200 ;
        RECT 3305.7200 1948.9800 3307.3200 1949.4600 ;
        RECT 3305.7200 1954.4200 3307.3200 1954.9000 ;
        RECT 3305.7200 1959.8600 3307.3200 1960.3400 ;
        RECT 3305.7200 1965.3000 3307.3200 1965.7800 ;
        RECT 3361.4200 1921.7800 3364.4200 1922.2600 ;
        RECT 3361.4200 1927.2200 3364.4200 1927.7000 ;
        RECT 3361.4200 1932.6600 3364.4200 1933.1400 ;
        RECT 3361.4200 1938.1000 3364.4200 1938.5800 ;
        RECT 3361.4200 1943.5400 3364.4200 1944.0200 ;
        RECT 3361.4200 1948.9800 3364.4200 1949.4600 ;
        RECT 3361.4200 1954.4200 3364.4200 1954.9000 ;
        RECT 3361.4200 1959.8600 3364.4200 1960.3400 ;
        RECT 3361.4200 1965.3000 3364.4200 1965.7800 ;
        RECT 3305.7200 1970.7400 3307.3200 1971.2200 ;
        RECT 3305.7200 1976.1800 3307.3200 1976.6600 ;
        RECT 3305.7200 1981.6200 3307.3200 1982.1000 ;
        RECT 3305.7200 1987.0600 3307.3200 1987.5400 ;
        RECT 3305.7200 1992.5000 3307.3200 1992.9800 ;
        RECT 3305.7200 2008.8200 3307.3200 2009.3000 ;
        RECT 3305.7200 2003.3800 3307.3200 2003.8600 ;
        RECT 3305.7200 1997.9400 3307.3200 1998.4200 ;
        RECT 3305.7200 2014.2600 3307.3200 2014.7400 ;
        RECT 3305.7200 2019.7000 3307.3200 2020.1800 ;
        RECT 3361.4200 1970.7400 3364.4200 1971.2200 ;
        RECT 3361.4200 1976.1800 3364.4200 1976.6600 ;
        RECT 3361.4200 1981.6200 3364.4200 1982.1000 ;
        RECT 3361.4200 1987.0600 3364.4200 1987.5400 ;
        RECT 3361.4200 1992.5000 3364.4200 1992.9800 ;
        RECT 3361.4200 2008.8200 3364.4200 2009.3000 ;
        RECT 3361.4200 1997.9400 3364.4200 1998.4200 ;
        RECT 3361.4200 2003.3800 3364.4200 2003.8600 ;
        RECT 3361.4200 2014.2600 3364.4200 2014.7400 ;
        RECT 3361.4200 2019.7000 3364.4200 2020.1800 ;
        RECT 3305.7200 2025.1400 3307.3200 2025.6200 ;
        RECT 3305.7200 2030.5800 3307.3200 2031.0600 ;
        RECT 3305.7200 2036.0200 3307.3200 2036.5000 ;
        RECT 3305.7200 2041.4600 3307.3200 2041.9400 ;
        RECT 3305.7200 2046.9000 3307.3200 2047.3800 ;
        RECT 3305.7200 2052.3400 3307.3200 2052.8200 ;
        RECT 3305.7200 2057.7800 3307.3200 2058.2600 ;
        RECT 3305.7200 2063.2200 3307.3200 2063.7000 ;
        RECT 3305.7200 2068.6600 3307.3200 2069.1400 ;
        RECT 3305.7200 2074.1000 3307.3200 2074.5800 ;
        RECT 3361.4200 2025.1400 3364.4200 2025.6200 ;
        RECT 3361.4200 2030.5800 3364.4200 2031.0600 ;
        RECT 3361.4200 2036.0200 3364.4200 2036.5000 ;
        RECT 3361.4200 2041.4600 3364.4200 2041.9400 ;
        RECT 3361.4200 2046.9000 3364.4200 2047.3800 ;
        RECT 3361.4200 2052.3400 3364.4200 2052.8200 ;
        RECT 3361.4200 2057.7800 3364.4200 2058.2600 ;
        RECT 3361.4200 2063.2200 3364.4200 2063.7000 ;
        RECT 3361.4200 2068.6600 3364.4200 2069.1400 ;
        RECT 3361.4200 2074.1000 3364.4200 2074.5800 ;
        RECT 3305.7200 2084.9800 3307.3200 2085.4600 ;
        RECT 3305.7200 2079.5400 3307.3200 2080.0200 ;
        RECT 3305.7200 2090.4200 3307.3200 2090.9000 ;
        RECT 3305.7200 2095.8600 3307.3200 2096.3400 ;
        RECT 3305.7200 2101.3000 3307.3200 2101.7800 ;
        RECT 3305.7200 2106.7400 3307.3200 2107.2200 ;
        RECT 3305.7200 2112.1800 3307.3200 2112.6600 ;
        RECT 3305.7200 2117.6200 3307.3200 2118.1000 ;
        RECT 3305.7200 2123.0600 3307.3200 2123.5400 ;
        RECT 3361.4200 2079.5400 3364.4200 2080.0200 ;
        RECT 3361.4200 2084.9800 3364.4200 2085.4600 ;
        RECT 3361.4200 2090.4200 3364.4200 2090.9000 ;
        RECT 3361.4200 2095.8600 3364.4200 2096.3400 ;
        RECT 3361.4200 2101.3000 3364.4200 2101.7800 ;
        RECT 3361.4200 2106.7400 3364.4200 2107.2200 ;
        RECT 3361.4200 2112.1800 3364.4200 2112.6600 ;
        RECT 3361.4200 2117.6200 3364.4200 2118.1000 ;
        RECT 3361.4200 2123.0600 3364.4200 2123.5400 ;
        RECT 1733.7400 2228.5000 1735.3400 2228.9800 ;
        RECT 1733.8400 2489.2200 1735.4400 2489.7000 ;
        RECT 1740.9000 2458.1400 1742.5000 2458.6200 ;
        RECT 1716.1200 2520.1800 1717.7200 2520.6600 ;
        RECT 1726.3800 2520.1800 1727.9800 2520.6600 ;
        RECT 1733.8400 2520.1800 1735.4400 2520.6600 ;
        RECT 1716.1200 2525.6200 1717.7200 2526.1000 ;
        RECT 1716.1200 2531.0600 1717.7200 2531.5400 ;
        RECT 1733.8400 2525.6200 1735.4400 2526.1000 ;
        RECT 1726.3800 2525.6200 1727.9800 2526.1000 ;
        RECT 1726.3800 2531.0600 1727.9800 2531.5400 ;
        RECT 1733.8400 2531.0600 1735.4400 2531.5400 ;
        RECT 1716.1200 2536.5000 1717.7200 2536.9800 ;
        RECT 1716.1200 2541.9400 1717.7200 2542.4200 ;
        RECT 1716.1200 2547.3800 1717.7200 2547.8600 ;
        RECT 1726.3800 2541.9400 1727.9800 2542.4200 ;
        RECT 1733.8400 2541.9400 1735.4400 2542.4200 ;
        RECT 1726.3800 2536.5000 1727.9800 2536.9800 ;
        RECT 1733.8400 2536.5000 1735.4400 2536.9800 ;
        RECT 1726.3800 2547.3800 1727.9800 2547.8600 ;
        RECT 1733.8400 2547.3800 1735.4400 2547.8600 ;
        RECT 1941.3000 2464.4900 1942.9000 2466.0900 ;
        RECT 1953.9600 2456.9800 1955.5600 2457.4600 ;
        RECT 1954.0600 2489.2200 1955.6600 2489.7000 ;
        RECT 1936.3400 2520.1800 1937.9400 2520.6600 ;
        RECT 1946.6000 2520.1800 1948.2000 2520.6600 ;
        RECT 1946.6000 2525.6200 1948.2000 2526.1000 ;
        RECT 1936.3400 2525.6200 1937.9400 2526.1000 ;
        RECT 1936.3400 2531.0600 1937.9400 2531.5400 ;
        RECT 1946.6000 2531.0600 1948.2000 2531.5400 ;
        RECT 1936.3400 2541.9400 1937.9400 2542.4200 ;
        RECT 1946.6000 2541.9400 1948.2000 2542.4200 ;
        RECT 1936.3400 2536.5000 1937.9400 2536.9800 ;
        RECT 1946.6000 2536.5000 1948.2000 2536.9800 ;
        RECT 1936.3400 2547.3800 1937.9400 2547.8600 ;
        RECT 1946.6000 2547.3800 1948.2000 2547.8600 ;
        RECT 1954.0600 2520.1800 1955.6600 2520.6600 ;
        RECT 1954.0600 2525.6200 1955.6600 2526.1000 ;
        RECT 1954.0600 2531.0600 1955.6600 2531.5400 ;
        RECT 1954.0600 2536.5000 1955.6600 2536.9800 ;
        RECT 1954.0600 2541.9400 1955.6600 2542.4200 ;
        RECT 1954.0600 2547.3800 1955.6600 2547.8600 ;
        RECT 2174.1800 2228.5000 2175.7800 2228.9800 ;
        RECT 2394.4000 2228.5000 2396.0000 2228.9800 ;
        RECT 2447.1800 2128.5000 2448.7800 2128.9800 ;
        RECT 2447.1800 2133.9400 2448.7800 2134.4200 ;
        RECT 2447.1800 2139.3800 2448.7800 2139.8600 ;
        RECT 2447.1800 2144.8200 2448.7800 2145.3000 ;
        RECT 2447.1800 2150.2600 2448.7800 2150.7400 ;
        RECT 2447.1800 2166.5800 2448.7800 2167.0600 ;
        RECT 2447.1800 2155.7000 2448.7800 2156.1800 ;
        RECT 2447.1800 2161.1400 2448.7800 2161.6200 ;
        RECT 2447.1800 2172.0200 2448.7800 2172.5000 ;
        RECT 2447.1800 2177.4600 2448.7800 2177.9400 ;
        RECT 2492.9200 2128.5000 2494.5200 2128.9800 ;
        RECT 2492.9200 2133.9400 2494.5200 2134.4200 ;
        RECT 2492.9200 2139.3800 2494.5200 2139.8600 ;
        RECT 2492.9200 2144.8200 2494.5200 2145.3000 ;
        RECT 2492.9200 2150.2600 2494.5200 2150.7400 ;
        RECT 2492.9200 2166.5800 2494.5200 2167.0600 ;
        RECT 2492.9200 2161.1400 2494.5200 2161.6200 ;
        RECT 2492.9200 2155.7000 2494.5200 2156.1800 ;
        RECT 2492.9200 2172.0200 2494.5200 2172.5000 ;
        RECT 2492.9200 2177.4600 2494.5200 2177.9400 ;
        RECT 2447.1800 2182.9000 2448.7800 2183.3800 ;
        RECT 2447.1800 2188.3400 2448.7800 2188.8200 ;
        RECT 2447.1800 2193.7800 2448.7800 2194.2600 ;
        RECT 2447.1800 2199.2200 2448.7800 2199.7000 ;
        RECT 2447.1800 2204.6600 2448.7800 2205.1400 ;
        RECT 2447.1800 2210.1000 2448.7800 2210.5800 ;
        RECT 2447.1800 2215.5400 2448.7800 2216.0200 ;
        RECT 2447.1800 2220.9800 2448.7800 2221.4600 ;
        RECT 2447.1800 2226.4200 2448.7800 2226.9000 ;
        RECT 2447.1800 2231.8600 2448.7800 2232.3400 ;
        RECT 2492.9200 2182.9000 2494.5200 2183.3800 ;
        RECT 2492.9200 2188.3400 2494.5200 2188.8200 ;
        RECT 2492.9200 2193.7800 2494.5200 2194.2600 ;
        RECT 2492.9200 2199.2200 2494.5200 2199.7000 ;
        RECT 2492.9200 2204.6600 2494.5200 2205.1400 ;
        RECT 2492.9200 2210.1000 2494.5200 2210.5800 ;
        RECT 2492.9200 2215.5400 2494.5200 2216.0200 ;
        RECT 2492.9200 2220.9800 2494.5200 2221.4600 ;
        RECT 2492.9200 2226.4200 2494.5200 2226.9000 ;
        RECT 2492.9200 2231.8600 2494.5200 2232.3400 ;
        RECT 2394.4000 2262.3000 2396.0000 2262.7800 ;
        RECT 2447.1800 2259.0600 2448.7800 2259.5400 ;
        RECT 2447.1800 2237.3000 2448.7800 2237.7800 ;
        RECT 2447.1800 2242.7400 2448.7800 2244.3600 ;
        RECT 2447.1800 2248.1800 2448.7800 2248.6600 ;
        RECT 2447.1800 2264.5000 2448.7800 2264.9800 ;
        RECT 2447.1800 2269.9400 2448.7800 2270.4200 ;
        RECT 2447.1800 2275.3800 2448.7800 2275.8600 ;
        RECT 2447.1800 2280.8200 2448.7800 2281.3000 ;
        RECT 2492.9200 2259.0600 2494.5200 2259.5400 ;
        RECT 2492.9200 2242.7400 2494.5200 2243.2200 ;
        RECT 2492.9200 2237.3000 2494.5200 2237.7800 ;
        RECT 2492.9200 2248.1800 2494.5200 2248.6600 ;
        RECT 2492.9200 2253.6200 2494.5200 2254.1000 ;
        RECT 2492.9200 2269.9400 2494.5200 2270.4200 ;
        RECT 2492.9200 2264.5000 2494.5200 2264.9800 ;
        RECT 2492.9200 2275.3800 2494.5200 2275.8600 ;
        RECT 2492.9200 2280.8200 2494.5200 2281.3000 ;
        RECT 2447.1800 2286.2600 2448.7800 2286.7400 ;
        RECT 2447.1800 2291.7000 2448.7800 2292.1800 ;
        RECT 2447.1800 2297.1400 2448.7800 2297.6200 ;
        RECT 2447.1800 2302.5800 2448.7800 2303.0600 ;
        RECT 2447.1800 2308.0200 2448.7800 2308.5000 ;
        RECT 2447.1800 2313.4600 2448.7800 2313.9400 ;
        RECT 2447.1800 2318.9000 2448.7800 2319.3800 ;
        RECT 2447.1800 2324.3400 2448.7800 2324.8200 ;
        RECT 2447.1800 2329.7800 2448.7800 2330.2600 ;
        RECT 2447.1800 2335.2200 2448.7800 2335.7000 ;
        RECT 2492.9200 2286.2600 2494.5200 2286.7400 ;
        RECT 2492.9200 2291.7000 2494.5200 2292.1800 ;
        RECT 2492.9200 2297.1400 2494.5200 2297.6200 ;
        RECT 2492.9200 2302.5800 2494.5200 2303.0600 ;
        RECT 2492.9200 2308.0200 2494.5200 2308.5000 ;
        RECT 2492.9200 2318.9000 2494.5200 2319.3800 ;
        RECT 2492.9200 2313.4600 2494.5200 2313.9400 ;
        RECT 2492.9200 2324.3400 2494.5200 2324.8200 ;
        RECT 2492.9200 2329.7800 2494.5200 2330.2600 ;
        RECT 2492.9200 2335.2200 2494.5200 2335.7000 ;
        RECT 2166.8200 2464.4900 2168.4200 2467.1400 ;
        RECT 2181.3400 2458.1400 2182.9400 2458.6200 ;
        RECT 2174.2800 2489.2200 2175.8800 2489.7000 ;
        RECT 2156.5600 2520.1800 2158.1600 2520.6600 ;
        RECT 2156.5600 2525.6200 2158.1600 2526.1000 ;
        RECT 2156.5600 2531.0600 2158.1600 2531.5400 ;
        RECT 2156.5600 2536.5000 2158.1600 2536.9800 ;
        RECT 2156.5600 2541.9400 2158.1600 2542.4200 ;
        RECT 2156.5600 2547.3800 2158.1600 2547.8600 ;
        RECT 2166.8200 2520.1800 2168.4200 2520.6600 ;
        RECT 2174.2800 2520.1800 2175.8800 2520.6600 ;
        RECT 2166.8200 2525.6200 2168.4200 2526.1000 ;
        RECT 2166.8200 2531.0600 2168.4200 2531.5400 ;
        RECT 2174.2800 2525.6200 2175.8800 2526.1000 ;
        RECT 2174.2800 2531.0600 2175.8800 2531.5400 ;
        RECT 2166.8200 2536.5000 2168.4200 2536.9800 ;
        RECT 2166.8200 2541.9400 2168.4200 2542.4200 ;
        RECT 2166.8200 2547.3800 2168.4200 2547.8600 ;
        RECT 2174.2800 2536.5000 2175.8800 2536.9800 ;
        RECT 2174.2800 2541.9400 2175.8800 2542.4200 ;
        RECT 2174.2800 2547.3800 2175.8800 2547.8600 ;
        RECT 2447.1800 2340.6600 2448.7800 2341.1400 ;
        RECT 2447.1800 2346.1000 2448.7800 2346.5800 ;
        RECT 2447.1800 2351.5400 2448.7800 2352.0200 ;
        RECT 2447.1800 2356.9800 2448.7800 2357.4600 ;
        RECT 2447.1800 2362.4200 2448.7800 2362.9000 ;
        RECT 2447.1800 2367.8600 2448.7800 2368.3400 ;
        RECT 2447.1800 2373.3000 2448.7800 2373.7800 ;
        RECT 2447.1800 2378.7400 2448.7800 2379.2200 ;
        RECT 2447.1800 2384.1800 2448.7800 2384.6600 ;
        RECT 2447.1800 2389.6200 2448.7800 2390.1000 ;
        RECT 2492.9200 2346.1000 2494.5200 2346.5800 ;
        RECT 2492.9200 2340.6600 2494.5200 2341.1400 ;
        RECT 2492.9200 2351.5400 2494.5200 2352.0200 ;
        RECT 2492.9200 2356.9800 2494.5200 2357.4600 ;
        RECT 2492.9200 2362.4200 2494.5200 2362.9000 ;
        RECT 2492.9200 2367.8600 2494.5200 2368.3400 ;
        RECT 2492.9200 2373.3000 2494.5200 2373.7800 ;
        RECT 2492.9200 2378.7400 2494.5200 2379.2200 ;
        RECT 2492.9200 2384.1800 2494.5200 2384.6600 ;
        RECT 2492.9200 2389.6200 2494.5200 2390.1000 ;
        RECT 2447.1800 2416.8200 2448.7800 2417.3000 ;
        RECT 2447.1800 2395.0600 2448.7800 2395.5400 ;
        RECT 2447.1800 2400.5000 2448.7800 2400.9800 ;
        RECT 2447.1800 2405.9400 2448.7800 2406.4200 ;
        RECT 2447.1800 2411.3800 2448.7800 2411.8600 ;
        RECT 2447.1800 2422.2600 2448.7800 2422.7400 ;
        RECT 2447.1800 2427.7000 2448.7800 2428.1800 ;
        RECT 2447.1800 2433.1400 2448.7800 2433.6200 ;
        RECT 2447.1800 2438.5800 2448.7800 2439.0600 ;
        RECT 2492.9200 2416.8200 2494.5200 2417.3000 ;
        RECT 2492.9200 2400.5000 2494.5200 2400.9800 ;
        RECT 2492.9200 2395.0600 2494.5200 2395.5400 ;
        RECT 2492.9200 2405.9400 2494.5200 2406.4200 ;
        RECT 2492.9200 2411.3800 2494.5200 2411.8600 ;
        RECT 2492.9200 2427.7000 2494.5200 2428.1800 ;
        RECT 2492.9200 2422.2600 2494.5200 2422.7400 ;
        RECT 2492.9200 2433.1400 2494.5200 2433.6200 ;
        RECT 2492.9200 2438.5800 2494.5200 2439.0600 ;
        RECT 2387.0400 2482.1000 2388.6400 2482.5800 ;
        RECT 2387.0400 2487.5400 2388.6400 2488.0200 ;
        RECT 2387.0400 2492.9800 2388.6400 2493.4600 ;
        RECT 2387.0400 2498.4200 2388.6400 2498.9000 ;
        RECT 2387.0400 2503.8600 2388.6400 2504.3400 ;
        RECT 2376.7800 2520.1800 2378.3800 2520.6600 ;
        RECT 2387.0400 2514.7400 2388.6400 2515.2200 ;
        RECT 2387.0400 2509.3000 2388.6400 2509.7800 ;
        RECT 2387.0400 2520.1800 2388.6400 2520.6600 ;
        RECT 2376.7800 2525.6200 2378.3800 2526.1000 ;
        RECT 2376.7800 2531.0600 2378.3800 2531.5400 ;
        RECT 2387.0400 2525.6200 2388.6400 2526.1000 ;
        RECT 2387.0400 2531.0600 2388.6400 2531.5400 ;
        RECT 2376.7800 2536.5000 2378.3800 2536.9800 ;
        RECT 2376.7800 2541.9400 2378.3800 2542.4200 ;
        RECT 2376.7800 2547.3800 2378.3800 2547.8600 ;
        RECT 2387.0400 2536.5000 2388.6400 2536.9800 ;
        RECT 2387.0400 2541.9400 2388.6400 2542.4200 ;
        RECT 2387.0400 2547.3800 2388.6400 2547.8600 ;
        RECT 2447.1800 2444.0200 2448.7800 2444.5000 ;
        RECT 2447.1800 2449.4600 2448.7800 2449.9400 ;
        RECT 2447.1800 2454.9000 2448.7800 2455.3800 ;
        RECT 2447.1800 2460.3400 2448.7800 2460.8200 ;
        RECT 2447.1800 2464.4900 2448.7800 2466.2600 ;
        RECT 2447.1800 2471.2200 2448.7800 2471.7000 ;
        RECT 2447.1800 2482.1000 2448.7800 2482.5800 ;
        RECT 2437.0200 2482.1000 2438.6200 2482.5800 ;
        RECT 2447.1800 2476.6600 2448.7800 2477.1400 ;
        RECT 2447.1800 2487.5400 2448.7800 2488.0200 ;
        RECT 2437.0200 2487.5400 2438.6200 2488.0200 ;
        RECT 2447.1800 2492.9800 2448.7800 2493.4600 ;
        RECT 2437.0200 2492.9800 2438.6200 2493.4600 ;
        RECT 2492.9200 2444.0200 2494.5200 2444.5000 ;
        RECT 2492.9200 2449.4600 2494.5200 2449.9400 ;
        RECT 2492.9200 2454.9000 2494.5200 2455.3800 ;
        RECT 2492.9200 2460.3400 2494.5200 2460.8200 ;
        RECT 2492.9200 2465.7800 2494.5200 2466.2600 ;
        RECT 2492.9200 2476.6600 2494.5200 2477.1400 ;
        RECT 2492.9200 2471.2200 2494.5200 2471.7000 ;
        RECT 2492.9200 2482.1000 2494.5200 2482.5800 ;
        RECT 2492.9200 2487.5400 2494.5200 2488.0200 ;
        RECT 2492.9200 2492.9800 2494.5200 2493.4600 ;
        RECT 2447.1800 2498.4200 2448.7800 2498.9000 ;
        RECT 2437.0200 2498.4200 2438.6200 2498.9000 ;
        RECT 2447.1800 2503.8600 2448.7800 2504.3400 ;
        RECT 2437.0200 2503.8600 2438.6200 2504.3400 ;
        RECT 2437.0200 2514.7400 2438.6200 2515.2200 ;
        RECT 2437.0200 2509.3000 2438.6200 2509.7800 ;
        RECT 2447.1800 2509.3000 2448.7800 2509.7800 ;
        RECT 2447.1800 2514.7400 2448.7800 2515.2200 ;
        RECT 2437.0200 2520.1800 2438.6200 2520.6600 ;
        RECT 2447.1800 2520.1800 2448.7800 2520.6600 ;
        RECT 2447.1800 2525.6200 2448.7800 2526.1000 ;
        RECT 2437.0200 2525.6200 2438.6200 2526.1000 ;
        RECT 2437.0200 2531.0600 2438.6200 2531.5400 ;
        RECT 2447.1800 2531.0600 2448.7800 2531.5400 ;
        RECT 2437.0200 2541.9400 2438.6200 2542.4200 ;
        RECT 2447.1800 2541.9400 2448.7800 2542.4200 ;
        RECT 2437.0200 2536.5000 2438.6200 2536.9800 ;
        RECT 2447.1800 2536.5000 2448.7800 2536.9800 ;
        RECT 2437.0200 2547.3800 2438.6200 2547.8600 ;
        RECT 2447.1800 2547.3800 2448.7800 2547.8600 ;
        RECT 2492.9200 2503.8600 2494.5200 2504.3400 ;
        RECT 2492.9200 2498.4200 2494.5200 2498.9000 ;
        RECT 2492.9200 2509.3000 2494.5200 2509.7800 ;
        RECT 2492.9200 2514.7400 2494.5200 2515.2200 ;
        RECT 2492.9200 2520.1800 2494.5200 2520.6600 ;
        RECT 2492.9200 2525.6200 2494.5200 2526.1000 ;
        RECT 2492.9200 2531.0600 2494.5200 2531.5400 ;
        RECT 2492.9200 2536.5000 2494.5200 2536.9800 ;
        RECT 2492.9200 2541.9400 2494.5200 2542.4200 ;
        RECT 2492.9200 2547.3800 2494.5200 2547.8600 ;
        RECT 1716.1200 2552.8200 1717.7200 2553.3000 ;
        RECT 1716.1200 2558.2600 1717.7200 2558.7400 ;
        RECT 1733.8400 2552.8200 1735.4400 2553.3000 ;
        RECT 1726.3800 2552.8200 1727.9800 2553.3000 ;
        RECT 1733.8400 2558.2600 1735.4400 2558.7400 ;
        RECT 1726.3800 2558.2600 1727.9800 2558.7400 ;
        RECT 1946.6000 2552.8200 1948.2000 2553.3000 ;
        RECT 1936.3400 2552.8200 1937.9400 2553.3000 ;
        RECT 1946.6000 2558.2600 1948.2000 2558.7400 ;
        RECT 1936.3400 2558.2600 1937.9400 2558.7400 ;
        RECT 1954.0600 2552.8200 1955.6600 2553.3000 ;
        RECT 1954.0600 2558.2600 1955.6600 2558.7400 ;
        RECT 2156.5600 2552.8200 2158.1600 2553.3000 ;
        RECT 2156.5600 2558.2600 2158.1600 2558.7400 ;
        RECT 2166.8200 2552.8200 2168.4200 2553.3000 ;
        RECT 2166.8200 2558.2600 2168.4200 2558.7400 ;
        RECT 2174.2800 2552.8200 2175.8800 2553.3000 ;
        RECT 2174.2800 2558.2600 2175.8800 2558.7400 ;
        RECT 2376.7800 2558.2600 2378.3800 2558.7400 ;
        RECT 2376.7800 2552.8200 2378.3800 2553.3000 ;
        RECT 2387.0400 2552.8200 2388.6400 2553.3000 ;
        RECT 2387.0400 2558.2600 2388.6400 2558.7400 ;
        RECT 2447.1800 2552.8200 2448.7800 2553.3000 ;
        RECT 2437.0200 2552.8200 2438.6200 2553.3000 ;
        RECT 2447.1800 2558.2600 2448.7800 2558.7400 ;
        RECT 2437.0200 2558.2600 2438.6200 2558.7400 ;
        RECT 2492.9200 2552.8200 2494.5200 2553.3000 ;
        RECT 2492.9200 2558.2600 2494.5200 2558.7400 ;
        RECT 3305.7200 2128.5000 3307.3200 2128.9800 ;
        RECT 3305.7200 2133.9400 3307.3200 2134.4200 ;
        RECT 3305.7200 2139.3800 3307.3200 2139.8600 ;
        RECT 3305.7200 2144.8200 3307.3200 2145.3000 ;
        RECT 3305.7200 2150.2600 3307.3200 2150.7400 ;
        RECT 3305.7200 2166.5800 3307.3200 2167.0600 ;
        RECT 3305.7200 2161.1400 3307.3200 2161.6200 ;
        RECT 3305.7200 2155.7000 3307.3200 2156.1800 ;
        RECT 3305.7200 2172.0200 3307.3200 2172.5000 ;
        RECT 3305.7200 2177.4600 3307.3200 2177.9400 ;
        RECT 3361.4200 2128.5000 3364.4200 2128.9800 ;
        RECT 3361.4200 2133.9400 3364.4200 2134.4200 ;
        RECT 3361.4200 2139.3800 3364.4200 2139.8600 ;
        RECT 3361.4200 2144.8200 3364.4200 2145.3000 ;
        RECT 3361.4200 2150.2600 3364.4200 2150.7400 ;
        RECT 3361.4200 2166.5800 3364.4200 2167.0600 ;
        RECT 3361.4200 2155.7000 3364.4200 2156.1800 ;
        RECT 3361.4200 2161.1400 3364.4200 2161.6200 ;
        RECT 3361.4200 2172.0200 3364.4200 2172.5000 ;
        RECT 3361.4200 2177.4600 3364.4200 2177.9400 ;
        RECT 3305.7200 2182.9000 3307.3200 2183.3800 ;
        RECT 3305.7200 2188.3400 3307.3200 2188.8200 ;
        RECT 3305.7200 2193.7800 3307.3200 2194.2600 ;
        RECT 3305.7200 2199.2200 3307.3200 2199.7000 ;
        RECT 3305.7200 2204.6600 3307.3200 2205.1400 ;
        RECT 3305.7200 2210.1000 3307.3200 2210.5800 ;
        RECT 3305.7200 2215.5400 3307.3200 2216.0200 ;
        RECT 3305.7200 2220.9800 3307.3200 2221.4600 ;
        RECT 3305.7200 2226.4200 3307.3200 2226.9000 ;
        RECT 3305.7200 2231.8600 3307.3200 2232.3400 ;
        RECT 3361.4200 2182.9000 3364.4200 2183.3800 ;
        RECT 3361.4200 2188.3400 3364.4200 2188.8200 ;
        RECT 3361.4200 2193.7800 3364.4200 2194.2600 ;
        RECT 3361.4200 2199.2200 3364.4200 2199.7000 ;
        RECT 3361.4200 2204.6600 3364.4200 2205.1400 ;
        RECT 3361.4200 2210.1000 3364.4200 2210.5800 ;
        RECT 3361.4200 2215.5400 3364.4200 2216.0200 ;
        RECT 3361.4200 2220.9800 3364.4200 2221.4600 ;
        RECT 3361.4200 2226.4200 3364.4200 2226.9000 ;
        RECT 3361.4200 2231.8600 3364.4200 2232.3400 ;
        RECT 3305.7200 2259.0600 3307.3200 2259.5400 ;
        RECT 3305.7200 2242.7400 3307.3200 2243.2200 ;
        RECT 3305.7200 2237.3000 3307.3200 2237.7800 ;
        RECT 3305.7200 2248.1800 3307.3200 2248.6600 ;
        RECT 3305.7200 2253.6200 3307.3200 2254.1000 ;
        RECT 3305.7200 2269.9400 3307.3200 2270.4200 ;
        RECT 3305.7200 2264.5000 3307.3200 2264.9800 ;
        RECT 3305.7200 2275.3800 3307.3200 2275.8600 ;
        RECT 3305.7200 2280.8200 3307.3200 2281.3000 ;
        RECT 3361.4200 2259.0600 3364.4200 2259.5400 ;
        RECT 3361.4200 2237.3000 3364.4200 2237.7800 ;
        RECT 3361.4200 2242.7400 3364.4200 2243.2200 ;
        RECT 3361.4200 2248.1800 3364.4200 2248.6600 ;
        RECT 3361.4200 2253.6200 3364.4200 2254.1000 ;
        RECT 3361.4200 2264.5000 3364.4200 2264.9800 ;
        RECT 3361.4200 2269.9400 3364.4200 2270.4200 ;
        RECT 3361.4200 2275.3800 3364.4200 2275.8600 ;
        RECT 3361.4200 2280.8200 3364.4200 2281.3000 ;
        RECT 3305.7200 2286.2600 3307.3200 2286.7400 ;
        RECT 3305.7200 2291.7000 3307.3200 2292.1800 ;
        RECT 3305.7200 2297.1400 3307.3200 2297.6200 ;
        RECT 3305.7200 2302.5800 3307.3200 2303.0600 ;
        RECT 3305.7200 2308.0200 3307.3200 2308.5000 ;
        RECT 3305.7200 2318.9000 3307.3200 2319.3800 ;
        RECT 3305.7200 2313.4600 3307.3200 2313.9400 ;
        RECT 3305.7200 2324.3400 3307.3200 2324.8200 ;
        RECT 3305.7200 2329.7800 3307.3200 2330.2600 ;
        RECT 3305.7200 2335.2200 3307.3200 2335.7000 ;
        RECT 3361.4200 2286.2600 3364.4200 2286.7400 ;
        RECT 3361.4200 2291.7000 3364.4200 2292.1800 ;
        RECT 3361.4200 2297.1400 3364.4200 2297.6200 ;
        RECT 3361.4200 2302.5800 3364.4200 2303.0600 ;
        RECT 3361.4200 2308.0200 3364.4200 2308.5000 ;
        RECT 3361.4200 2313.4600 3364.4200 2313.9400 ;
        RECT 3361.4200 2318.9000 3364.4200 2319.3800 ;
        RECT 3361.4200 2324.3400 3364.4200 2324.8200 ;
        RECT 3361.4200 2329.7800 3364.4200 2330.2600 ;
        RECT 3361.4200 2335.2200 3364.4200 2335.7000 ;
        RECT 3305.7200 2346.1000 3307.3200 2346.5800 ;
        RECT 3305.7200 2340.6600 3307.3200 2341.1400 ;
        RECT 3305.7200 2351.5400 3307.3200 2352.0200 ;
        RECT 3305.7200 2356.9800 3307.3200 2357.4600 ;
        RECT 3305.7200 2362.4200 3307.3200 2362.9000 ;
        RECT 3305.7200 2367.8600 3307.3200 2368.3400 ;
        RECT 3305.7200 2373.3000 3307.3200 2373.7800 ;
        RECT 3305.7200 2378.7400 3307.3200 2379.2200 ;
        RECT 3305.7200 2384.1800 3307.3200 2384.6600 ;
        RECT 3305.7200 2389.6200 3307.3200 2390.1000 ;
        RECT 3361.4200 2340.6600 3364.4200 2341.1400 ;
        RECT 3361.4200 2346.1000 3364.4200 2346.5800 ;
        RECT 3361.4200 2351.5400 3364.4200 2352.0200 ;
        RECT 3361.4200 2356.9800 3364.4200 2357.4600 ;
        RECT 3361.4200 2362.4200 3364.4200 2362.9000 ;
        RECT 3361.4200 2367.8600 3364.4200 2368.3400 ;
        RECT 3361.4200 2373.3000 3364.4200 2373.7800 ;
        RECT 3361.4200 2378.7400 3364.4200 2379.2200 ;
        RECT 3361.4200 2384.1800 3364.4200 2384.6600 ;
        RECT 3361.4200 2389.6200 3364.4200 2390.1000 ;
        RECT 3305.7200 2416.8200 3307.3200 2417.3000 ;
        RECT 3305.7200 2400.5000 3307.3200 2400.9800 ;
        RECT 3305.7200 2395.0600 3307.3200 2395.5400 ;
        RECT 3305.7200 2405.9400 3307.3200 2406.4200 ;
        RECT 3305.7200 2411.3800 3307.3200 2411.8600 ;
        RECT 3305.7200 2427.7000 3307.3200 2428.1800 ;
        RECT 3305.7200 2422.2600 3307.3200 2422.7400 ;
        RECT 3305.7200 2433.1400 3307.3200 2433.6200 ;
        RECT 3305.7200 2438.5800 3307.3200 2439.0600 ;
        RECT 3361.4200 2416.8200 3364.4200 2417.3000 ;
        RECT 3361.4200 2395.0600 3364.4200 2395.5400 ;
        RECT 3361.4200 2400.5000 3364.4200 2400.9800 ;
        RECT 3361.4200 2405.9400 3364.4200 2406.4200 ;
        RECT 3361.4200 2411.3800 3364.4200 2411.8600 ;
        RECT 3361.4200 2422.2600 3364.4200 2422.7400 ;
        RECT 3361.4200 2427.7000 3364.4200 2428.1800 ;
        RECT 3361.4200 2433.1400 3364.4200 2433.6200 ;
        RECT 3361.4200 2438.5800 3364.4200 2439.0600 ;
        RECT 3305.7200 2444.0200 3307.3200 2444.5000 ;
        RECT 3305.7200 2449.4600 3307.3200 2449.9400 ;
        RECT 3305.7200 2454.9000 3307.3200 2455.3800 ;
        RECT 3305.7200 2460.3400 3307.3200 2460.8200 ;
        RECT 3305.7200 2465.7800 3307.3200 2466.2600 ;
        RECT 3305.7200 2476.6600 3307.3200 2477.1400 ;
        RECT 3305.7200 2471.2200 3307.3200 2471.7000 ;
        RECT 3305.7200 2482.1000 3307.3200 2482.5800 ;
        RECT 3305.7200 2487.5400 3307.3200 2488.0200 ;
        RECT 3305.7200 2492.9800 3307.3200 2493.4600 ;
        RECT 3361.4200 2444.0200 3364.4200 2444.5000 ;
        RECT 3361.4200 2449.4600 3364.4200 2449.9400 ;
        RECT 3361.4200 2454.9000 3364.4200 2455.3800 ;
        RECT 3361.4200 2460.3400 3364.4200 2460.8200 ;
        RECT 3361.4200 2465.7800 3364.4200 2466.2600 ;
        RECT 3361.4200 2471.2200 3364.4200 2471.7000 ;
        RECT 3361.4200 2476.6600 3364.4200 2477.1400 ;
        RECT 3361.4200 2482.1000 3364.4200 2482.5800 ;
        RECT 3361.4200 2487.5400 3364.4200 2488.0200 ;
        RECT 3361.4200 2492.9800 3364.4200 2493.4600 ;
        RECT 3305.7200 2503.8600 3307.3200 2504.3400 ;
        RECT 3305.7200 2498.4200 3307.3200 2498.9000 ;
        RECT 3305.7200 2509.3000 3307.3200 2509.7800 ;
        RECT 3305.7200 2514.7400 3307.3200 2515.2200 ;
        RECT 3305.7200 2520.1800 3307.3200 2520.6600 ;
        RECT 3305.7200 2525.6200 3307.3200 2526.1000 ;
        RECT 3305.7200 2531.0600 3307.3200 2531.5400 ;
        RECT 3305.7200 2536.5000 3307.3200 2536.9800 ;
        RECT 3305.7200 2541.9400 3307.3200 2542.4200 ;
        RECT 3305.7200 2547.3800 3307.3200 2547.8600 ;
        RECT 3361.4200 2498.4200 3364.4200 2498.9000 ;
        RECT 3361.4200 2503.8600 3364.4200 2504.3400 ;
        RECT 3361.4200 2509.3000 3364.4200 2509.7800 ;
        RECT 3361.4200 2514.7400 3364.4200 2515.2200 ;
        RECT 3361.4200 2520.1800 3364.4200 2520.6600 ;
        RECT 3361.4200 2525.6200 3364.4200 2526.1000 ;
        RECT 3361.4200 2531.0600 3364.4200 2531.5400 ;
        RECT 3361.4200 2536.5000 3364.4200 2536.9800 ;
        RECT 3361.4200 2541.9400 3364.4200 2542.4200 ;
        RECT 3361.4200 2547.3800 3364.4200 2547.8600 ;
        RECT 3305.7200 2552.8200 3307.3200 2553.3000 ;
        RECT 3305.7200 2558.2600 3307.3200 2558.7400 ;
        RECT 3361.4200 2558.2600 3364.4200 2558.7400 ;
        RECT 3361.4200 2552.8200 3364.4200 2553.3000 ;
      LAYER met4 ;
        RECT 1002.9200 176.2600 1004.5200 2563.7200 ;
        RECT 1065.8600 6.0000 1067.4600 2563.7200 ;
        RECT 1285.9400 6.0000 1287.5400 2563.7200 ;
        RECT 1286.0800 6.0000 1287.6800 2563.7200 ;
        RECT 1506.1600 6.0000 1507.7600 2563.7200 ;
        RECT 6.0000 6.0000 9.0000 2563.7200 ;
        RECT 965.7200 635.5400 967.3200 2014.9800 ;
        RECT 152.9200 635.5400 154.5200 2014.9800 ;
        RECT 1726.3800 6.0000 1727.9800 2563.7200 ;
        RECT 1946.6000 6.0000 1948.2000 2563.7200 ;
        RECT 2166.8200 6.0000 2168.4200 2563.7200 ;
        RECT 2387.0400 6.0000 2388.6400 2563.7200 ;
        RECT 2447.1800 6.0000 2448.7800 2563.7200 ;
        RECT 2492.9200 6.0000 2494.5200 2563.7200 ;
        RECT 3305.7200 6.0000 3307.3200 2563.7200 ;
        RECT 3361.4200 6.0000 3364.4200 2563.7200 ;
        RECT 502.9200 176.2600 504.5200 637.1400 ;
        RECT 665.7200 176.2600 667.3200 637.1400 ;
        RECT 1013.1800 176.2600 1014.7800 184.2600 ;
        RECT 1073.2200 177.7800 1074.8200 184.2600 ;
        RECT 1055.6000 176.2600 1057.2000 184.2600 ;
        RECT 1073.3200 136.0000 1074.9200 144.0000 ;
        RECT 1073.3200 163.9400 1074.9200 177.8600 ;
        RECT 1073.3200 172.6600 1074.9200 177.8600 ;
        RECT 1013.1800 402.3000 1014.7800 407.5000 ;
        RECT 1013.1800 391.8800 1014.7800 407.5000 ;
        RECT 1013.1800 405.9000 1014.7800 413.9000 ;
        RECT 1055.6000 402.3000 1057.2000 407.5000 ;
        RECT 1055.6000 405.9000 1057.2000 413.9000 ;
        RECT 1293.3000 177.3100 1294.9000 184.0000 ;
        RECT 1275.9200 177.7800 1277.5200 184.2600 ;
        RECT 1275.8200 136.0000 1277.4200 144.0000 ;
        RECT 1293.4000 135.7400 1295.0000 143.7400 ;
        RECT 1293.4000 163.6800 1295.0000 177.6000 ;
        RECT 1293.4000 172.4000 1295.0000 177.6000 ;
        RECT 1275.8200 172.6600 1277.4200 177.8600 ;
        RECT 1496.0000 177.3100 1497.6000 184.0000 ;
        RECT 1513.5200 177.3100 1515.1200 184.0000 ;
        RECT 1495.9000 135.7400 1497.5000 143.7400 ;
        RECT 1513.6200 135.7400 1515.2200 143.7400 ;
        RECT 1495.9000 172.4000 1497.5000 177.6000 ;
        RECT 1513.6200 163.6800 1515.2200 177.6000 ;
        RECT 1513.6200 172.4000 1515.2200 177.6000 ;
        RECT 1293.3000 391.6200 1294.9000 407.2400 ;
        RECT 1293.3000 402.0400 1294.9000 407.2400 ;
        RECT 1293.3000 405.6400 1294.9000 413.6400 ;
        RECT 1496.0000 405.6400 1497.6000 413.6400 ;
        RECT 1513.5200 402.0400 1515.1200 407.2400 ;
        RECT 1496.0000 402.0400 1497.6000 407.2400 ;
        RECT 1513.5200 391.6200 1515.1200 407.2400 ;
        RECT 1513.5200 405.6400 1515.1200 413.6400 ;
        RECT 1513.5200 850.9000 1515.1200 866.5200 ;
        RECT 1293.3000 850.9000 1294.9000 866.5200 ;
        RECT 1496.0000 861.3200 1497.6000 866.5200 ;
        RECT 1513.5200 861.3200 1515.1200 866.5200 ;
        RECT 1293.3000 861.3200 1294.9000 866.5200 ;
        RECT 1013.1800 851.1600 1014.7800 866.7800 ;
        RECT 1055.6000 861.5800 1057.2000 866.7800 ;
        RECT 1013.1800 861.5800 1014.7800 866.7800 ;
        RECT 1013.1800 635.5400 1014.7800 643.5400 ;
        RECT 1013.1800 631.9400 1014.7800 637.1400 ;
        RECT 1055.6000 621.5200 1057.2000 637.1400 ;
        RECT 1073.2200 620.3600 1074.8200 637.1400 ;
        RECT 1055.6000 635.5400 1057.2000 643.5400 ;
        RECT 1073.2200 635.5400 1074.8200 643.5400 ;
        RECT 1073.2200 632.4800 1074.8200 637.1400 ;
        RECT 1055.6000 631.9400 1057.2000 637.1400 ;
        RECT 1293.3000 621.2600 1294.9000 636.8800 ;
        RECT 1275.9200 635.5400 1277.5200 643.5400 ;
        RECT 1275.9200 632.4800 1277.5200 637.1400 ;
        RECT 1293.3000 631.6800 1294.9000 636.8800 ;
        RECT 1293.3000 635.2800 1294.9000 643.2800 ;
        RECT 1513.5200 621.2600 1515.1200 636.8800 ;
        RECT 1496.0000 635.2800 1497.6000 643.2800 ;
        RECT 1496.0000 631.6800 1497.6000 636.8800 ;
        RECT 1513.5200 635.2800 1515.1200 643.2800 ;
        RECT 1513.5200 631.6800 1515.1200 636.8800 ;
        RECT 1055.6000 865.1800 1057.2000 873.1800 ;
        RECT 1013.1800 865.1800 1014.7800 873.1800 ;
        RECT 1013.1800 1094.8200 1014.7800 1102.8200 ;
        RECT 1013.1800 1091.2200 1014.7800 1096.4200 ;
        RECT 1073.2200 1094.8200 1074.8200 1102.8200 ;
        RECT 1055.6000 1094.8200 1057.2000 1102.8200 ;
        RECT 1055.6000 1091.2200 1057.2000 1096.4200 ;
        RECT 1055.6000 1080.8000 1057.2000 1096.4200 ;
        RECT 1073.2200 1091.7600 1074.8200 1096.4200 ;
        RECT 1073.2200 1079.6400 1074.8200 1096.4200 ;
        RECT 1293.3000 864.9200 1294.9000 872.9200 ;
        RECT 1496.0000 864.9200 1497.6000 872.9200 ;
        RECT 1513.5200 864.9200 1515.1200 872.9200 ;
        RECT 1293.3000 1094.5600 1294.9000 1102.5600 ;
        RECT 1275.9200 1094.8200 1277.5200 1102.8200 ;
        RECT 1293.3000 1080.5400 1294.9000 1096.1600 ;
        RECT 1293.3000 1090.9600 1294.9000 1096.1600 ;
        RECT 1275.9200 1091.7600 1277.5200 1096.4200 ;
        RECT 1496.0000 1094.5600 1497.6000 1102.5600 ;
        RECT 1513.5200 1094.5600 1515.1200 1102.5600 ;
        RECT 1513.5200 1080.5400 1515.1200 1096.1600 ;
        RECT 1496.0000 1090.9600 1497.6000 1096.1600 ;
        RECT 1513.5200 1090.9600 1515.1200 1096.1600 ;
        RECT 1733.7400 177.3100 1735.3400 184.0000 ;
        RECT 1716.2200 177.3100 1717.8200 184.0000 ;
        RECT 1716.1200 135.7400 1717.7200 143.7400 ;
        RECT 1733.8400 135.7400 1735.4400 143.7400 ;
        RECT 1733.8400 163.6800 1735.4400 177.6000 ;
        RECT 1733.8400 172.4000 1735.4400 177.6000 ;
        RECT 1716.1200 172.4000 1717.7200 177.6000 ;
        RECT 1936.4400 177.3100 1938.0400 184.0000 ;
        RECT 1953.9600 177.3100 1955.5600 184.0000 ;
        RECT 1936.3400 135.7400 1937.9400 143.7400 ;
        RECT 1936.3400 172.4000 1937.9400 177.6000 ;
        RECT 1954.0600 172.4000 1955.6600 177.6000 ;
        RECT 1954.0600 163.6800 1955.6600 177.6000 ;
        RECT 1954.0600 135.7400 1955.6600 143.7400 ;
        RECT 1716.2200 405.6400 1717.8200 413.6400 ;
        RECT 1733.7400 405.6400 1735.3400 413.6400 ;
        RECT 1733.7400 391.6200 1735.3400 407.2400 ;
        RECT 1733.7400 402.0400 1735.3400 407.2400 ;
        RECT 1716.2200 402.0400 1717.8200 407.2400 ;
        RECT 1936.4400 402.0400 1938.0400 407.2400 ;
        RECT 1936.4400 405.6400 1938.0400 413.6400 ;
        RECT 2156.6600 177.3100 2158.2600 184.0000 ;
        RECT 2174.1800 177.3100 2175.7800 184.0000 ;
        RECT 2156.5600 135.7400 2158.1600 143.7400 ;
        RECT 2156.5600 172.4000 2158.1600 177.6000 ;
        RECT 2174.2800 135.7400 2175.8800 143.7400 ;
        RECT 2174.2800 172.4000 2175.8800 177.6000 ;
        RECT 2174.2800 163.6800 2175.8800 177.6000 ;
        RECT 2394.4000 176.0000 2396.0000 184.0000 ;
        RECT 2376.8800 177.3100 2378.4800 184.0000 ;
        RECT 2376.7800 135.7400 2378.3800 143.7400 ;
        RECT 2387.0400 137.4600 2389.7500 137.9400 ;
        RECT 2376.7800 172.4000 2378.3800 177.6000 ;
        RECT 2437.0200 176.0000 2438.6200 184.0000 ;
        RECT 2174.1800 391.6200 2175.7800 407.2400 ;
        RECT 2174.1800 402.0400 2175.7800 407.2400 ;
        RECT 2174.1800 405.6400 2175.7800 413.6400 ;
        RECT 2394.4000 402.0400 2396.0000 407.2400 ;
        RECT 2394.4000 391.6200 2396.0000 407.2400 ;
        RECT 2376.8800 402.0400 2378.4800 407.2400 ;
        RECT 2394.4000 405.6400 2396.0000 413.6400 ;
        RECT 2376.8800 405.6400 2378.4800 413.6400 ;
        RECT 2447.1800 414.9000 2449.8900 415.3800 ;
        RECT 2437.0200 402.0400 2438.6200 407.2400 ;
        RECT 2437.0200 405.6400 2438.6200 413.6400 ;
        RECT 1733.7400 850.9000 1735.3400 866.5200 ;
        RECT 1936.4400 861.3200 1938.0400 866.5200 ;
        RECT 1733.7400 861.3200 1735.3400 866.5200 ;
        RECT 1716.2200 861.3200 1717.8200 866.5200 ;
        RECT 2394.4000 861.3200 2396.0000 866.5200 ;
        RECT 2437.0200 861.3200 2438.6200 866.5200 ;
        RECT 2394.4000 850.9000 2396.0000 866.5200 ;
        RECT 2174.1800 850.9000 2175.7800 866.5200 ;
        RECT 2376.8800 861.3200 2378.4800 866.5200 ;
        RECT 2174.1800 861.3200 2175.7800 866.5200 ;
        RECT 1733.7400 635.2800 1735.3400 643.2800 ;
        RECT 1733.7400 621.2600 1735.3400 636.8800 ;
        RECT 1733.7400 631.6800 1735.3400 636.8800 ;
        RECT 1716.2200 635.2800 1717.8200 643.2800 ;
        RECT 1716.2200 631.6800 1717.8200 636.8800 ;
        RECT 1936.4400 635.2800 1938.0400 643.2800 ;
        RECT 1936.4400 631.6800 1938.0400 636.8800 ;
        RECT 1953.9600 620.1000 1955.5600 636.8800 ;
        RECT 1953.9600 635.2800 1955.5600 643.2800 ;
        RECT 1953.9600 632.2200 1955.5600 636.8800 ;
        RECT 2156.6600 635.2800 2158.2600 643.2800 ;
        RECT 2156.6600 632.2200 2158.2600 636.8800 ;
        RECT 2174.1800 621.2600 2175.7800 636.8800 ;
        RECT 2174.1800 631.6800 2175.7800 636.8800 ;
        RECT 2174.1800 635.2800 2175.7800 643.2800 ;
        RECT 2394.4000 631.6800 2396.0000 636.8800 ;
        RECT 2394.4000 621.2600 2396.0000 636.8800 ;
        RECT 2394.4000 635.2800 2396.0000 643.2800 ;
        RECT 2376.8800 635.2800 2378.4800 643.2800 ;
        RECT 2376.8800 631.6800 2378.4800 636.8800 ;
        RECT 2437.0200 635.2800 2438.6200 643.2800 ;
        RECT 2437.0200 631.6800 2438.6200 636.8800 ;
        RECT 1716.2200 864.9200 1717.8200 872.9200 ;
        RECT 1733.7400 864.9200 1735.3400 872.9200 ;
        RECT 1936.4400 864.9200 1938.0400 872.9200 ;
        RECT 1733.7400 1094.5600 1735.3400 1102.5600 ;
        RECT 1716.2200 1094.5600 1717.8200 1102.5600 ;
        RECT 1733.7400 1080.5400 1735.3400 1096.1600 ;
        RECT 1733.7400 1090.9600 1735.3400 1096.1600 ;
        RECT 1716.2200 1090.9600 1717.8200 1096.1600 ;
        RECT 1936.4400 1094.5600 1938.0400 1102.5600 ;
        RECT 1936.4400 1090.9600 1938.0400 1096.1600 ;
        RECT 1953.9600 1094.5600 1955.5600 1102.5600 ;
        RECT 1953.9600 1079.3800 1955.5600 1096.1600 ;
        RECT 1953.9600 1091.5000 1955.5600 1096.1600 ;
        RECT 2174.1800 864.9200 2175.7800 872.9200 ;
        RECT 2394.4000 864.9200 2396.0000 872.9200 ;
        RECT 2437.0200 864.9200 2438.6200 872.9200 ;
        RECT 2376.8800 864.9200 2378.4800 872.9200 ;
        RECT 2156.6600 1094.5600 2158.2600 1102.5600 ;
        RECT 2156.6600 1091.5000 2158.2600 1096.1600 ;
        RECT 2174.1800 1094.5600 2175.7800 1102.5600 ;
        RECT 2174.1800 1090.9600 2175.7800 1096.1600 ;
        RECT 2174.1800 1080.5400 2175.7800 1096.1600 ;
        RECT 2376.8800 1094.5600 2378.4800 1102.5600 ;
        RECT 2394.4000 1094.5600 2396.0000 1102.5600 ;
        RECT 2394.4000 1090.9600 2396.0000 1096.1600 ;
        RECT 2394.4000 1080.5400 2396.0000 1096.1600 ;
        RECT 2376.8800 1090.9600 2378.4800 1096.1600 ;
        RECT 2437.0200 1094.5600 2438.6200 1102.5600 ;
        RECT 2437.0200 1090.9600 2438.6200 1096.1600 ;
        RECT 1013.1800 1310.4400 1014.7800 1326.0600 ;
        RECT 1013.1800 1324.4600 1014.7800 1332.4600 ;
        RECT 1013.1800 1320.8600 1014.7800 1326.0600 ;
        RECT 1055.6000 1324.4600 1057.2000 1332.4600 ;
        RECT 1055.6000 1320.8600 1057.2000 1326.0600 ;
        RECT 1013.1800 1554.1000 1014.7800 1562.1000 ;
        RECT 1013.1800 1550.5000 1014.7800 1555.7000 ;
        RECT 1073.2200 1538.9200 1074.8200 1555.7000 ;
        RECT 1055.6000 1540.0800 1057.2000 1555.7000 ;
        RECT 1055.6000 1550.5000 1057.2000 1555.7000 ;
        RECT 1055.6000 1554.1000 1057.2000 1562.1000 ;
        RECT 1073.2200 1554.1000 1074.8200 1562.1000 ;
        RECT 1073.2200 1551.0400 1074.8200 1555.7000 ;
        RECT 1293.3000 1310.1800 1294.9000 1325.8000 ;
        RECT 1293.3000 1324.2000 1294.9000 1332.2000 ;
        RECT 1293.3000 1320.6000 1294.9000 1325.8000 ;
        RECT 1513.5200 1320.6000 1515.1200 1325.8000 ;
        RECT 1496.0000 1320.6000 1497.6000 1325.8000 ;
        RECT 1513.5200 1310.1800 1515.1200 1325.8000 ;
        RECT 1496.0000 1324.2000 1497.6000 1332.2000 ;
        RECT 1513.5200 1324.2000 1515.1200 1332.2000 ;
        RECT 1293.3000 1539.8200 1294.9000 1555.4400 ;
        RECT 1293.3000 1553.8400 1294.9000 1561.8400 ;
        RECT 1293.3000 1550.2400 1294.9000 1555.4400 ;
        RECT 1275.9200 1554.1000 1277.5200 1562.1000 ;
        RECT 1275.9200 1551.0400 1277.5200 1555.7000 ;
        RECT 1513.5200 1539.8200 1515.1200 1555.4400 ;
        RECT 1496.0000 1550.2400 1497.6000 1555.4400 ;
        RECT 1513.5200 1553.8400 1515.1200 1561.8400 ;
        RECT 1496.0000 1553.8400 1497.6000 1561.8400 ;
        RECT 1513.5200 1550.2400 1515.1200 1555.4400 ;
        RECT 1013.1800 1769.7200 1014.7800 1785.3400 ;
        RECT 1013.1800 1780.1400 1014.7800 1785.3400 ;
        RECT 1013.1800 1783.7400 1014.7800 1791.7400 ;
        RECT 1055.6000 1780.1400 1057.2000 1785.3400 ;
        RECT 1055.6000 1783.7400 1057.2000 1791.7400 ;
        RECT 1013.1800 2013.3800 1014.7800 2021.3800 ;
        RECT 1013.1800 2009.7800 1014.7800 2014.9800 ;
        RECT 1001.5800 2025.1400 1004.5200 2025.6200 ;
        RECT 1055.6000 1999.3600 1057.2000 2014.9800 ;
        RECT 1073.2200 1998.2000 1074.8200 2014.9800 ;
        RECT 1073.2200 2013.3800 1074.8200 2021.3800 ;
        RECT 1073.2200 2010.3200 1074.8200 2014.9800 ;
        RECT 1055.6000 2013.3800 1057.2000 2021.3800 ;
        RECT 1055.6000 2009.7800 1057.2000 2014.9800 ;
        RECT 1293.3000 1769.4600 1294.9000 1785.0800 ;
        RECT 1293.3000 1783.4800 1294.9000 1791.4800 ;
        RECT 1293.3000 1779.8800 1294.9000 1785.0800 ;
        RECT 1496.0000 1783.4800 1497.6000 1791.4800 ;
        RECT 1513.5200 1783.4800 1515.1200 1791.4800 ;
        RECT 1513.5200 1779.8800 1515.1200 1785.0800 ;
        RECT 1513.5200 1769.4600 1515.1200 1785.0800 ;
        RECT 1496.0000 1779.8800 1497.6000 1785.0800 ;
        RECT 1293.3000 2013.1200 1294.9000 2021.1200 ;
        RECT 1293.3000 1999.1000 1294.9000 2014.7200 ;
        RECT 1293.3000 2009.5200 1294.9000 2014.7200 ;
        RECT 1275.9200 2013.3800 1277.5200 2021.3800 ;
        RECT 1275.9200 2010.3200 1277.5200 2014.9800 ;
        RECT 1496.0000 2013.1200 1497.6000 2021.1200 ;
        RECT 1513.5200 1999.1000 1515.1200 2014.7200 ;
        RECT 1513.5200 2013.1200 1515.1200 2021.1200 ;
        RECT 1496.0000 2009.5200 1497.6000 2014.7200 ;
        RECT 1513.5200 2009.5200 1515.1200 2014.7200 ;
        RECT 1293.4000 2509.0600 1295.0000 2563.7200 ;
        RECT 1495.9000 2509.0600 1497.5000 2563.7200 ;
        RECT 1513.6200 2509.0600 1515.2200 2563.7200 ;
        RECT 1275.6800 2509.0600 1277.2800 2563.7200 ;
        RECT 1073.1800 2509.0600 1074.7800 2563.7200 ;
        RECT 1013.1800 2469.0600 1014.7800 2563.7200 ;
        RECT 1055.6000 2469.0600 1057.2000 2563.7200 ;
        RECT 1013.1800 2243.0200 1014.7800 2251.0200 ;
        RECT 1013.1800 2239.4200 1014.7800 2244.6200 ;
        RECT 1055.6000 2243.0200 1057.2000 2251.0200 ;
        RECT 1055.6000 2243.0200 1057.2000 2262.8000 ;
        RECT 1055.6000 2239.4200 1057.2000 2244.6200 ;
        RECT 1055.6000 2229.0000 1057.2000 2244.6200 ;
        RECT 1073.2200 2469.6000 1074.8200 2474.0000 ;
        RECT 1073.2200 2457.4800 1074.8200 2474.0000 ;
        RECT 1073.1800 2472.4000 1074.7800 2489.4600 ;
        RECT 1073.1800 2473.8200 1074.7800 2480.4000 ;
        RECT 1293.3000 2228.7400 1294.9000 2244.3600 ;
        RECT 1293.3000 2242.7600 1294.9000 2250.7600 ;
        RECT 1293.3000 2239.1600 1294.9000 2244.3600 ;
        RECT 1513.5200 2228.7400 1515.1200 2244.3600 ;
        RECT 1513.5200 2239.1600 1515.1200 2244.3600 ;
        RECT 1496.0000 2239.1600 1497.6000 2244.3600 ;
        RECT 1496.0000 2242.7600 1497.6000 2250.7600 ;
        RECT 1513.5200 2242.7600 1515.1200 2250.7600 ;
        RECT 1293.3000 2468.8000 1294.9000 2474.0000 ;
        RECT 1275.9200 2469.6000 1277.5200 2474.0000 ;
        RECT 1300.4600 2458.6200 1302.0600 2462.7250 ;
        RECT 1293.4000 2473.8200 1295.0000 2480.4000 ;
        RECT 1293.4000 2472.4000 1295.0000 2489.4600 ;
        RECT 1275.6800 2473.8200 1277.2800 2480.4000 ;
        RECT 1496.0000 2468.8000 1497.6000 2474.0000 ;
        RECT 1513.5200 2468.8000 1515.1200 2474.0000 ;
        RECT 1520.6800 2458.6200 1522.2800 2462.7250 ;
        RECT 1495.9000 2473.8200 1497.5000 2480.4000 ;
        RECT 1513.6200 2473.8200 1515.2200 2480.4000 ;
        RECT 1513.6200 2472.4000 1515.2200 2489.4600 ;
        RECT 1716.2200 1320.6000 1717.8200 1325.8000 ;
        RECT 1733.7400 1310.1800 1735.3400 1325.8000 ;
        RECT 1733.7400 1324.2000 1735.3400 1332.2000 ;
        RECT 1733.7400 1320.6000 1735.3400 1325.8000 ;
        RECT 1716.2200 1324.2000 1717.8200 1332.2000 ;
        RECT 1936.4400 1324.2000 1938.0400 1332.2000 ;
        RECT 1936.4400 1320.6000 1938.0400 1325.8000 ;
        RECT 1733.7400 1539.8200 1735.3400 1555.4400 ;
        RECT 1716.2200 1553.8400 1717.8200 1561.8400 ;
        RECT 1733.7400 1550.2400 1735.3400 1555.4400 ;
        RECT 1733.7400 1553.8400 1735.3400 1561.8400 ;
        RECT 1716.2200 1550.2400 1717.8200 1555.4400 ;
        RECT 1953.9600 1538.6600 1955.5600 1555.4400 ;
        RECT 1936.4400 1553.8400 1938.0400 1561.8400 ;
        RECT 1936.4400 1550.2400 1938.0400 1555.4400 ;
        RECT 1953.9600 1550.7800 1955.5600 1555.4400 ;
        RECT 1953.9600 1553.8400 1955.5600 1561.8400 ;
        RECT 2174.1800 1310.1800 2175.7800 1325.8000 ;
        RECT 2174.1800 1324.2000 2175.7800 1332.2000 ;
        RECT 2174.1800 1320.6000 2175.7800 1325.8000 ;
        RECT 2376.8800 1324.2000 2378.4800 1332.2000 ;
        RECT 2376.8800 1320.6000 2378.4800 1325.8000 ;
        RECT 2394.4000 1310.1800 2396.0000 1325.8000 ;
        RECT 2394.4000 1324.2000 2396.0000 1332.2000 ;
        RECT 2394.4000 1320.6000 2396.0000 1325.8000 ;
        RECT 2437.0200 1320.6000 2438.6200 1325.8000 ;
        RECT 2437.0200 1324.2000 2438.6200 1332.2000 ;
        RECT 2174.1800 1539.8200 2175.7800 1555.4400 ;
        RECT 2156.6600 1553.8400 2158.2600 1561.8400 ;
        RECT 2174.1800 1553.8400 2175.7800 1561.8400 ;
        RECT 2174.1800 1550.2400 2175.7800 1555.4400 ;
        RECT 2156.6600 1550.7800 2158.2600 1555.4400 ;
        RECT 2376.8800 1553.8400 2378.4800 1561.8400 ;
        RECT 2394.4000 1553.8400 2396.0000 1561.8400 ;
        RECT 2376.8800 1550.2400 2378.4800 1555.4400 ;
        RECT 2394.4000 1550.2400 2396.0000 1555.4400 ;
        RECT 2394.4000 1539.8200 2396.0000 1555.4400 ;
        RECT 2437.0200 1553.8400 2438.6200 1561.8400 ;
        RECT 2437.0200 1550.2400 2438.6200 1555.4400 ;
        RECT 1733.7400 1769.4600 1735.3400 1785.0800 ;
        RECT 1733.7400 1783.4800 1735.3400 1791.4800 ;
        RECT 1733.7400 1779.8800 1735.3400 1785.0800 ;
        RECT 1716.2200 1783.4800 1717.8200 1791.4800 ;
        RECT 1716.2200 1779.8800 1717.8200 1785.0800 ;
        RECT 1936.4400 1783.4800 1938.0400 1791.4800 ;
        RECT 1936.4400 1779.8800 1938.0400 1785.0800 ;
        RECT 1733.7400 2009.5200 1735.3400 2014.7200 ;
        RECT 1733.7400 2013.1200 1735.3400 2021.1200 ;
        RECT 1733.7400 1999.1000 1735.3400 2014.7200 ;
        RECT 1716.2200 2013.1200 1717.8200 2021.1200 ;
        RECT 1716.2200 2009.5200 1717.8200 2014.7200 ;
        RECT 1936.4400 2013.1200 1938.0400 2021.1200 ;
        RECT 1936.4400 2009.5200 1938.0400 2014.7200 ;
        RECT 1953.9600 2010.0600 1955.5600 2014.7200 ;
        RECT 1953.9600 2013.1200 1955.5600 2021.1200 ;
        RECT 1953.9600 1997.9400 1955.5600 2014.7200 ;
        RECT 2174.1800 1769.4600 2175.7800 1785.0800 ;
        RECT 2174.1800 1783.4800 2175.7800 1791.4800 ;
        RECT 2174.1800 1779.8800 2175.7800 1785.0800 ;
        RECT 2376.8800 1783.4800 2378.4800 1791.4800 ;
        RECT 2376.8800 1779.8800 2378.4800 1785.0800 ;
        RECT 2394.4000 1783.4800 2396.0000 1791.4800 ;
        RECT 2394.4000 1779.8800 2396.0000 1785.0800 ;
        RECT 2394.4000 1769.4600 2396.0000 1785.0800 ;
        RECT 2437.0200 1779.8800 2438.6200 1785.0800 ;
        RECT 2437.0200 1783.4800 2438.6200 1791.4800 ;
        RECT 2156.6600 2013.1200 2158.2600 2021.1200 ;
        RECT 2174.1800 1999.1000 2175.7800 2014.7200 ;
        RECT 2174.1800 2013.1200 2175.7800 2021.1200 ;
        RECT 2174.1800 2009.5200 2175.7800 2014.7200 ;
        RECT 2156.6600 2010.0600 2158.2600 2014.7200 ;
        RECT 2394.4000 1999.1000 2396.0000 2014.7200 ;
        RECT 2394.4000 2013.1200 2396.0000 2021.1200 ;
        RECT 2394.4000 2009.5200 2396.0000 2014.7200 ;
        RECT 2376.8800 2013.1200 2378.4800 2021.1200 ;
        RECT 2376.8800 2009.5200 2378.4800 2014.7200 ;
        RECT 2437.0200 2013.1200 2438.6200 2021.1200 ;
        RECT 2437.0200 2009.5200 2438.6200 2014.7200 ;
        RECT 1936.3400 2509.0600 1937.9400 2563.7200 ;
        RECT 1733.8400 2509.0600 1735.4400 2563.7200 ;
        RECT 1716.1200 2509.0600 1717.7200 2563.7200 ;
        RECT 2437.0200 2468.8000 2438.6200 2563.7200 ;
        RECT 1954.0600 2509.0600 1955.6600 2563.7200 ;
        RECT 2156.5600 2509.0600 2158.1600 2563.7200 ;
        RECT 2376.7800 2509.0600 2378.3800 2563.7200 ;
        RECT 2174.2800 2509.0600 2175.8800 2563.7200 ;
        RECT 1733.7400 2228.7400 1735.3400 2244.3600 ;
        RECT 1716.2200 2239.1600 1717.8200 2244.3600 ;
        RECT 1733.7400 2242.7600 1735.3400 2250.7600 ;
        RECT 1733.7400 2239.1600 1735.3400 2244.3600 ;
        RECT 1716.2200 2242.7600 1717.8200 2250.7600 ;
        RECT 1936.4400 2242.7600 1938.0400 2250.7600 ;
        RECT 1936.4400 2239.1600 1938.0400 2244.3600 ;
        RECT 1733.7400 2468.8000 1735.3400 2474.0000 ;
        RECT 1716.2200 2468.8000 1717.8200 2474.0000 ;
        RECT 1716.1200 2473.8200 1717.7200 2480.4000 ;
        RECT 1733.8400 2473.8200 1735.4400 2480.4000 ;
        RECT 1733.8400 2472.4000 1735.4400 2489.4600 ;
        RECT 1740.9000 2458.6200 1742.5000 2462.7250 ;
        RECT 1936.4400 2468.8000 1938.0400 2474.0000 ;
        RECT 1936.3400 2473.8200 1937.9400 2480.4000 ;
        RECT 1954.0600 2473.8200 1955.6600 2480.4000 ;
        RECT 1953.9600 2457.2200 1955.5600 2474.0000 ;
        RECT 1953.9600 2469.3400 1955.5600 2474.0000 ;
        RECT 1954.0600 2472.4000 1955.6600 2489.4600 ;
        RECT 2174.1800 2228.7400 2175.7800 2244.3600 ;
        RECT 2174.1800 2242.7600 2175.7800 2250.7600 ;
        RECT 2174.1800 2239.1600 2175.7800 2244.3600 ;
        RECT 2394.4000 2228.7400 2396.0000 2244.3600 ;
        RECT 2394.4000 2242.7600 2396.0000 2262.5400 ;
        RECT 2394.4000 2242.7600 2396.0000 2250.7600 ;
        RECT 2394.4000 2239.1600 2396.0000 2244.3600 ;
        RECT 2376.8800 2242.7600 2378.4800 2250.7600 ;
        RECT 2376.8800 2239.1600 2378.4800 2244.3600 ;
        RECT 2437.0200 2242.7600 2438.6200 2250.7600 ;
        RECT 2437.0200 2239.1600 2438.6200 2244.3600 ;
        RECT 2156.6600 2469.3400 2158.2600 2474.0000 ;
        RECT 2156.5600 2473.8200 2158.1600 2480.4000 ;
        RECT 2174.1800 2468.8000 2175.7800 2474.0000 ;
        RECT 2181.3400 2458.6200 2182.9400 2462.7250 ;
        RECT 2174.2800 2473.8200 2175.8800 2480.4000 ;
        RECT 2174.2800 2472.4000 2175.8800 2489.4600 ;
        RECT 2394.4000 2467.6600 2396.0000 2470.1600 ;
        RECT 2376.8800 2468.8000 2378.4800 2474.0000 ;
        RECT 2394.4000 2468.8000 2396.0000 2468.9100 ;
        RECT 2376.7800 2473.8200 2378.3800 2480.4000 ;
        RECT 1285.9400 6.0000 1287.6800 9.0000 ;
        RECT 1285.9400 12.3400 1287.6800 12.8200 ;
        RECT 1285.9400 17.7800 1287.6800 18.2600 ;
        RECT 1073.3200 163.7000 1074.9200 164.1800 ;
        RECT 1013.1800 391.6400 1014.7800 392.1200 ;
        RECT 1285.9400 34.1000 1287.6800 34.5800 ;
        RECT 1285.9400 28.6600 1287.6800 29.1400 ;
        RECT 1285.9400 23.2200 1287.6800 23.7000 ;
        RECT 1285.9400 39.5400 1287.6800 40.0200 ;
        RECT 1285.9400 44.9800 1287.6800 45.4600 ;
        RECT 1285.9400 50.4200 1287.6800 50.9000 ;
        RECT 1285.9400 55.8600 1287.6800 56.3400 ;
        RECT 1285.9400 61.3000 1287.6800 61.7800 ;
        RECT 1285.9400 66.7400 1287.6800 67.2200 ;
        RECT 1285.9400 72.1800 1287.6800 72.6600 ;
        RECT 1285.9400 77.6200 1287.6800 78.1000 ;
        RECT 1285.9400 83.0600 1287.6800 83.5400 ;
        RECT 1285.9400 88.5000 1287.6800 88.9800 ;
        RECT 1285.9400 93.9400 1287.6800 94.4200 ;
        RECT 1285.9400 99.3800 1287.6800 99.8600 ;
        RECT 1285.9400 110.2600 1287.6800 110.7400 ;
        RECT 1285.9400 104.8200 1287.6800 105.3000 ;
        RECT 1285.9400 115.7000 1287.6800 116.1800 ;
        RECT 1285.9400 121.1400 1287.6800 121.6200 ;
        RECT 1285.9400 126.5800 1287.6800 127.0600 ;
        RECT 1285.9400 144.5100 1287.6800 146.1100 ;
        RECT 1285.9400 135.7400 1287.6800 137.6000 ;
        RECT 1285.9400 132.0200 1287.6800 132.5000 ;
        RECT 1285.9400 176.0000 1287.6800 177.8600 ;
        RECT 1285.9400 168.8400 1287.6800 170.7000 ;
        RECT 1293.4000 163.4400 1295.0000 163.9200 ;
        RECT 1285.9400 186.0300 1287.6800 187.8900 ;
        RECT 1513.6200 163.4400 1515.2200 163.9200 ;
        RECT 1285.9400 405.6400 1287.6800 407.2400 ;
        RECT 1285.9400 397.7300 1287.6800 399.3300 ;
        RECT 1285.9400 415.6700 1287.6800 417.2700 ;
        RECT 1293.3000 391.3800 1294.9000 391.8600 ;
        RECT 1513.5200 391.3800 1515.1200 391.8600 ;
        RECT 1055.6000 621.2800 1057.2000 621.7600 ;
        RECT 1073.2200 620.1200 1074.8200 620.6000 ;
        RECT 1013.1800 850.9200 1014.7800 851.4000 ;
        RECT 1293.3000 621.0200 1294.9000 621.5000 ;
        RECT 1285.9400 635.2800 1287.6800 637.1400 ;
        RECT 1285.9400 627.3700 1287.6800 630.2800 ;
        RECT 1285.9400 645.3100 1287.6800 647.1700 ;
        RECT 1513.5200 621.0200 1515.1200 621.5000 ;
        RECT 1285.9400 857.0100 1287.6800 858.6100 ;
        RECT 1293.3000 850.6600 1294.9000 851.1400 ;
        RECT 1513.5200 850.6600 1515.1200 851.1400 ;
        RECT 1073.2200 1079.4000 1074.8200 1079.8800 ;
        RECT 1055.6000 1080.5600 1057.2000 1081.0400 ;
        RECT 1285.9400 864.9200 1287.6800 866.5200 ;
        RECT 1285.9400 874.9500 1287.6800 876.5500 ;
        RECT 1285.9400 1094.5600 1287.6800 1096.4200 ;
        RECT 1285.9400 1086.6500 1287.6800 1089.5600 ;
        RECT 1293.3000 1080.3000 1294.9000 1080.7800 ;
        RECT 1285.9400 1104.5900 1287.6800 1106.4500 ;
        RECT 1513.5200 1080.3000 1515.1200 1080.7800 ;
        RECT 1733.8400 163.4400 1735.4400 163.9200 ;
        RECT 1954.0600 163.4400 1955.6600 163.9200 ;
        RECT 1733.7400 391.3800 1735.3400 391.8600 ;
        RECT 2174.2800 163.4400 2175.8800 163.9200 ;
        RECT 2389.5000 137.4600 2390.0000 137.9400 ;
        RECT 2174.1800 391.3800 2175.7800 391.8600 ;
        RECT 2394.4000 391.3800 2396.0000 391.8600 ;
        RECT 2449.6400 414.9000 2450.1400 415.3800 ;
        RECT 1733.7400 621.0200 1735.3400 621.5000 ;
        RECT 1953.9600 619.8600 1955.5600 620.3400 ;
        RECT 1733.7400 850.6600 1735.3400 851.1400 ;
        RECT 2174.1800 621.0200 2175.7800 621.5000 ;
        RECT 2394.4000 621.0200 2396.0000 621.5000 ;
        RECT 2174.1800 850.6600 2175.7800 851.1400 ;
        RECT 2394.4000 850.6600 2396.0000 851.1400 ;
        RECT 1733.7400 1080.3000 1735.3400 1080.7800 ;
        RECT 1953.9600 1079.1400 1955.5600 1079.6200 ;
        RECT 2174.1800 1080.3000 2175.7800 1080.7800 ;
        RECT 2394.4000 1080.3000 2396.0000 1080.7800 ;
        RECT 1013.1800 1310.2000 1014.7800 1310.6800 ;
        RECT 1055.6000 1539.8400 1057.2000 1540.3200 ;
        RECT 1073.2200 1538.6800 1074.8200 1539.1600 ;
        RECT 1285.9400 1324.2000 1287.6800 1325.8000 ;
        RECT 1285.9400 1334.2300 1287.6800 1335.8300 ;
        RECT 1285.9400 1316.2900 1287.6800 1317.8900 ;
        RECT 1293.3000 1309.9400 1294.9000 1310.4200 ;
        RECT 1513.5200 1309.9400 1515.1200 1310.4200 ;
        RECT 1285.9400 1545.9300 1287.6800 1548.8400 ;
        RECT 1293.3000 1539.5800 1294.9000 1540.0600 ;
        RECT 1285.9400 1553.8400 1287.6800 1555.7000 ;
        RECT 1285.9400 1563.8700 1287.6800 1565.7300 ;
        RECT 1513.5200 1539.5800 1515.1200 1540.0600 ;
        RECT 1013.1800 1769.4800 1014.7800 1769.9600 ;
        RECT 1001.3300 2025.1400 1001.8300 2025.6200 ;
        RECT 1073.2200 1997.9600 1074.8200 1998.4400 ;
        RECT 1055.6000 1999.1200 1057.2000 1999.6000 ;
        RECT 1285.9400 1783.4800 1287.6800 1785.0800 ;
        RECT 1285.9400 1793.5100 1287.6800 1795.1100 ;
        RECT 1285.9400 1775.5700 1287.6800 1777.1700 ;
        RECT 1293.3000 1769.2200 1294.9000 1769.7000 ;
        RECT 1513.5200 1769.2200 1515.1200 1769.7000 ;
        RECT 1285.9400 2013.1200 1287.6800 2014.9800 ;
        RECT 1285.9400 2005.2100 1287.6800 2008.1200 ;
        RECT 1293.3000 1998.8600 1294.9000 1999.3400 ;
        RECT 1285.9400 2023.1500 1287.6800 2025.0100 ;
        RECT 1513.5200 1998.8600 1515.1200 1999.3400 ;
        RECT 1055.6000 2228.7600 1057.2000 2229.2400 ;
        RECT 1055.6000 2262.5600 1057.2000 2263.0400 ;
        RECT 1073.2200 2457.2400 1074.8200 2457.7200 ;
        RECT 1073.1800 2472.4000 1074.8200 2474.0000 ;
        RECT 1073.1800 2489.2200 1074.7800 2489.7000 ;
        RECT 1285.9400 2242.7600 1287.6800 2244.3600 ;
        RECT 1285.9400 2252.7900 1287.6800 2254.3900 ;
        RECT 1285.9400 2234.8500 1287.6800 2236.4500 ;
        RECT 1293.3000 2228.5000 1294.9000 2228.9800 ;
        RECT 1513.5200 2228.5000 1515.1200 2228.9800 ;
        RECT 1285.9400 2464.4900 1287.6800 2467.4000 ;
        RECT 1300.4600 2458.1400 1302.0600 2458.6200 ;
        RECT 1285.9400 2472.4000 1287.6800 2474.0000 ;
        RECT 1285.9400 2481.1700 1287.6800 2482.7700 ;
        RECT 1293.3000 2472.4000 1295.0000 2474.0000 ;
        RECT 1293.4000 2489.2200 1295.0000 2489.7000 ;
        RECT 1285.9400 2505.5000 1287.6800 2507.1000 ;
        RECT 1285.9400 2520.1800 1287.6800 2520.6600 ;
        RECT 1285.9400 2525.6200 1287.6800 2526.1000 ;
        RECT 1285.9400 2531.0600 1287.6800 2531.5400 ;
        RECT 1285.9400 2536.5000 1287.6800 2536.9800 ;
        RECT 1285.9400 2541.9400 1287.6800 2542.4200 ;
        RECT 1285.9400 2547.3800 1287.6800 2547.8600 ;
        RECT 1520.6800 2458.1400 1522.2800 2458.6200 ;
        RECT 1513.5200 2472.4000 1515.2200 2474.0000 ;
        RECT 1513.6200 2489.2200 1515.2200 2489.7000 ;
        RECT 1285.9400 2560.7200 1287.6800 2563.7200 ;
        RECT 1285.9400 2552.8200 1287.6800 2553.3000 ;
        RECT 1285.9400 2558.2600 1287.6800 2558.7400 ;
        RECT 1733.7400 1309.9400 1735.3400 1310.4200 ;
        RECT 1733.7400 1539.5800 1735.3400 1540.0600 ;
        RECT 1953.9600 1538.4200 1955.5600 1538.9000 ;
        RECT 2174.1800 1309.9400 2175.7800 1310.4200 ;
        RECT 2394.4000 1309.9400 2396.0000 1310.4200 ;
        RECT 2174.1800 1539.5800 2175.7800 1540.0600 ;
        RECT 2394.4000 1539.5800 2396.0000 1540.0600 ;
        RECT 1733.7400 1769.2200 1735.3400 1769.7000 ;
        RECT 1733.7400 1998.8600 1735.3400 1999.3400 ;
        RECT 1953.9600 1997.7000 1955.5600 1998.1800 ;
        RECT 2174.1800 1769.2200 2175.7800 1769.7000 ;
        RECT 2394.4000 1769.2200 2396.0000 1769.7000 ;
        RECT 2174.1800 1998.8600 2175.7800 1999.3400 ;
        RECT 2394.4000 1998.8600 2396.0000 1999.3400 ;
        RECT 1733.7400 2228.5000 1735.3400 2228.9800 ;
        RECT 1733.7400 2472.4000 1735.4400 2474.0000 ;
        RECT 1733.8400 2489.2200 1735.4400 2489.7000 ;
        RECT 1740.9000 2458.1400 1742.5000 2458.6200 ;
        RECT 1953.9600 2456.9800 1955.5600 2457.4600 ;
        RECT 1953.9600 2472.4000 1955.6600 2474.0000 ;
        RECT 1954.0600 2489.2200 1955.6600 2489.7000 ;
        RECT 2174.1800 2228.5000 2175.7800 2228.9800 ;
        RECT 2394.4000 2228.5000 2396.0000 2228.9800 ;
        RECT 2394.4000 2262.3000 2396.0000 2262.7800 ;
        RECT 2181.3400 2458.1400 2182.9400 2458.6200 ;
        RECT 2174.1800 2472.4000 2175.8800 2474.0000 ;
        RECT 2174.2800 2489.2200 2175.8800 2489.7000 ;
        RECT 647.8800 457.2200 649.4800 458.8200 ;
        RECT 1060.5600 627.5300 1062.1600 629.1300 ;
        RECT 1060.5600 1086.8100 1062.1600 1088.4100 ;
        RECT 1941.3000 627.3700 1942.9000 628.9700 ;
        RECT 1941.3000 1086.6500 1942.9000 1088.2500 ;
        RECT 1060.5600 1546.0900 1062.1600 1547.6900 ;
        RECT 947.8800 1905.9000 949.4800 1907.5000 ;
        RECT 1060.5600 2005.3700 1062.1600 2006.9700 ;
        RECT 1060.5600 2464.6500 1062.1600 2466.2500 ;
        RECT 1300.4600 2461.9250 1302.0600 2463.5250 ;
        RECT 1300.4600 2472.4000 1302.0600 2474.0000 ;
        RECT 1520.6800 2461.9250 1522.2800 2463.5250 ;
        RECT 1520.6800 2472.4000 1522.2800 2474.0000 ;
        RECT 1941.3000 1545.9300 1942.9000 1547.5300 ;
        RECT 1941.3000 2005.2100 1942.9000 2006.8100 ;
        RECT 3287.8800 1905.9000 3289.4800 1907.5000 ;
        RECT 1740.9000 2461.9250 1742.5000 2463.5250 ;
        RECT 1740.9000 2472.4000 1742.5000 2474.0000 ;
        RECT 1941.3000 2464.4900 1942.9000 2466.0900 ;
        RECT 2181.3400 2461.9250 2182.9400 2463.5250 ;
        RECT 2181.3400 2472.4000 2182.9400 2474.0000 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'core_sram'
    PORT
      LAYER met4 ;
        RECT 171.0800 1905.9000 949.4800 1907.5000 ;
    END
# end of P/G pin shape extracted from block 'core_sram'


# P/G pin shape extracted from block 'core_sram'
    PORT
      LAYER met4 ;
        RECT 2511.0800 1905.9000 3289.4800 1907.5000 ;
    END
# end of P/G pin shape extracted from block 'core_sram'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 183.4600 1057.2000 403.1000 ;
        RECT 1013.1800 183.4600 1014.7800 403.1000 ;
      LAYER met3 ;
        RECT 1055.6000 391.6400 1057.2000 392.1200 ;
        RECT 1055.6000 380.7600 1057.2000 381.2400 ;
        RECT 1055.6000 386.2000 1057.2000 386.6800 ;
        RECT 1055.6000 364.4400 1057.2000 364.9200 ;
        RECT 1055.6000 369.8800 1057.2000 370.3600 ;
        RECT 1055.6000 353.5600 1057.2000 354.0400 ;
        RECT 1055.6000 359.0000 1057.2000 359.4800 ;
        RECT 1055.6000 375.3200 1057.2000 375.8000 ;
        RECT 1055.6000 337.2400 1057.2000 337.7200 ;
        RECT 1055.6000 342.6800 1057.2000 343.1600 ;
        RECT 1055.6000 320.9200 1057.2000 321.4000 ;
        RECT 1055.6000 326.3600 1057.2000 326.8400 ;
        RECT 1055.6000 331.8000 1057.2000 332.2800 ;
        RECT 1055.6000 310.0400 1057.2000 310.5200 ;
        RECT 1055.6000 315.4800 1057.2000 315.9600 ;
        RECT 1055.6000 293.7200 1057.2000 294.2000 ;
        RECT 1055.6000 299.1600 1057.2000 299.6400 ;
        RECT 1055.6000 304.6000 1057.2000 305.0800 ;
        RECT 1055.6000 348.1200 1057.2000 348.6000 ;
        RECT 1013.1800 391.6400 1014.7800 392.1200 ;
        RECT 1013.1800 380.7600 1014.7800 381.2400 ;
        RECT 1013.1800 386.2000 1014.7800 386.6800 ;
        RECT 1013.1800 364.4400 1014.7800 364.9200 ;
        RECT 1013.1800 369.8800 1014.7800 370.3600 ;
        RECT 1013.1800 353.5600 1014.7800 354.0400 ;
        RECT 1013.1800 359.0000 1014.7800 359.4800 ;
        RECT 1013.1800 375.3200 1014.7800 375.8000 ;
        RECT 1013.1800 337.2400 1014.7800 337.7200 ;
        RECT 1013.1800 342.6800 1014.7800 343.1600 ;
        RECT 1013.1800 320.9200 1014.7800 321.4000 ;
        RECT 1013.1800 326.3600 1014.7800 326.8400 ;
        RECT 1013.1800 331.8000 1014.7800 332.2800 ;
        RECT 1013.1800 310.0400 1014.7800 310.5200 ;
        RECT 1013.1800 315.4800 1014.7800 315.9600 ;
        RECT 1013.1800 293.7200 1014.7800 294.2000 ;
        RECT 1013.1800 299.1600 1014.7800 299.6400 ;
        RECT 1013.1800 304.6000 1014.7800 305.0800 ;
        RECT 1013.1800 348.1200 1014.7800 348.6000 ;
        RECT 1055.6000 282.8400 1057.2000 283.3200 ;
        RECT 1055.6000 288.2800 1057.2000 288.7600 ;
        RECT 1055.6000 266.5200 1057.2000 267.0000 ;
        RECT 1055.6000 271.9600 1057.2000 272.4400 ;
        RECT 1055.6000 277.4000 1057.2000 277.8800 ;
        RECT 1055.6000 255.6400 1057.2000 256.1200 ;
        RECT 1055.6000 261.0800 1057.2000 261.5600 ;
        RECT 1055.6000 239.3200 1057.2000 239.8000 ;
        RECT 1055.6000 244.7600 1057.2000 245.2400 ;
        RECT 1055.6000 250.2000 1057.2000 250.6800 ;
        RECT 1055.6000 228.4400 1057.2000 228.9200 ;
        RECT 1055.6000 233.8800 1057.2000 234.3600 ;
        RECT 1055.6000 212.1200 1057.2000 212.6000 ;
        RECT 1055.6000 217.5600 1057.2000 218.0400 ;
        RECT 1055.6000 223.0000 1057.2000 223.4800 ;
        RECT 1055.6000 201.2400 1057.2000 201.7200 ;
        RECT 1055.6000 206.6800 1057.2000 207.1600 ;
        RECT 1055.6000 195.8000 1057.2000 196.2800 ;
        RECT 1013.1800 282.8400 1014.7800 283.3200 ;
        RECT 1013.1800 288.2800 1014.7800 288.7600 ;
        RECT 1013.1800 266.5200 1014.7800 267.0000 ;
        RECT 1013.1800 271.9600 1014.7800 272.4400 ;
        RECT 1013.1800 277.4000 1014.7800 277.8800 ;
        RECT 1013.1800 255.6400 1014.7800 256.1200 ;
        RECT 1013.1800 261.0800 1014.7800 261.5600 ;
        RECT 1013.1800 239.3200 1014.7800 239.8000 ;
        RECT 1013.1800 244.7600 1014.7800 245.2400 ;
        RECT 1013.1800 250.2000 1014.7800 250.6800 ;
        RECT 1013.1800 228.4400 1014.7800 228.9200 ;
        RECT 1013.1800 233.8800 1014.7800 234.3600 ;
        RECT 1013.1800 212.1200 1014.7800 212.6000 ;
        RECT 1013.1800 217.5600 1014.7800 218.0400 ;
        RECT 1013.1800 223.0000 1014.7800 223.4800 ;
        RECT 1013.1800 201.2400 1014.7800 201.7200 ;
        RECT 1013.1800 206.6800 1014.7800 207.1600 ;
        RECT 1013.1800 195.8000 1014.7800 196.2800 ;
        RECT 1010.1200 397.8900 1060.2600 399.4900 ;
        RECT 1010.1200 186.3900 1060.2600 187.9900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 183.4600 1014.7800 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 401.5000 1014.7800 403.1000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 183.4600 1057.2000 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 401.5000 1057.2000 403.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 186.3900 1011.7200 187.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 186.3900 1060.2600 187.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 397.8900 1011.7200 399.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 397.8900 1060.2600 399.4900 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 2250.2200 1057.2000 2469.8600 ;
        RECT 1013.1800 2250.2200 1014.7800 2469.8600 ;
      LAYER met3 ;
        RECT 1055.6000 2458.4000 1057.2000 2458.8800 ;
        RECT 1055.6000 2447.5200 1057.2000 2448.0000 ;
        RECT 1055.6000 2452.9600 1057.2000 2453.4400 ;
        RECT 1055.6000 2431.2000 1057.2000 2431.6800 ;
        RECT 1055.6000 2436.6400 1057.2000 2437.1200 ;
        RECT 1055.6000 2420.3200 1057.2000 2420.8000 ;
        RECT 1055.6000 2425.7600 1057.2000 2426.2400 ;
        RECT 1055.6000 2442.0800 1057.2000 2442.5600 ;
        RECT 1055.6000 2404.0000 1057.2000 2404.4800 ;
        RECT 1055.6000 2409.4400 1057.2000 2409.9200 ;
        RECT 1055.6000 2387.6800 1057.2000 2388.1600 ;
        RECT 1055.6000 2393.1200 1057.2000 2393.6000 ;
        RECT 1055.6000 2398.5600 1057.2000 2399.0400 ;
        RECT 1055.6000 2376.8000 1057.2000 2377.2800 ;
        RECT 1055.6000 2382.2400 1057.2000 2382.7200 ;
        RECT 1055.6000 2360.4800 1057.2000 2360.9600 ;
        RECT 1055.6000 2365.9200 1057.2000 2366.4000 ;
        RECT 1055.6000 2371.3600 1057.2000 2371.8400 ;
        RECT 1055.6000 2414.8800 1057.2000 2415.3600 ;
        RECT 1013.1800 2458.4000 1014.7800 2458.8800 ;
        RECT 1013.1800 2447.5200 1014.7800 2448.0000 ;
        RECT 1013.1800 2452.9600 1014.7800 2453.4400 ;
        RECT 1013.1800 2431.2000 1014.7800 2431.6800 ;
        RECT 1013.1800 2436.6400 1014.7800 2437.1200 ;
        RECT 1013.1800 2420.3200 1014.7800 2420.8000 ;
        RECT 1013.1800 2425.7600 1014.7800 2426.2400 ;
        RECT 1013.1800 2442.0800 1014.7800 2442.5600 ;
        RECT 1013.1800 2404.0000 1014.7800 2404.4800 ;
        RECT 1013.1800 2409.4400 1014.7800 2409.9200 ;
        RECT 1013.1800 2387.6800 1014.7800 2388.1600 ;
        RECT 1013.1800 2393.1200 1014.7800 2393.6000 ;
        RECT 1013.1800 2398.5600 1014.7800 2399.0400 ;
        RECT 1013.1800 2376.8000 1014.7800 2377.2800 ;
        RECT 1013.1800 2382.2400 1014.7800 2382.7200 ;
        RECT 1013.1800 2360.4800 1014.7800 2360.9600 ;
        RECT 1013.1800 2365.9200 1014.7800 2366.4000 ;
        RECT 1013.1800 2371.3600 1014.7800 2371.8400 ;
        RECT 1013.1800 2414.8800 1014.7800 2415.3600 ;
        RECT 1055.6000 2349.6000 1057.2000 2350.0800 ;
        RECT 1055.6000 2355.0400 1057.2000 2355.5200 ;
        RECT 1055.6000 2333.2800 1057.2000 2333.7600 ;
        RECT 1055.6000 2338.7200 1057.2000 2339.2000 ;
        RECT 1055.6000 2344.1600 1057.2000 2344.6400 ;
        RECT 1055.6000 2322.4000 1057.2000 2322.8800 ;
        RECT 1055.6000 2327.8400 1057.2000 2328.3200 ;
        RECT 1055.6000 2306.0800 1057.2000 2306.5600 ;
        RECT 1055.6000 2311.5200 1057.2000 2312.0000 ;
        RECT 1055.6000 2316.9600 1057.2000 2317.4400 ;
        RECT 1055.6000 2295.2000 1057.2000 2295.6800 ;
        RECT 1055.6000 2300.6400 1057.2000 2301.1200 ;
        RECT 1055.6000 2278.8800 1057.2000 2279.3600 ;
        RECT 1055.6000 2284.3200 1057.2000 2284.8000 ;
        RECT 1055.6000 2289.7600 1057.2000 2290.2400 ;
        RECT 1055.6000 2268.0000 1057.2000 2268.4800 ;
        RECT 1055.6000 2273.4400 1057.2000 2273.9200 ;
        RECT 1055.6000 2262.5600 1057.2000 2263.0400 ;
        RECT 1013.1800 2349.6000 1014.7800 2350.0800 ;
        RECT 1013.1800 2355.0400 1014.7800 2355.5200 ;
        RECT 1013.1800 2333.2800 1014.7800 2333.7600 ;
        RECT 1013.1800 2338.7200 1014.7800 2339.2000 ;
        RECT 1013.1800 2344.1600 1014.7800 2344.6400 ;
        RECT 1013.1800 2322.4000 1014.7800 2322.8800 ;
        RECT 1013.1800 2327.8400 1014.7800 2328.3200 ;
        RECT 1013.1800 2306.0800 1014.7800 2306.5600 ;
        RECT 1013.1800 2311.5200 1014.7800 2312.0000 ;
        RECT 1013.1800 2316.9600 1014.7800 2317.4400 ;
        RECT 1013.1800 2295.2000 1014.7800 2295.6800 ;
        RECT 1013.1800 2300.6400 1014.7800 2301.1200 ;
        RECT 1013.1800 2278.8800 1014.7800 2279.3600 ;
        RECT 1013.1800 2284.3200 1014.7800 2284.8000 ;
        RECT 1013.1800 2289.7600 1014.7800 2290.2400 ;
        RECT 1013.1800 2268.0000 1014.7800 2268.4800 ;
        RECT 1013.1800 2273.4400 1014.7800 2273.9200 ;
        RECT 1013.1800 2262.5600 1014.7800 2263.0400 ;
        RECT 1010.1200 2464.6500 1060.2600 2466.2500 ;
        RECT 1010.1200 2253.1500 1060.2600 2254.7500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 2250.2200 1014.7800 2251.8200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 2468.2600 1014.7800 2469.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 2250.2200 1057.2000 2251.8200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 2468.2600 1057.2000 2469.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2253.1500 1011.7200 2254.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2253.1500 1060.2600 2254.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2464.6500 1011.7200 2466.2500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2464.6500 1060.2600 2466.2500 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 2020.5800 1057.2000 2240.2200 ;
        RECT 1013.1800 2020.5800 1014.7800 2240.2200 ;
      LAYER met3 ;
        RECT 1055.6000 2228.7600 1057.2000 2229.2400 ;
        RECT 1055.6000 2217.8800 1057.2000 2218.3600 ;
        RECT 1055.6000 2223.3200 1057.2000 2223.8000 ;
        RECT 1055.6000 2201.5600 1057.2000 2202.0400 ;
        RECT 1055.6000 2207.0000 1057.2000 2207.4800 ;
        RECT 1055.6000 2190.6800 1057.2000 2191.1600 ;
        RECT 1055.6000 2196.1200 1057.2000 2196.6000 ;
        RECT 1055.6000 2212.4400 1057.2000 2212.9200 ;
        RECT 1055.6000 2174.3600 1057.2000 2174.8400 ;
        RECT 1055.6000 2179.8000 1057.2000 2180.2800 ;
        RECT 1055.6000 2158.0400 1057.2000 2158.5200 ;
        RECT 1055.6000 2163.4800 1057.2000 2163.9600 ;
        RECT 1055.6000 2168.9200 1057.2000 2169.4000 ;
        RECT 1055.6000 2147.1600 1057.2000 2147.6400 ;
        RECT 1055.6000 2152.6000 1057.2000 2153.0800 ;
        RECT 1055.6000 2130.8400 1057.2000 2131.3200 ;
        RECT 1055.6000 2136.2800 1057.2000 2136.7600 ;
        RECT 1055.6000 2141.7200 1057.2000 2142.2000 ;
        RECT 1055.6000 2185.2400 1057.2000 2185.7200 ;
        RECT 1013.1800 2228.7600 1014.7800 2229.2400 ;
        RECT 1013.1800 2217.8800 1014.7800 2218.3600 ;
        RECT 1013.1800 2223.3200 1014.7800 2223.8000 ;
        RECT 1013.1800 2201.5600 1014.7800 2202.0400 ;
        RECT 1013.1800 2207.0000 1014.7800 2207.4800 ;
        RECT 1013.1800 2190.6800 1014.7800 2191.1600 ;
        RECT 1013.1800 2196.1200 1014.7800 2196.6000 ;
        RECT 1013.1800 2212.4400 1014.7800 2212.9200 ;
        RECT 1013.1800 2174.3600 1014.7800 2174.8400 ;
        RECT 1013.1800 2179.8000 1014.7800 2180.2800 ;
        RECT 1013.1800 2158.0400 1014.7800 2158.5200 ;
        RECT 1013.1800 2163.4800 1014.7800 2163.9600 ;
        RECT 1013.1800 2168.9200 1014.7800 2169.4000 ;
        RECT 1013.1800 2147.1600 1014.7800 2147.6400 ;
        RECT 1013.1800 2152.6000 1014.7800 2153.0800 ;
        RECT 1013.1800 2130.8400 1014.7800 2131.3200 ;
        RECT 1013.1800 2136.2800 1014.7800 2136.7600 ;
        RECT 1013.1800 2141.7200 1014.7800 2142.2000 ;
        RECT 1013.1800 2185.2400 1014.7800 2185.7200 ;
        RECT 1055.6000 2119.9600 1057.2000 2120.4400 ;
        RECT 1055.6000 2125.4000 1057.2000 2125.8800 ;
        RECT 1055.6000 2103.6400 1057.2000 2104.1200 ;
        RECT 1055.6000 2109.0800 1057.2000 2109.5600 ;
        RECT 1055.6000 2114.5200 1057.2000 2115.0000 ;
        RECT 1055.6000 2092.7600 1057.2000 2093.2400 ;
        RECT 1055.6000 2098.2000 1057.2000 2098.6800 ;
        RECT 1055.6000 2076.4400 1057.2000 2076.9200 ;
        RECT 1055.6000 2081.8800 1057.2000 2082.3600 ;
        RECT 1055.6000 2087.3200 1057.2000 2087.8000 ;
        RECT 1055.6000 2065.5600 1057.2000 2066.0400 ;
        RECT 1055.6000 2071.0000 1057.2000 2071.4800 ;
        RECT 1055.6000 2049.2400 1057.2000 2049.7200 ;
        RECT 1055.6000 2054.6800 1057.2000 2055.1600 ;
        RECT 1055.6000 2060.1200 1057.2000 2060.6000 ;
        RECT 1055.6000 2038.3600 1057.2000 2038.8400 ;
        RECT 1055.6000 2043.8000 1057.2000 2044.2800 ;
        RECT 1055.6000 2032.9200 1057.2000 2033.4000 ;
        RECT 1013.1800 2119.9600 1014.7800 2120.4400 ;
        RECT 1013.1800 2125.4000 1014.7800 2125.8800 ;
        RECT 1013.1800 2103.6400 1014.7800 2104.1200 ;
        RECT 1013.1800 2109.0800 1014.7800 2109.5600 ;
        RECT 1013.1800 2114.5200 1014.7800 2115.0000 ;
        RECT 1013.1800 2092.7600 1014.7800 2093.2400 ;
        RECT 1013.1800 2098.2000 1014.7800 2098.6800 ;
        RECT 1013.1800 2076.4400 1014.7800 2076.9200 ;
        RECT 1013.1800 2081.8800 1014.7800 2082.3600 ;
        RECT 1013.1800 2087.3200 1014.7800 2087.8000 ;
        RECT 1013.1800 2065.5600 1014.7800 2066.0400 ;
        RECT 1013.1800 2071.0000 1014.7800 2071.4800 ;
        RECT 1013.1800 2049.2400 1014.7800 2049.7200 ;
        RECT 1013.1800 2054.6800 1014.7800 2055.1600 ;
        RECT 1013.1800 2060.1200 1014.7800 2060.6000 ;
        RECT 1013.1800 2038.3600 1014.7800 2038.8400 ;
        RECT 1013.1800 2043.8000 1014.7800 2044.2800 ;
        RECT 1013.1800 2032.9200 1014.7800 2033.4000 ;
        RECT 1010.1200 2235.0100 1060.2600 2236.6100 ;
        RECT 1010.1200 2023.5100 1060.2600 2025.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 2020.5800 1014.7800 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 2238.6200 1014.7800 2240.2200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 2020.5800 1057.2000 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 2238.6200 1057.2000 2240.2200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2023.5100 1011.7200 2025.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2023.5100 1060.2600 2025.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2235.0100 1011.7200 2236.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2235.0100 1060.2600 2236.6100 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 1790.9400 1057.2000 2010.5800 ;
        RECT 1013.1800 1790.9400 1014.7800 2010.5800 ;
      LAYER met3 ;
        RECT 1055.6000 1999.1200 1057.2000 1999.6000 ;
        RECT 1055.6000 1988.2400 1057.2000 1988.7200 ;
        RECT 1055.6000 1993.6800 1057.2000 1994.1600 ;
        RECT 1055.6000 1971.9200 1057.2000 1972.4000 ;
        RECT 1055.6000 1977.3600 1057.2000 1977.8400 ;
        RECT 1055.6000 1961.0400 1057.2000 1961.5200 ;
        RECT 1055.6000 1966.4800 1057.2000 1966.9600 ;
        RECT 1055.6000 1982.8000 1057.2000 1983.2800 ;
        RECT 1055.6000 1944.7200 1057.2000 1945.2000 ;
        RECT 1055.6000 1950.1600 1057.2000 1950.6400 ;
        RECT 1055.6000 1928.4000 1057.2000 1928.8800 ;
        RECT 1055.6000 1933.8400 1057.2000 1934.3200 ;
        RECT 1055.6000 1939.2800 1057.2000 1939.7600 ;
        RECT 1055.6000 1917.5200 1057.2000 1918.0000 ;
        RECT 1055.6000 1922.9600 1057.2000 1923.4400 ;
        RECT 1055.6000 1901.2000 1057.2000 1901.6800 ;
        RECT 1055.6000 1906.6400 1057.2000 1907.1200 ;
        RECT 1055.6000 1912.0800 1057.2000 1912.5600 ;
        RECT 1055.6000 1955.6000 1057.2000 1956.0800 ;
        RECT 1013.1800 1999.1200 1014.7800 1999.6000 ;
        RECT 1013.1800 1988.2400 1014.7800 1988.7200 ;
        RECT 1013.1800 1993.6800 1014.7800 1994.1600 ;
        RECT 1013.1800 1971.9200 1014.7800 1972.4000 ;
        RECT 1013.1800 1977.3600 1014.7800 1977.8400 ;
        RECT 1013.1800 1961.0400 1014.7800 1961.5200 ;
        RECT 1013.1800 1966.4800 1014.7800 1966.9600 ;
        RECT 1013.1800 1982.8000 1014.7800 1983.2800 ;
        RECT 1013.1800 1944.7200 1014.7800 1945.2000 ;
        RECT 1013.1800 1950.1600 1014.7800 1950.6400 ;
        RECT 1013.1800 1928.4000 1014.7800 1928.8800 ;
        RECT 1013.1800 1933.8400 1014.7800 1934.3200 ;
        RECT 1013.1800 1939.2800 1014.7800 1939.7600 ;
        RECT 1013.1800 1917.5200 1014.7800 1918.0000 ;
        RECT 1013.1800 1922.9600 1014.7800 1923.4400 ;
        RECT 1013.1800 1901.2000 1014.7800 1901.6800 ;
        RECT 1013.1800 1906.6400 1014.7800 1907.1200 ;
        RECT 1013.1800 1912.0800 1014.7800 1912.5600 ;
        RECT 1013.1800 1955.6000 1014.7800 1956.0800 ;
        RECT 1055.6000 1890.3200 1057.2000 1890.8000 ;
        RECT 1055.6000 1895.7600 1057.2000 1896.2400 ;
        RECT 1055.6000 1874.0000 1057.2000 1874.4800 ;
        RECT 1055.6000 1879.4400 1057.2000 1879.9200 ;
        RECT 1055.6000 1884.8800 1057.2000 1885.3600 ;
        RECT 1055.6000 1863.1200 1057.2000 1863.6000 ;
        RECT 1055.6000 1868.5600 1057.2000 1869.0400 ;
        RECT 1055.6000 1846.8000 1057.2000 1847.2800 ;
        RECT 1055.6000 1852.2400 1057.2000 1852.7200 ;
        RECT 1055.6000 1857.6800 1057.2000 1858.1600 ;
        RECT 1055.6000 1835.9200 1057.2000 1836.4000 ;
        RECT 1055.6000 1841.3600 1057.2000 1841.8400 ;
        RECT 1055.6000 1819.6000 1057.2000 1820.0800 ;
        RECT 1055.6000 1825.0400 1057.2000 1825.5200 ;
        RECT 1055.6000 1830.4800 1057.2000 1830.9600 ;
        RECT 1055.6000 1808.7200 1057.2000 1809.2000 ;
        RECT 1055.6000 1814.1600 1057.2000 1814.6400 ;
        RECT 1055.6000 1803.2800 1057.2000 1803.7600 ;
        RECT 1013.1800 1890.3200 1014.7800 1890.8000 ;
        RECT 1013.1800 1895.7600 1014.7800 1896.2400 ;
        RECT 1013.1800 1874.0000 1014.7800 1874.4800 ;
        RECT 1013.1800 1879.4400 1014.7800 1879.9200 ;
        RECT 1013.1800 1884.8800 1014.7800 1885.3600 ;
        RECT 1013.1800 1863.1200 1014.7800 1863.6000 ;
        RECT 1013.1800 1868.5600 1014.7800 1869.0400 ;
        RECT 1013.1800 1846.8000 1014.7800 1847.2800 ;
        RECT 1013.1800 1852.2400 1014.7800 1852.7200 ;
        RECT 1013.1800 1857.6800 1014.7800 1858.1600 ;
        RECT 1013.1800 1835.9200 1014.7800 1836.4000 ;
        RECT 1013.1800 1841.3600 1014.7800 1841.8400 ;
        RECT 1013.1800 1819.6000 1014.7800 1820.0800 ;
        RECT 1013.1800 1825.0400 1014.7800 1825.5200 ;
        RECT 1013.1800 1830.4800 1014.7800 1830.9600 ;
        RECT 1013.1800 1808.7200 1014.7800 1809.2000 ;
        RECT 1013.1800 1814.1600 1014.7800 1814.6400 ;
        RECT 1013.1800 1803.2800 1014.7800 1803.7600 ;
        RECT 1010.1200 2005.3700 1060.2600 2006.9700 ;
        RECT 1010.1200 1793.8700 1060.2600 1795.4700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1790.9400 1014.7800 1792.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 2008.9800 1014.7800 2010.5800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1790.9400 1057.2000 1792.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 2008.9800 1057.2000 2010.5800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1793.8700 1011.7200 1795.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1793.8700 1060.2600 1795.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2005.3700 1011.7200 2006.9700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2005.3700 1060.2600 2006.9700 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 1561.3000 1057.2000 1780.9400 ;
        RECT 1013.1800 1561.3000 1014.7800 1780.9400 ;
      LAYER met3 ;
        RECT 1055.6000 1769.4800 1057.2000 1769.9600 ;
        RECT 1055.6000 1758.6000 1057.2000 1759.0800 ;
        RECT 1055.6000 1764.0400 1057.2000 1764.5200 ;
        RECT 1055.6000 1742.2800 1057.2000 1742.7600 ;
        RECT 1055.6000 1747.7200 1057.2000 1748.2000 ;
        RECT 1055.6000 1731.4000 1057.2000 1731.8800 ;
        RECT 1055.6000 1736.8400 1057.2000 1737.3200 ;
        RECT 1055.6000 1753.1600 1057.2000 1753.6400 ;
        RECT 1055.6000 1715.0800 1057.2000 1715.5600 ;
        RECT 1055.6000 1720.5200 1057.2000 1721.0000 ;
        RECT 1055.6000 1698.7600 1057.2000 1699.2400 ;
        RECT 1055.6000 1704.2000 1057.2000 1704.6800 ;
        RECT 1055.6000 1709.6400 1057.2000 1710.1200 ;
        RECT 1055.6000 1687.8800 1057.2000 1688.3600 ;
        RECT 1055.6000 1693.3200 1057.2000 1693.8000 ;
        RECT 1055.6000 1671.5600 1057.2000 1672.0400 ;
        RECT 1055.6000 1677.0000 1057.2000 1677.4800 ;
        RECT 1055.6000 1682.4400 1057.2000 1682.9200 ;
        RECT 1055.6000 1725.9600 1057.2000 1726.4400 ;
        RECT 1013.1800 1769.4800 1014.7800 1769.9600 ;
        RECT 1013.1800 1758.6000 1014.7800 1759.0800 ;
        RECT 1013.1800 1764.0400 1014.7800 1764.5200 ;
        RECT 1013.1800 1742.2800 1014.7800 1742.7600 ;
        RECT 1013.1800 1747.7200 1014.7800 1748.2000 ;
        RECT 1013.1800 1731.4000 1014.7800 1731.8800 ;
        RECT 1013.1800 1736.8400 1014.7800 1737.3200 ;
        RECT 1013.1800 1753.1600 1014.7800 1753.6400 ;
        RECT 1013.1800 1715.0800 1014.7800 1715.5600 ;
        RECT 1013.1800 1720.5200 1014.7800 1721.0000 ;
        RECT 1013.1800 1698.7600 1014.7800 1699.2400 ;
        RECT 1013.1800 1704.2000 1014.7800 1704.6800 ;
        RECT 1013.1800 1709.6400 1014.7800 1710.1200 ;
        RECT 1013.1800 1687.8800 1014.7800 1688.3600 ;
        RECT 1013.1800 1693.3200 1014.7800 1693.8000 ;
        RECT 1013.1800 1671.5600 1014.7800 1672.0400 ;
        RECT 1013.1800 1677.0000 1014.7800 1677.4800 ;
        RECT 1013.1800 1682.4400 1014.7800 1682.9200 ;
        RECT 1013.1800 1725.9600 1014.7800 1726.4400 ;
        RECT 1055.6000 1660.6800 1057.2000 1661.1600 ;
        RECT 1055.6000 1666.1200 1057.2000 1666.6000 ;
        RECT 1055.6000 1644.3600 1057.2000 1644.8400 ;
        RECT 1055.6000 1649.8000 1057.2000 1650.2800 ;
        RECT 1055.6000 1655.2400 1057.2000 1655.7200 ;
        RECT 1055.6000 1633.4800 1057.2000 1633.9600 ;
        RECT 1055.6000 1638.9200 1057.2000 1639.4000 ;
        RECT 1055.6000 1617.1600 1057.2000 1617.6400 ;
        RECT 1055.6000 1622.6000 1057.2000 1623.0800 ;
        RECT 1055.6000 1628.0400 1057.2000 1628.5200 ;
        RECT 1055.6000 1606.2800 1057.2000 1606.7600 ;
        RECT 1055.6000 1611.7200 1057.2000 1612.2000 ;
        RECT 1055.6000 1589.9600 1057.2000 1590.4400 ;
        RECT 1055.6000 1595.4000 1057.2000 1595.8800 ;
        RECT 1055.6000 1600.8400 1057.2000 1601.3200 ;
        RECT 1055.6000 1579.0800 1057.2000 1579.5600 ;
        RECT 1055.6000 1584.5200 1057.2000 1585.0000 ;
        RECT 1055.6000 1573.6400 1057.2000 1574.1200 ;
        RECT 1013.1800 1660.6800 1014.7800 1661.1600 ;
        RECT 1013.1800 1666.1200 1014.7800 1666.6000 ;
        RECT 1013.1800 1644.3600 1014.7800 1644.8400 ;
        RECT 1013.1800 1649.8000 1014.7800 1650.2800 ;
        RECT 1013.1800 1655.2400 1014.7800 1655.7200 ;
        RECT 1013.1800 1633.4800 1014.7800 1633.9600 ;
        RECT 1013.1800 1638.9200 1014.7800 1639.4000 ;
        RECT 1013.1800 1617.1600 1014.7800 1617.6400 ;
        RECT 1013.1800 1622.6000 1014.7800 1623.0800 ;
        RECT 1013.1800 1628.0400 1014.7800 1628.5200 ;
        RECT 1013.1800 1606.2800 1014.7800 1606.7600 ;
        RECT 1013.1800 1611.7200 1014.7800 1612.2000 ;
        RECT 1013.1800 1589.9600 1014.7800 1590.4400 ;
        RECT 1013.1800 1595.4000 1014.7800 1595.8800 ;
        RECT 1013.1800 1600.8400 1014.7800 1601.3200 ;
        RECT 1013.1800 1579.0800 1014.7800 1579.5600 ;
        RECT 1013.1800 1584.5200 1014.7800 1585.0000 ;
        RECT 1013.1800 1573.6400 1014.7800 1574.1200 ;
        RECT 1010.1200 1775.7300 1060.2600 1777.3300 ;
        RECT 1010.1200 1564.2300 1060.2600 1565.8300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1561.3000 1014.7800 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1779.3400 1014.7800 1780.9400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1561.3000 1057.2000 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1779.3400 1057.2000 1780.9400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1564.2300 1011.7200 1565.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1564.2300 1060.2600 1565.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1775.7300 1011.7200 1777.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1775.7300 1060.2600 1777.3300 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 1331.6600 1057.2000 1551.3000 ;
        RECT 1013.1800 1331.6600 1014.7800 1551.3000 ;
      LAYER met3 ;
        RECT 1055.6000 1539.8400 1057.2000 1540.3200 ;
        RECT 1055.6000 1528.9600 1057.2000 1529.4400 ;
        RECT 1055.6000 1534.4000 1057.2000 1534.8800 ;
        RECT 1055.6000 1512.6400 1057.2000 1513.1200 ;
        RECT 1055.6000 1518.0800 1057.2000 1518.5600 ;
        RECT 1055.6000 1501.7600 1057.2000 1502.2400 ;
        RECT 1055.6000 1507.2000 1057.2000 1507.6800 ;
        RECT 1055.6000 1523.5200 1057.2000 1524.0000 ;
        RECT 1055.6000 1485.4400 1057.2000 1485.9200 ;
        RECT 1055.6000 1490.8800 1057.2000 1491.3600 ;
        RECT 1055.6000 1469.1200 1057.2000 1469.6000 ;
        RECT 1055.6000 1474.5600 1057.2000 1475.0400 ;
        RECT 1055.6000 1480.0000 1057.2000 1480.4800 ;
        RECT 1055.6000 1458.2400 1057.2000 1458.7200 ;
        RECT 1055.6000 1463.6800 1057.2000 1464.1600 ;
        RECT 1055.6000 1441.9200 1057.2000 1442.4000 ;
        RECT 1055.6000 1447.3600 1057.2000 1447.8400 ;
        RECT 1055.6000 1452.8000 1057.2000 1453.2800 ;
        RECT 1055.6000 1496.3200 1057.2000 1496.8000 ;
        RECT 1013.1800 1539.8400 1014.7800 1540.3200 ;
        RECT 1013.1800 1528.9600 1014.7800 1529.4400 ;
        RECT 1013.1800 1534.4000 1014.7800 1534.8800 ;
        RECT 1013.1800 1512.6400 1014.7800 1513.1200 ;
        RECT 1013.1800 1518.0800 1014.7800 1518.5600 ;
        RECT 1013.1800 1501.7600 1014.7800 1502.2400 ;
        RECT 1013.1800 1507.2000 1014.7800 1507.6800 ;
        RECT 1013.1800 1523.5200 1014.7800 1524.0000 ;
        RECT 1013.1800 1485.4400 1014.7800 1485.9200 ;
        RECT 1013.1800 1490.8800 1014.7800 1491.3600 ;
        RECT 1013.1800 1469.1200 1014.7800 1469.6000 ;
        RECT 1013.1800 1474.5600 1014.7800 1475.0400 ;
        RECT 1013.1800 1480.0000 1014.7800 1480.4800 ;
        RECT 1013.1800 1458.2400 1014.7800 1458.7200 ;
        RECT 1013.1800 1463.6800 1014.7800 1464.1600 ;
        RECT 1013.1800 1441.9200 1014.7800 1442.4000 ;
        RECT 1013.1800 1447.3600 1014.7800 1447.8400 ;
        RECT 1013.1800 1452.8000 1014.7800 1453.2800 ;
        RECT 1013.1800 1496.3200 1014.7800 1496.8000 ;
        RECT 1055.6000 1431.0400 1057.2000 1431.5200 ;
        RECT 1055.6000 1436.4800 1057.2000 1436.9600 ;
        RECT 1055.6000 1414.7200 1057.2000 1415.2000 ;
        RECT 1055.6000 1420.1600 1057.2000 1420.6400 ;
        RECT 1055.6000 1425.6000 1057.2000 1426.0800 ;
        RECT 1055.6000 1403.8400 1057.2000 1404.3200 ;
        RECT 1055.6000 1409.2800 1057.2000 1409.7600 ;
        RECT 1055.6000 1387.5200 1057.2000 1388.0000 ;
        RECT 1055.6000 1392.9600 1057.2000 1393.4400 ;
        RECT 1055.6000 1398.4000 1057.2000 1398.8800 ;
        RECT 1055.6000 1376.6400 1057.2000 1377.1200 ;
        RECT 1055.6000 1382.0800 1057.2000 1382.5600 ;
        RECT 1055.6000 1360.3200 1057.2000 1360.8000 ;
        RECT 1055.6000 1365.7600 1057.2000 1366.2400 ;
        RECT 1055.6000 1371.2000 1057.2000 1371.6800 ;
        RECT 1055.6000 1349.4400 1057.2000 1349.9200 ;
        RECT 1055.6000 1354.8800 1057.2000 1355.3600 ;
        RECT 1055.6000 1344.0000 1057.2000 1344.4800 ;
        RECT 1013.1800 1431.0400 1014.7800 1431.5200 ;
        RECT 1013.1800 1436.4800 1014.7800 1436.9600 ;
        RECT 1013.1800 1414.7200 1014.7800 1415.2000 ;
        RECT 1013.1800 1420.1600 1014.7800 1420.6400 ;
        RECT 1013.1800 1425.6000 1014.7800 1426.0800 ;
        RECT 1013.1800 1403.8400 1014.7800 1404.3200 ;
        RECT 1013.1800 1409.2800 1014.7800 1409.7600 ;
        RECT 1013.1800 1387.5200 1014.7800 1388.0000 ;
        RECT 1013.1800 1392.9600 1014.7800 1393.4400 ;
        RECT 1013.1800 1398.4000 1014.7800 1398.8800 ;
        RECT 1013.1800 1376.6400 1014.7800 1377.1200 ;
        RECT 1013.1800 1382.0800 1014.7800 1382.5600 ;
        RECT 1013.1800 1360.3200 1014.7800 1360.8000 ;
        RECT 1013.1800 1365.7600 1014.7800 1366.2400 ;
        RECT 1013.1800 1371.2000 1014.7800 1371.6800 ;
        RECT 1013.1800 1349.4400 1014.7800 1349.9200 ;
        RECT 1013.1800 1354.8800 1014.7800 1355.3600 ;
        RECT 1013.1800 1344.0000 1014.7800 1344.4800 ;
        RECT 1010.1200 1546.0900 1060.2600 1547.6900 ;
        RECT 1010.1200 1334.5900 1060.2600 1336.1900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1331.6600 1014.7800 1333.2600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1549.7000 1014.7800 1551.3000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1331.6600 1057.2000 1333.2600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1549.7000 1057.2000 1551.3000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1334.5900 1011.7200 1336.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1334.5900 1060.2600 1336.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1546.0900 1011.7200 1547.6900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1546.0900 1060.2600 1547.6900 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 1102.0200 1057.2000 1321.6600 ;
        RECT 1013.1800 1102.0200 1014.7800 1321.6600 ;
      LAYER met3 ;
        RECT 1055.6000 1310.2000 1057.2000 1310.6800 ;
        RECT 1055.6000 1299.3200 1057.2000 1299.8000 ;
        RECT 1055.6000 1304.7600 1057.2000 1305.2400 ;
        RECT 1055.6000 1283.0000 1057.2000 1283.4800 ;
        RECT 1055.6000 1288.4400 1057.2000 1288.9200 ;
        RECT 1055.6000 1272.1200 1057.2000 1272.6000 ;
        RECT 1055.6000 1277.5600 1057.2000 1278.0400 ;
        RECT 1055.6000 1293.8800 1057.2000 1294.3600 ;
        RECT 1055.6000 1255.8000 1057.2000 1256.2800 ;
        RECT 1055.6000 1261.2400 1057.2000 1261.7200 ;
        RECT 1055.6000 1239.4800 1057.2000 1239.9600 ;
        RECT 1055.6000 1244.9200 1057.2000 1245.4000 ;
        RECT 1055.6000 1250.3600 1057.2000 1250.8400 ;
        RECT 1055.6000 1228.6000 1057.2000 1229.0800 ;
        RECT 1055.6000 1234.0400 1057.2000 1234.5200 ;
        RECT 1055.6000 1212.2800 1057.2000 1212.7600 ;
        RECT 1055.6000 1217.7200 1057.2000 1218.2000 ;
        RECT 1055.6000 1223.1600 1057.2000 1223.6400 ;
        RECT 1055.6000 1266.6800 1057.2000 1267.1600 ;
        RECT 1013.1800 1310.2000 1014.7800 1310.6800 ;
        RECT 1013.1800 1299.3200 1014.7800 1299.8000 ;
        RECT 1013.1800 1304.7600 1014.7800 1305.2400 ;
        RECT 1013.1800 1283.0000 1014.7800 1283.4800 ;
        RECT 1013.1800 1288.4400 1014.7800 1288.9200 ;
        RECT 1013.1800 1272.1200 1014.7800 1272.6000 ;
        RECT 1013.1800 1277.5600 1014.7800 1278.0400 ;
        RECT 1013.1800 1293.8800 1014.7800 1294.3600 ;
        RECT 1013.1800 1255.8000 1014.7800 1256.2800 ;
        RECT 1013.1800 1261.2400 1014.7800 1261.7200 ;
        RECT 1013.1800 1239.4800 1014.7800 1239.9600 ;
        RECT 1013.1800 1244.9200 1014.7800 1245.4000 ;
        RECT 1013.1800 1250.3600 1014.7800 1250.8400 ;
        RECT 1013.1800 1228.6000 1014.7800 1229.0800 ;
        RECT 1013.1800 1234.0400 1014.7800 1234.5200 ;
        RECT 1013.1800 1212.2800 1014.7800 1212.7600 ;
        RECT 1013.1800 1217.7200 1014.7800 1218.2000 ;
        RECT 1013.1800 1223.1600 1014.7800 1223.6400 ;
        RECT 1013.1800 1266.6800 1014.7800 1267.1600 ;
        RECT 1055.6000 1201.4000 1057.2000 1201.8800 ;
        RECT 1055.6000 1206.8400 1057.2000 1207.3200 ;
        RECT 1055.6000 1185.0800 1057.2000 1185.5600 ;
        RECT 1055.6000 1190.5200 1057.2000 1191.0000 ;
        RECT 1055.6000 1195.9600 1057.2000 1196.4400 ;
        RECT 1055.6000 1174.2000 1057.2000 1174.6800 ;
        RECT 1055.6000 1179.6400 1057.2000 1180.1200 ;
        RECT 1055.6000 1157.8800 1057.2000 1158.3600 ;
        RECT 1055.6000 1163.3200 1057.2000 1163.8000 ;
        RECT 1055.6000 1168.7600 1057.2000 1169.2400 ;
        RECT 1055.6000 1147.0000 1057.2000 1147.4800 ;
        RECT 1055.6000 1152.4400 1057.2000 1152.9200 ;
        RECT 1055.6000 1130.6800 1057.2000 1131.1600 ;
        RECT 1055.6000 1136.1200 1057.2000 1136.6000 ;
        RECT 1055.6000 1141.5600 1057.2000 1142.0400 ;
        RECT 1055.6000 1119.8000 1057.2000 1120.2800 ;
        RECT 1055.6000 1125.2400 1057.2000 1125.7200 ;
        RECT 1055.6000 1114.3600 1057.2000 1114.8400 ;
        RECT 1013.1800 1201.4000 1014.7800 1201.8800 ;
        RECT 1013.1800 1206.8400 1014.7800 1207.3200 ;
        RECT 1013.1800 1185.0800 1014.7800 1185.5600 ;
        RECT 1013.1800 1190.5200 1014.7800 1191.0000 ;
        RECT 1013.1800 1195.9600 1014.7800 1196.4400 ;
        RECT 1013.1800 1174.2000 1014.7800 1174.6800 ;
        RECT 1013.1800 1179.6400 1014.7800 1180.1200 ;
        RECT 1013.1800 1157.8800 1014.7800 1158.3600 ;
        RECT 1013.1800 1163.3200 1014.7800 1163.8000 ;
        RECT 1013.1800 1168.7600 1014.7800 1169.2400 ;
        RECT 1013.1800 1147.0000 1014.7800 1147.4800 ;
        RECT 1013.1800 1152.4400 1014.7800 1152.9200 ;
        RECT 1013.1800 1130.6800 1014.7800 1131.1600 ;
        RECT 1013.1800 1136.1200 1014.7800 1136.6000 ;
        RECT 1013.1800 1141.5600 1014.7800 1142.0400 ;
        RECT 1013.1800 1119.8000 1014.7800 1120.2800 ;
        RECT 1013.1800 1125.2400 1014.7800 1125.7200 ;
        RECT 1013.1800 1114.3600 1014.7800 1114.8400 ;
        RECT 1010.1200 1316.4500 1060.2600 1318.0500 ;
        RECT 1010.1200 1104.9500 1060.2600 1106.5500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1102.0200 1014.7800 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1320.0600 1014.7800 1321.6600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1102.0200 1057.2000 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1320.0600 1057.2000 1321.6600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1104.9500 1011.7200 1106.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1104.9500 1060.2600 1106.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1316.4500 1011.7200 1318.0500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1316.4500 1060.2600 1318.0500 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 872.3800 1057.2000 1092.0200 ;
        RECT 1013.1800 872.3800 1014.7800 1092.0200 ;
      LAYER met3 ;
        RECT 1055.6000 1080.5600 1057.2000 1081.0400 ;
        RECT 1055.6000 1069.6800 1057.2000 1070.1600 ;
        RECT 1055.6000 1075.1200 1057.2000 1075.6000 ;
        RECT 1055.6000 1053.3600 1057.2000 1053.8400 ;
        RECT 1055.6000 1058.8000 1057.2000 1059.2800 ;
        RECT 1055.6000 1042.4800 1057.2000 1042.9600 ;
        RECT 1055.6000 1047.9200 1057.2000 1048.4000 ;
        RECT 1055.6000 1064.2400 1057.2000 1064.7200 ;
        RECT 1055.6000 1026.1600 1057.2000 1026.6400 ;
        RECT 1055.6000 1031.6000 1057.2000 1032.0800 ;
        RECT 1055.6000 1009.8400 1057.2000 1010.3200 ;
        RECT 1055.6000 1015.2800 1057.2000 1015.7600 ;
        RECT 1055.6000 1020.7200 1057.2000 1021.2000 ;
        RECT 1055.6000 998.9600 1057.2000 999.4400 ;
        RECT 1055.6000 1004.4000 1057.2000 1004.8800 ;
        RECT 1055.6000 982.6400 1057.2000 983.1200 ;
        RECT 1055.6000 988.0800 1057.2000 988.5600 ;
        RECT 1055.6000 993.5200 1057.2000 994.0000 ;
        RECT 1055.6000 1037.0400 1057.2000 1037.5200 ;
        RECT 1013.1800 1080.5600 1014.7800 1081.0400 ;
        RECT 1013.1800 1069.6800 1014.7800 1070.1600 ;
        RECT 1013.1800 1075.1200 1014.7800 1075.6000 ;
        RECT 1013.1800 1053.3600 1014.7800 1053.8400 ;
        RECT 1013.1800 1058.8000 1014.7800 1059.2800 ;
        RECT 1013.1800 1042.4800 1014.7800 1042.9600 ;
        RECT 1013.1800 1047.9200 1014.7800 1048.4000 ;
        RECT 1013.1800 1064.2400 1014.7800 1064.7200 ;
        RECT 1013.1800 1026.1600 1014.7800 1026.6400 ;
        RECT 1013.1800 1031.6000 1014.7800 1032.0800 ;
        RECT 1013.1800 1009.8400 1014.7800 1010.3200 ;
        RECT 1013.1800 1015.2800 1014.7800 1015.7600 ;
        RECT 1013.1800 1020.7200 1014.7800 1021.2000 ;
        RECT 1013.1800 998.9600 1014.7800 999.4400 ;
        RECT 1013.1800 1004.4000 1014.7800 1004.8800 ;
        RECT 1013.1800 982.6400 1014.7800 983.1200 ;
        RECT 1013.1800 988.0800 1014.7800 988.5600 ;
        RECT 1013.1800 993.5200 1014.7800 994.0000 ;
        RECT 1013.1800 1037.0400 1014.7800 1037.5200 ;
        RECT 1055.6000 971.7600 1057.2000 972.2400 ;
        RECT 1055.6000 977.2000 1057.2000 977.6800 ;
        RECT 1055.6000 955.4400 1057.2000 955.9200 ;
        RECT 1055.6000 960.8800 1057.2000 961.3600 ;
        RECT 1055.6000 966.3200 1057.2000 966.8000 ;
        RECT 1055.6000 944.5600 1057.2000 945.0400 ;
        RECT 1055.6000 950.0000 1057.2000 950.4800 ;
        RECT 1055.6000 928.2400 1057.2000 928.7200 ;
        RECT 1055.6000 933.6800 1057.2000 934.1600 ;
        RECT 1055.6000 939.1200 1057.2000 939.6000 ;
        RECT 1055.6000 917.3600 1057.2000 917.8400 ;
        RECT 1055.6000 922.8000 1057.2000 923.2800 ;
        RECT 1055.6000 901.0400 1057.2000 901.5200 ;
        RECT 1055.6000 906.4800 1057.2000 906.9600 ;
        RECT 1055.6000 911.9200 1057.2000 912.4000 ;
        RECT 1055.6000 890.1600 1057.2000 890.6400 ;
        RECT 1055.6000 895.6000 1057.2000 896.0800 ;
        RECT 1055.6000 884.7200 1057.2000 885.2000 ;
        RECT 1013.1800 971.7600 1014.7800 972.2400 ;
        RECT 1013.1800 977.2000 1014.7800 977.6800 ;
        RECT 1013.1800 955.4400 1014.7800 955.9200 ;
        RECT 1013.1800 960.8800 1014.7800 961.3600 ;
        RECT 1013.1800 966.3200 1014.7800 966.8000 ;
        RECT 1013.1800 944.5600 1014.7800 945.0400 ;
        RECT 1013.1800 950.0000 1014.7800 950.4800 ;
        RECT 1013.1800 928.2400 1014.7800 928.7200 ;
        RECT 1013.1800 933.6800 1014.7800 934.1600 ;
        RECT 1013.1800 939.1200 1014.7800 939.6000 ;
        RECT 1013.1800 917.3600 1014.7800 917.8400 ;
        RECT 1013.1800 922.8000 1014.7800 923.2800 ;
        RECT 1013.1800 901.0400 1014.7800 901.5200 ;
        RECT 1013.1800 906.4800 1014.7800 906.9600 ;
        RECT 1013.1800 911.9200 1014.7800 912.4000 ;
        RECT 1013.1800 890.1600 1014.7800 890.6400 ;
        RECT 1013.1800 895.6000 1014.7800 896.0800 ;
        RECT 1013.1800 884.7200 1014.7800 885.2000 ;
        RECT 1010.1200 1086.8100 1060.2600 1088.4100 ;
        RECT 1010.1200 875.3100 1060.2600 876.9100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 872.3800 1014.7800 873.9800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 1090.4200 1014.7800 1092.0200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 872.3800 1057.2000 873.9800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 1090.4200 1057.2000 1092.0200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 875.3100 1011.7200 876.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 875.3100 1060.2600 876.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1086.8100 1011.7200 1088.4100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1086.8100 1060.2600 1088.4100 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 642.7400 1057.2000 862.3800 ;
        RECT 1013.1800 642.7400 1014.7800 862.3800 ;
      LAYER met3 ;
        RECT 1055.6000 850.9200 1057.2000 851.4000 ;
        RECT 1055.6000 840.0400 1057.2000 840.5200 ;
        RECT 1055.6000 845.4800 1057.2000 845.9600 ;
        RECT 1055.6000 823.7200 1057.2000 824.2000 ;
        RECT 1055.6000 829.1600 1057.2000 829.6400 ;
        RECT 1055.6000 812.8400 1057.2000 813.3200 ;
        RECT 1055.6000 818.2800 1057.2000 818.7600 ;
        RECT 1055.6000 834.6000 1057.2000 835.0800 ;
        RECT 1055.6000 796.5200 1057.2000 797.0000 ;
        RECT 1055.6000 801.9600 1057.2000 802.4400 ;
        RECT 1055.6000 780.2000 1057.2000 780.6800 ;
        RECT 1055.6000 785.6400 1057.2000 786.1200 ;
        RECT 1055.6000 791.0800 1057.2000 791.5600 ;
        RECT 1055.6000 769.3200 1057.2000 769.8000 ;
        RECT 1055.6000 774.7600 1057.2000 775.2400 ;
        RECT 1055.6000 753.0000 1057.2000 753.4800 ;
        RECT 1055.6000 758.4400 1057.2000 758.9200 ;
        RECT 1055.6000 763.8800 1057.2000 764.3600 ;
        RECT 1055.6000 807.4000 1057.2000 807.8800 ;
        RECT 1013.1800 850.9200 1014.7800 851.4000 ;
        RECT 1013.1800 840.0400 1014.7800 840.5200 ;
        RECT 1013.1800 845.4800 1014.7800 845.9600 ;
        RECT 1013.1800 823.7200 1014.7800 824.2000 ;
        RECT 1013.1800 829.1600 1014.7800 829.6400 ;
        RECT 1013.1800 812.8400 1014.7800 813.3200 ;
        RECT 1013.1800 818.2800 1014.7800 818.7600 ;
        RECT 1013.1800 834.6000 1014.7800 835.0800 ;
        RECT 1013.1800 796.5200 1014.7800 797.0000 ;
        RECT 1013.1800 801.9600 1014.7800 802.4400 ;
        RECT 1013.1800 780.2000 1014.7800 780.6800 ;
        RECT 1013.1800 785.6400 1014.7800 786.1200 ;
        RECT 1013.1800 791.0800 1014.7800 791.5600 ;
        RECT 1013.1800 769.3200 1014.7800 769.8000 ;
        RECT 1013.1800 774.7600 1014.7800 775.2400 ;
        RECT 1013.1800 753.0000 1014.7800 753.4800 ;
        RECT 1013.1800 758.4400 1014.7800 758.9200 ;
        RECT 1013.1800 763.8800 1014.7800 764.3600 ;
        RECT 1013.1800 807.4000 1014.7800 807.8800 ;
        RECT 1055.6000 742.1200 1057.2000 742.6000 ;
        RECT 1055.6000 747.5600 1057.2000 748.0400 ;
        RECT 1055.6000 725.8000 1057.2000 726.2800 ;
        RECT 1055.6000 731.2400 1057.2000 731.7200 ;
        RECT 1055.6000 736.6800 1057.2000 737.1600 ;
        RECT 1055.6000 714.9200 1057.2000 715.4000 ;
        RECT 1055.6000 720.3600 1057.2000 720.8400 ;
        RECT 1055.6000 698.6000 1057.2000 699.0800 ;
        RECT 1055.6000 704.0400 1057.2000 704.5200 ;
        RECT 1055.6000 709.4800 1057.2000 709.9600 ;
        RECT 1055.6000 687.7200 1057.2000 688.2000 ;
        RECT 1055.6000 693.1600 1057.2000 693.6400 ;
        RECT 1055.6000 671.4000 1057.2000 671.8800 ;
        RECT 1055.6000 676.8400 1057.2000 677.3200 ;
        RECT 1055.6000 682.2800 1057.2000 682.7600 ;
        RECT 1055.6000 660.5200 1057.2000 661.0000 ;
        RECT 1055.6000 665.9600 1057.2000 666.4400 ;
        RECT 1055.6000 655.0800 1057.2000 655.5600 ;
        RECT 1013.1800 742.1200 1014.7800 742.6000 ;
        RECT 1013.1800 747.5600 1014.7800 748.0400 ;
        RECT 1013.1800 725.8000 1014.7800 726.2800 ;
        RECT 1013.1800 731.2400 1014.7800 731.7200 ;
        RECT 1013.1800 736.6800 1014.7800 737.1600 ;
        RECT 1013.1800 714.9200 1014.7800 715.4000 ;
        RECT 1013.1800 720.3600 1014.7800 720.8400 ;
        RECT 1013.1800 698.6000 1014.7800 699.0800 ;
        RECT 1013.1800 704.0400 1014.7800 704.5200 ;
        RECT 1013.1800 709.4800 1014.7800 709.9600 ;
        RECT 1013.1800 687.7200 1014.7800 688.2000 ;
        RECT 1013.1800 693.1600 1014.7800 693.6400 ;
        RECT 1013.1800 671.4000 1014.7800 671.8800 ;
        RECT 1013.1800 676.8400 1014.7800 677.3200 ;
        RECT 1013.1800 682.2800 1014.7800 682.7600 ;
        RECT 1013.1800 660.5200 1014.7800 661.0000 ;
        RECT 1013.1800 665.9600 1014.7800 666.4400 ;
        RECT 1013.1800 655.0800 1014.7800 655.5600 ;
        RECT 1010.1200 857.1700 1060.2600 858.7700 ;
        RECT 1010.1200 645.6700 1060.2600 647.2700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 642.7400 1014.7800 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 860.7800 1014.7800 862.3800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 642.7400 1057.2000 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 860.7800 1057.2000 862.3800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 645.6700 1011.7200 647.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 645.6700 1060.2600 647.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 857.1700 1011.7200 858.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 857.1700 1060.2600 858.7700 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1055.6000 413.1000 1057.2000 632.7400 ;
        RECT 1013.1800 413.1000 1014.7800 632.7400 ;
      LAYER met3 ;
        RECT 1055.6000 621.2800 1057.2000 621.7600 ;
        RECT 1055.6000 610.4000 1057.2000 610.8800 ;
        RECT 1055.6000 615.8400 1057.2000 616.3200 ;
        RECT 1055.6000 594.0800 1057.2000 594.5600 ;
        RECT 1055.6000 599.5200 1057.2000 600.0000 ;
        RECT 1055.6000 583.2000 1057.2000 583.6800 ;
        RECT 1055.6000 588.6400 1057.2000 589.1200 ;
        RECT 1055.6000 604.9600 1057.2000 605.4400 ;
        RECT 1055.6000 566.8800 1057.2000 567.3600 ;
        RECT 1055.6000 572.3200 1057.2000 572.8000 ;
        RECT 1055.6000 550.5600 1057.2000 551.0400 ;
        RECT 1055.6000 556.0000 1057.2000 556.4800 ;
        RECT 1055.6000 561.4400 1057.2000 561.9200 ;
        RECT 1055.6000 539.6800 1057.2000 540.1600 ;
        RECT 1055.6000 545.1200 1057.2000 545.6000 ;
        RECT 1055.6000 523.3600 1057.2000 523.8400 ;
        RECT 1055.6000 528.8000 1057.2000 529.2800 ;
        RECT 1055.6000 534.2400 1057.2000 534.7200 ;
        RECT 1055.6000 577.7600 1057.2000 578.2400 ;
        RECT 1013.1800 621.2800 1014.7800 621.7600 ;
        RECT 1013.1800 610.4000 1014.7800 610.8800 ;
        RECT 1013.1800 615.8400 1014.7800 616.3200 ;
        RECT 1013.1800 594.0800 1014.7800 594.5600 ;
        RECT 1013.1800 599.5200 1014.7800 600.0000 ;
        RECT 1013.1800 583.2000 1014.7800 583.6800 ;
        RECT 1013.1800 588.6400 1014.7800 589.1200 ;
        RECT 1013.1800 604.9600 1014.7800 605.4400 ;
        RECT 1013.1800 566.8800 1014.7800 567.3600 ;
        RECT 1013.1800 572.3200 1014.7800 572.8000 ;
        RECT 1013.1800 550.5600 1014.7800 551.0400 ;
        RECT 1013.1800 556.0000 1014.7800 556.4800 ;
        RECT 1013.1800 561.4400 1014.7800 561.9200 ;
        RECT 1013.1800 539.6800 1014.7800 540.1600 ;
        RECT 1013.1800 545.1200 1014.7800 545.6000 ;
        RECT 1013.1800 523.3600 1014.7800 523.8400 ;
        RECT 1013.1800 528.8000 1014.7800 529.2800 ;
        RECT 1013.1800 534.2400 1014.7800 534.7200 ;
        RECT 1013.1800 577.7600 1014.7800 578.2400 ;
        RECT 1055.6000 512.4800 1057.2000 512.9600 ;
        RECT 1055.6000 517.9200 1057.2000 518.4000 ;
        RECT 1055.6000 496.1600 1057.2000 496.6400 ;
        RECT 1055.6000 501.6000 1057.2000 502.0800 ;
        RECT 1055.6000 507.0400 1057.2000 507.5200 ;
        RECT 1055.6000 485.2800 1057.2000 485.7600 ;
        RECT 1055.6000 490.7200 1057.2000 491.2000 ;
        RECT 1055.6000 468.9600 1057.2000 469.4400 ;
        RECT 1055.6000 474.4000 1057.2000 474.8800 ;
        RECT 1055.6000 479.8400 1057.2000 480.3200 ;
        RECT 1055.6000 458.0800 1057.2000 458.5600 ;
        RECT 1055.6000 463.5200 1057.2000 464.0000 ;
        RECT 1055.6000 441.7600 1057.2000 442.2400 ;
        RECT 1055.6000 447.2000 1057.2000 447.6800 ;
        RECT 1055.6000 452.6400 1057.2000 453.1200 ;
        RECT 1055.6000 430.8800 1057.2000 431.3600 ;
        RECT 1055.6000 436.3200 1057.2000 436.8000 ;
        RECT 1055.6000 425.4400 1057.2000 425.9200 ;
        RECT 1013.1800 512.4800 1014.7800 512.9600 ;
        RECT 1013.1800 517.9200 1014.7800 518.4000 ;
        RECT 1013.1800 496.1600 1014.7800 496.6400 ;
        RECT 1013.1800 501.6000 1014.7800 502.0800 ;
        RECT 1013.1800 507.0400 1014.7800 507.5200 ;
        RECT 1013.1800 485.2800 1014.7800 485.7600 ;
        RECT 1013.1800 490.7200 1014.7800 491.2000 ;
        RECT 1013.1800 468.9600 1014.7800 469.4400 ;
        RECT 1013.1800 474.4000 1014.7800 474.8800 ;
        RECT 1013.1800 479.8400 1014.7800 480.3200 ;
        RECT 1013.1800 458.0800 1014.7800 458.5600 ;
        RECT 1013.1800 463.5200 1014.7800 464.0000 ;
        RECT 1013.1800 441.7600 1014.7800 442.2400 ;
        RECT 1013.1800 447.2000 1014.7800 447.6800 ;
        RECT 1013.1800 452.6400 1014.7800 453.1200 ;
        RECT 1013.1800 430.8800 1014.7800 431.3600 ;
        RECT 1013.1800 436.3200 1014.7800 436.8000 ;
        RECT 1013.1800 425.4400 1014.7800 425.9200 ;
        RECT 1010.1200 627.5300 1060.2600 629.1300 ;
        RECT 1010.1200 416.0300 1060.2600 417.6300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 413.1000 1014.7800 414.7000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1013.1800 631.1400 1014.7800 632.7400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 413.1000 1057.2000 414.7000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.6000 631.1400 1057.2000 632.7400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 416.0300 1011.7200 417.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 416.0300 1060.2600 417.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 627.5300 1011.7200 629.1300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 627.5300 1060.2600 629.1300 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'N_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1073.1800 2479.6000 1074.7800 2509.8600 ;
        RECT 1275.6800 2479.6000 1277.2800 2509.8600 ;
      LAYER met3 ;
        RECT 1275.6800 2500.1000 1277.2800 2500.5800 ;
        RECT 1073.1800 2500.1000 1074.7800 2500.5800 ;
        RECT 1275.6800 2489.2200 1277.2800 2489.7000 ;
        RECT 1073.1800 2489.2200 1074.7800 2489.7000 ;
        RECT 1275.6800 2494.6600 1277.2800 2495.1400 ;
        RECT 1073.1800 2494.6600 1074.7800 2495.1400 ;
        RECT 1070.1200 2505.5000 1280.3400 2507.1000 ;
        RECT 1070.1200 2481.1700 1280.3400 2482.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.1800 2479.6000 1074.7800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.1800 2508.2600 1074.7800 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.6800 2479.6000 1277.2800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.6800 2508.2600 1277.2800 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.1200 2481.1700 1071.7200 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.7400 2481.1700 1280.3400 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.1200 2505.5000 1071.7200 2507.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.7400 2505.5000 1280.3400 2507.1000 ;
    END
# end of P/G pin shape extracted from block 'N_term_DSP'


# P/G pin shape extracted from block 'S_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1073.3200 143.2000 1074.9200 173.4600 ;
        RECT 1275.8200 143.2000 1277.4200 173.4600 ;
      LAYER met3 ;
        RECT 1275.8200 163.7000 1277.4200 164.1800 ;
        RECT 1073.3200 163.7000 1074.9200 164.1800 ;
        RECT 1275.8200 152.8200 1277.4200 153.3000 ;
        RECT 1073.3200 152.8200 1074.9200 153.3000 ;
        RECT 1275.8200 158.2600 1277.4200 158.7400 ;
        RECT 1073.3200 158.2600 1074.9200 158.7400 ;
        RECT 1070.2600 169.1000 1280.4800 170.7000 ;
        RECT 1070.2600 144.7700 1280.4800 146.3700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.3200 143.2000 1074.9200 144.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.3200 171.8600 1074.9200 173.4600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.8200 143.2000 1277.4200 144.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.8200 171.8600 1277.4200 173.4600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 144.7700 1071.8600 146.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 144.7700 1280.4800 146.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 169.1000 1071.8600 170.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 169.1000 1280.4800 170.7000 ;
    END
# end of P/G pin shape extracted from block 'S_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1073.2200 2020.5800 1074.8200 2470.4000 ;
        RECT 1275.9200 2020.5800 1277.5200 2470.4000 ;
        RECT 1080.3800 2023.4100 1081.9800 2467.4000 ;
        RECT 1125.3800 2023.4100 1126.9800 2467.4000 ;
        RECT 1170.3800 2023.4100 1171.9800 2467.4000 ;
        RECT 1215.3800 2023.4100 1216.9800 2467.4000 ;
        RECT 1260.3800 2023.4100 1261.9800 2467.4000 ;
      LAYER met3 ;
        RECT 1275.9200 2457.2400 1277.5200 2457.7200 ;
        RECT 1275.9200 2451.8000 1277.5200 2452.2800 ;
        RECT 1275.9200 2446.3600 1277.5200 2446.8400 ;
        RECT 1275.9200 2440.9200 1277.5200 2441.4000 ;
        RECT 1275.9200 2435.4800 1277.5200 2435.9600 ;
        RECT 1275.9200 2430.0400 1277.5200 2430.5200 ;
        RECT 1275.9200 2424.6000 1277.5200 2425.0800 ;
        RECT 1275.9200 2419.1600 1277.5200 2419.6400 ;
        RECT 1275.9200 2408.2800 1277.5200 2408.7600 ;
        RECT 1275.9200 2402.8400 1277.5200 2403.3200 ;
        RECT 1275.9200 2397.4000 1277.5200 2397.8800 ;
        RECT 1275.9200 2391.9600 1277.5200 2392.4400 ;
        RECT 1275.9200 2386.5200 1277.5200 2387.0000 ;
        RECT 1275.9200 2381.0800 1277.5200 2381.5600 ;
        RECT 1275.9200 2375.6400 1277.5200 2376.1200 ;
        RECT 1275.9200 2370.2000 1277.5200 2370.6800 ;
        RECT 1275.9200 2364.7600 1277.5200 2365.2400 ;
        RECT 1275.9200 2359.3200 1277.5200 2359.8000 ;
        RECT 1275.9200 2413.7200 1277.5200 2414.2000 ;
        RECT 1275.9200 2353.8800 1277.5200 2354.3600 ;
        RECT 1275.9200 2348.4400 1277.5200 2348.9200 ;
        RECT 1275.9200 2343.0000 1277.5200 2343.4800 ;
        RECT 1275.9200 2337.5600 1277.5200 2338.0400 ;
        RECT 1275.9200 2332.1200 1277.5200 2332.6000 ;
        RECT 1275.9200 2326.6800 1277.5200 2327.1600 ;
        RECT 1275.9200 2321.2400 1277.5200 2321.7200 ;
        RECT 1275.9200 2315.8000 1277.5200 2316.2800 ;
        RECT 1275.9200 2310.3600 1277.5200 2310.8400 ;
        RECT 1275.9200 2304.9200 1277.5200 2305.4000 ;
        RECT 1275.9200 2299.4800 1277.5200 2299.9600 ;
        RECT 1275.9200 2294.0400 1277.5200 2294.5200 ;
        RECT 1275.9200 2288.6000 1277.5200 2289.0800 ;
        RECT 1275.9200 2283.1600 1277.5200 2283.6400 ;
        RECT 1275.9200 2277.7200 1277.5200 2278.2000 ;
        RECT 1275.9200 2272.2800 1277.5200 2272.7600 ;
        RECT 1275.9200 2266.8400 1277.5200 2267.3200 ;
        RECT 1275.9200 2261.4000 1277.5200 2261.8800 ;
        RECT 1275.9200 2255.9600 1277.5200 2256.4400 ;
        RECT 1275.9200 2250.5200 1277.5200 2251.0000 ;
        RECT 1073.2200 2457.2400 1074.8200 2457.7200 ;
        RECT 1073.2200 2451.8000 1074.8200 2452.2800 ;
        RECT 1073.2200 2446.3600 1074.8200 2446.8400 ;
        RECT 1073.2200 2440.9200 1074.8200 2441.4000 ;
        RECT 1073.2200 2435.4800 1074.8200 2435.9600 ;
        RECT 1073.2200 2430.0400 1074.8200 2430.5200 ;
        RECT 1073.2200 2424.6000 1074.8200 2425.0800 ;
        RECT 1073.2200 2419.1600 1074.8200 2419.6400 ;
        RECT 1073.2200 2408.2800 1074.8200 2408.7600 ;
        RECT 1073.2200 2402.8400 1074.8200 2403.3200 ;
        RECT 1073.2200 2397.4000 1074.8200 2397.8800 ;
        RECT 1073.2200 2391.9600 1074.8200 2392.4400 ;
        RECT 1073.2200 2386.5200 1074.8200 2387.0000 ;
        RECT 1073.2200 2381.0800 1074.8200 2381.5600 ;
        RECT 1073.2200 2375.6400 1074.8200 2376.1200 ;
        RECT 1073.2200 2370.2000 1074.8200 2370.6800 ;
        RECT 1073.2200 2364.7600 1074.8200 2365.2400 ;
        RECT 1073.2200 2359.3200 1074.8200 2359.8000 ;
        RECT 1073.2200 2413.7200 1074.8200 2414.2000 ;
        RECT 1073.2200 2353.8800 1074.8200 2354.3600 ;
        RECT 1073.2200 2348.4400 1074.8200 2348.9200 ;
        RECT 1073.2200 2343.0000 1074.8200 2343.4800 ;
        RECT 1073.2200 2337.5600 1074.8200 2338.0400 ;
        RECT 1073.2200 2332.1200 1074.8200 2332.6000 ;
        RECT 1073.2200 2326.6800 1074.8200 2327.1600 ;
        RECT 1073.2200 2321.2400 1074.8200 2321.7200 ;
        RECT 1073.2200 2315.8000 1074.8200 2316.2800 ;
        RECT 1073.2200 2310.3600 1074.8200 2310.8400 ;
        RECT 1073.2200 2304.9200 1074.8200 2305.4000 ;
        RECT 1073.2200 2299.4800 1074.8200 2299.9600 ;
        RECT 1073.2200 2294.0400 1074.8200 2294.5200 ;
        RECT 1073.2200 2288.6000 1074.8200 2289.0800 ;
        RECT 1073.2200 2283.1600 1074.8200 2283.6400 ;
        RECT 1073.2200 2277.7200 1074.8200 2278.2000 ;
        RECT 1073.2200 2272.2800 1074.8200 2272.7600 ;
        RECT 1073.2200 2266.8400 1074.8200 2267.3200 ;
        RECT 1073.2200 2261.4000 1074.8200 2261.8800 ;
        RECT 1073.2200 2255.9600 1074.8200 2256.4400 ;
        RECT 1073.2200 2250.5200 1074.8200 2251.0000 ;
        RECT 1275.9200 2239.6400 1277.5200 2240.1200 ;
        RECT 1275.9200 2234.2000 1277.5200 2234.6800 ;
        RECT 1275.9200 2228.7600 1277.5200 2229.2400 ;
        RECT 1275.9200 2223.3200 1277.5200 2223.8000 ;
        RECT 1275.9200 2217.8800 1277.5200 2218.3600 ;
        RECT 1275.9200 2212.4400 1277.5200 2212.9200 ;
        RECT 1275.9200 2207.0000 1277.5200 2207.4800 ;
        RECT 1275.9200 2201.5600 1277.5200 2202.0400 ;
        RECT 1275.9200 2196.1200 1277.5200 2196.6000 ;
        RECT 1275.9200 2190.6800 1277.5200 2191.1600 ;
        RECT 1275.9200 2185.2400 1277.5200 2185.7200 ;
        RECT 1275.9200 2179.8000 1277.5200 2180.2800 ;
        RECT 1275.9200 2174.3600 1277.5200 2174.8400 ;
        RECT 1275.9200 2168.9200 1277.5200 2169.4000 ;
        RECT 1275.9200 2163.4800 1277.5200 2163.9600 ;
        RECT 1275.9200 2158.0400 1277.5200 2158.5200 ;
        RECT 1275.9200 2152.6000 1277.5200 2153.0800 ;
        RECT 1275.9200 2147.1600 1277.5200 2147.6400 ;
        RECT 1275.9200 2141.7200 1277.5200 2142.2000 ;
        RECT 1275.9200 2136.2800 1277.5200 2136.7600 ;
        RECT 1275.9200 2130.8400 1277.5200 2131.3200 ;
        RECT 1275.9200 2125.4000 1277.5200 2125.8800 ;
        RECT 1275.9200 2119.9600 1277.5200 2120.4400 ;
        RECT 1275.9200 2114.5200 1277.5200 2115.0000 ;
        RECT 1275.9200 2109.0800 1277.5200 2109.5600 ;
        RECT 1275.9200 2103.6400 1277.5200 2104.1200 ;
        RECT 1275.9200 2098.2000 1277.5200 2098.6800 ;
        RECT 1275.9200 2092.7600 1277.5200 2093.2400 ;
        RECT 1275.9200 2087.3200 1277.5200 2087.8000 ;
        RECT 1275.9200 2081.8800 1277.5200 2082.3600 ;
        RECT 1275.9200 2071.0000 1277.5200 2071.4800 ;
        RECT 1275.9200 2065.5600 1277.5200 2066.0400 ;
        RECT 1275.9200 2060.1200 1277.5200 2060.6000 ;
        RECT 1275.9200 2054.6800 1277.5200 2055.1600 ;
        RECT 1275.9200 2049.2400 1277.5200 2049.7200 ;
        RECT 1275.9200 2043.8000 1277.5200 2044.2800 ;
        RECT 1275.9200 2038.3600 1277.5200 2038.8400 ;
        RECT 1275.9200 2032.9200 1277.5200 2033.4000 ;
        RECT 1275.9200 2076.4400 1277.5200 2076.9200 ;
        RECT 1073.2200 2239.6400 1074.8200 2240.1200 ;
        RECT 1073.2200 2234.2000 1074.8200 2234.6800 ;
        RECT 1073.2200 2228.7600 1074.8200 2229.2400 ;
        RECT 1073.2200 2223.3200 1074.8200 2223.8000 ;
        RECT 1073.2200 2217.8800 1074.8200 2218.3600 ;
        RECT 1073.2200 2212.4400 1074.8200 2212.9200 ;
        RECT 1073.2200 2207.0000 1074.8200 2207.4800 ;
        RECT 1073.2200 2201.5600 1074.8200 2202.0400 ;
        RECT 1073.2200 2196.1200 1074.8200 2196.6000 ;
        RECT 1073.2200 2190.6800 1074.8200 2191.1600 ;
        RECT 1073.2200 2185.2400 1074.8200 2185.7200 ;
        RECT 1073.2200 2179.8000 1074.8200 2180.2800 ;
        RECT 1073.2200 2174.3600 1074.8200 2174.8400 ;
        RECT 1073.2200 2168.9200 1074.8200 2169.4000 ;
        RECT 1073.2200 2163.4800 1074.8200 2163.9600 ;
        RECT 1073.2200 2158.0400 1074.8200 2158.5200 ;
        RECT 1073.2200 2152.6000 1074.8200 2153.0800 ;
        RECT 1073.2200 2147.1600 1074.8200 2147.6400 ;
        RECT 1073.2200 2141.7200 1074.8200 2142.2000 ;
        RECT 1073.2200 2136.2800 1074.8200 2136.7600 ;
        RECT 1073.2200 2130.8400 1074.8200 2131.3200 ;
        RECT 1073.2200 2125.4000 1074.8200 2125.8800 ;
        RECT 1073.2200 2119.9600 1074.8200 2120.4400 ;
        RECT 1073.2200 2114.5200 1074.8200 2115.0000 ;
        RECT 1073.2200 2109.0800 1074.8200 2109.5600 ;
        RECT 1073.2200 2103.6400 1074.8200 2104.1200 ;
        RECT 1073.2200 2098.2000 1074.8200 2098.6800 ;
        RECT 1073.2200 2092.7600 1074.8200 2093.2400 ;
        RECT 1073.2200 2087.3200 1074.8200 2087.8000 ;
        RECT 1073.2200 2081.8800 1074.8200 2082.3600 ;
        RECT 1073.2200 2071.0000 1074.8200 2071.4800 ;
        RECT 1073.2200 2065.5600 1074.8200 2066.0400 ;
        RECT 1073.2200 2060.1200 1074.8200 2060.6000 ;
        RECT 1073.2200 2054.6800 1074.8200 2055.1600 ;
        RECT 1073.2200 2049.2400 1074.8200 2049.7200 ;
        RECT 1073.2200 2043.8000 1074.8200 2044.2800 ;
        RECT 1073.2200 2038.3600 1074.8200 2038.8400 ;
        RECT 1073.2200 2032.9200 1074.8200 2033.4000 ;
        RECT 1073.2200 2076.4400 1074.8200 2076.9200 ;
        RECT 1275.9200 2245.0800 1277.5200 2245.5600 ;
        RECT 1073.2200 2245.0800 1074.8200 2245.5600 ;
        RECT 1070.2600 2465.8000 1280.4800 2467.4000 ;
        RECT 1070.2600 2023.4100 1280.4800 2025.0100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 2020.5800 1074.8200 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 2468.8000 1074.8200 2470.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 2020.5800 1277.5200 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 2468.8000 1277.5200 2470.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 2023.4100 1071.8600 2025.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 2023.4100 1280.4800 2025.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 2465.8000 1071.8600 2467.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 2465.8000 1280.4800 2467.4000 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1073.2200 1561.3000 1074.8200 2011.1200 ;
        RECT 1275.9200 1561.3000 1277.5200 2011.1200 ;
        RECT 1080.3800 1564.1300 1081.9800 2008.1200 ;
        RECT 1125.3800 1564.1300 1126.9800 2008.1200 ;
        RECT 1170.3800 1564.1300 1171.9800 2008.1200 ;
        RECT 1215.3800 1564.1300 1216.9800 2008.1200 ;
        RECT 1260.3800 1564.1300 1261.9800 2008.1200 ;
      LAYER met3 ;
        RECT 1275.9200 1997.9600 1277.5200 1998.4400 ;
        RECT 1275.9200 1992.5200 1277.5200 1993.0000 ;
        RECT 1275.9200 1987.0800 1277.5200 1987.5600 ;
        RECT 1275.9200 1981.6400 1277.5200 1982.1200 ;
        RECT 1275.9200 1976.2000 1277.5200 1976.6800 ;
        RECT 1275.9200 1970.7600 1277.5200 1971.2400 ;
        RECT 1275.9200 1965.3200 1277.5200 1965.8000 ;
        RECT 1275.9200 1959.8800 1277.5200 1960.3600 ;
        RECT 1275.9200 1949.0000 1277.5200 1949.4800 ;
        RECT 1275.9200 1943.5600 1277.5200 1944.0400 ;
        RECT 1275.9200 1938.1200 1277.5200 1938.6000 ;
        RECT 1275.9200 1932.6800 1277.5200 1933.1600 ;
        RECT 1275.9200 1927.2400 1277.5200 1927.7200 ;
        RECT 1275.9200 1921.8000 1277.5200 1922.2800 ;
        RECT 1275.9200 1916.3600 1277.5200 1916.8400 ;
        RECT 1275.9200 1910.9200 1277.5200 1911.4000 ;
        RECT 1275.9200 1905.4800 1277.5200 1905.9600 ;
        RECT 1275.9200 1900.0400 1277.5200 1900.5200 ;
        RECT 1275.9200 1954.4400 1277.5200 1954.9200 ;
        RECT 1275.9200 1894.6000 1277.5200 1895.0800 ;
        RECT 1275.9200 1889.1600 1277.5200 1889.6400 ;
        RECT 1275.9200 1883.7200 1277.5200 1884.2000 ;
        RECT 1275.9200 1878.2800 1277.5200 1878.7600 ;
        RECT 1275.9200 1872.8400 1277.5200 1873.3200 ;
        RECT 1275.9200 1867.4000 1277.5200 1867.8800 ;
        RECT 1275.9200 1861.9600 1277.5200 1862.4400 ;
        RECT 1275.9200 1856.5200 1277.5200 1857.0000 ;
        RECT 1275.9200 1851.0800 1277.5200 1851.5600 ;
        RECT 1275.9200 1845.6400 1277.5200 1846.1200 ;
        RECT 1275.9200 1840.2000 1277.5200 1840.6800 ;
        RECT 1275.9200 1834.7600 1277.5200 1835.2400 ;
        RECT 1275.9200 1829.3200 1277.5200 1829.8000 ;
        RECT 1275.9200 1823.8800 1277.5200 1824.3600 ;
        RECT 1275.9200 1818.4400 1277.5200 1818.9200 ;
        RECT 1275.9200 1813.0000 1277.5200 1813.4800 ;
        RECT 1275.9200 1807.5600 1277.5200 1808.0400 ;
        RECT 1275.9200 1802.1200 1277.5200 1802.6000 ;
        RECT 1275.9200 1796.6800 1277.5200 1797.1600 ;
        RECT 1275.9200 1791.2400 1277.5200 1791.7200 ;
        RECT 1073.2200 1997.9600 1074.8200 1998.4400 ;
        RECT 1073.2200 1992.5200 1074.8200 1993.0000 ;
        RECT 1073.2200 1987.0800 1074.8200 1987.5600 ;
        RECT 1073.2200 1981.6400 1074.8200 1982.1200 ;
        RECT 1073.2200 1976.2000 1074.8200 1976.6800 ;
        RECT 1073.2200 1970.7600 1074.8200 1971.2400 ;
        RECT 1073.2200 1965.3200 1074.8200 1965.8000 ;
        RECT 1073.2200 1959.8800 1074.8200 1960.3600 ;
        RECT 1073.2200 1949.0000 1074.8200 1949.4800 ;
        RECT 1073.2200 1943.5600 1074.8200 1944.0400 ;
        RECT 1073.2200 1938.1200 1074.8200 1938.6000 ;
        RECT 1073.2200 1932.6800 1074.8200 1933.1600 ;
        RECT 1073.2200 1927.2400 1074.8200 1927.7200 ;
        RECT 1073.2200 1921.8000 1074.8200 1922.2800 ;
        RECT 1073.2200 1916.3600 1074.8200 1916.8400 ;
        RECT 1073.2200 1910.9200 1074.8200 1911.4000 ;
        RECT 1073.2200 1905.4800 1074.8200 1905.9600 ;
        RECT 1073.2200 1900.0400 1074.8200 1900.5200 ;
        RECT 1073.2200 1954.4400 1074.8200 1954.9200 ;
        RECT 1073.2200 1894.6000 1074.8200 1895.0800 ;
        RECT 1073.2200 1889.1600 1074.8200 1889.6400 ;
        RECT 1073.2200 1883.7200 1074.8200 1884.2000 ;
        RECT 1073.2200 1878.2800 1074.8200 1878.7600 ;
        RECT 1073.2200 1872.8400 1074.8200 1873.3200 ;
        RECT 1073.2200 1867.4000 1074.8200 1867.8800 ;
        RECT 1073.2200 1861.9600 1074.8200 1862.4400 ;
        RECT 1073.2200 1856.5200 1074.8200 1857.0000 ;
        RECT 1073.2200 1851.0800 1074.8200 1851.5600 ;
        RECT 1073.2200 1845.6400 1074.8200 1846.1200 ;
        RECT 1073.2200 1840.2000 1074.8200 1840.6800 ;
        RECT 1073.2200 1834.7600 1074.8200 1835.2400 ;
        RECT 1073.2200 1829.3200 1074.8200 1829.8000 ;
        RECT 1073.2200 1823.8800 1074.8200 1824.3600 ;
        RECT 1073.2200 1818.4400 1074.8200 1818.9200 ;
        RECT 1073.2200 1813.0000 1074.8200 1813.4800 ;
        RECT 1073.2200 1807.5600 1074.8200 1808.0400 ;
        RECT 1073.2200 1802.1200 1074.8200 1802.6000 ;
        RECT 1073.2200 1796.6800 1074.8200 1797.1600 ;
        RECT 1073.2200 1791.2400 1074.8200 1791.7200 ;
        RECT 1275.9200 1780.3600 1277.5200 1780.8400 ;
        RECT 1275.9200 1774.9200 1277.5200 1775.4000 ;
        RECT 1275.9200 1769.4800 1277.5200 1769.9600 ;
        RECT 1275.9200 1764.0400 1277.5200 1764.5200 ;
        RECT 1275.9200 1758.6000 1277.5200 1759.0800 ;
        RECT 1275.9200 1753.1600 1277.5200 1753.6400 ;
        RECT 1275.9200 1747.7200 1277.5200 1748.2000 ;
        RECT 1275.9200 1742.2800 1277.5200 1742.7600 ;
        RECT 1275.9200 1736.8400 1277.5200 1737.3200 ;
        RECT 1275.9200 1731.4000 1277.5200 1731.8800 ;
        RECT 1275.9200 1725.9600 1277.5200 1726.4400 ;
        RECT 1275.9200 1720.5200 1277.5200 1721.0000 ;
        RECT 1275.9200 1715.0800 1277.5200 1715.5600 ;
        RECT 1275.9200 1709.6400 1277.5200 1710.1200 ;
        RECT 1275.9200 1704.2000 1277.5200 1704.6800 ;
        RECT 1275.9200 1698.7600 1277.5200 1699.2400 ;
        RECT 1275.9200 1693.3200 1277.5200 1693.8000 ;
        RECT 1275.9200 1687.8800 1277.5200 1688.3600 ;
        RECT 1275.9200 1682.4400 1277.5200 1682.9200 ;
        RECT 1275.9200 1677.0000 1277.5200 1677.4800 ;
        RECT 1275.9200 1671.5600 1277.5200 1672.0400 ;
        RECT 1275.9200 1666.1200 1277.5200 1666.6000 ;
        RECT 1275.9200 1660.6800 1277.5200 1661.1600 ;
        RECT 1275.9200 1655.2400 1277.5200 1655.7200 ;
        RECT 1275.9200 1649.8000 1277.5200 1650.2800 ;
        RECT 1275.9200 1644.3600 1277.5200 1644.8400 ;
        RECT 1275.9200 1638.9200 1277.5200 1639.4000 ;
        RECT 1275.9200 1633.4800 1277.5200 1633.9600 ;
        RECT 1275.9200 1628.0400 1277.5200 1628.5200 ;
        RECT 1275.9200 1622.6000 1277.5200 1623.0800 ;
        RECT 1275.9200 1611.7200 1277.5200 1612.2000 ;
        RECT 1275.9200 1606.2800 1277.5200 1606.7600 ;
        RECT 1275.9200 1600.8400 1277.5200 1601.3200 ;
        RECT 1275.9200 1595.4000 1277.5200 1595.8800 ;
        RECT 1275.9200 1589.9600 1277.5200 1590.4400 ;
        RECT 1275.9200 1584.5200 1277.5200 1585.0000 ;
        RECT 1275.9200 1579.0800 1277.5200 1579.5600 ;
        RECT 1275.9200 1573.6400 1277.5200 1574.1200 ;
        RECT 1275.9200 1617.1600 1277.5200 1617.6400 ;
        RECT 1073.2200 1780.3600 1074.8200 1780.8400 ;
        RECT 1073.2200 1774.9200 1074.8200 1775.4000 ;
        RECT 1073.2200 1769.4800 1074.8200 1769.9600 ;
        RECT 1073.2200 1764.0400 1074.8200 1764.5200 ;
        RECT 1073.2200 1758.6000 1074.8200 1759.0800 ;
        RECT 1073.2200 1753.1600 1074.8200 1753.6400 ;
        RECT 1073.2200 1747.7200 1074.8200 1748.2000 ;
        RECT 1073.2200 1742.2800 1074.8200 1742.7600 ;
        RECT 1073.2200 1736.8400 1074.8200 1737.3200 ;
        RECT 1073.2200 1731.4000 1074.8200 1731.8800 ;
        RECT 1073.2200 1725.9600 1074.8200 1726.4400 ;
        RECT 1073.2200 1720.5200 1074.8200 1721.0000 ;
        RECT 1073.2200 1715.0800 1074.8200 1715.5600 ;
        RECT 1073.2200 1709.6400 1074.8200 1710.1200 ;
        RECT 1073.2200 1704.2000 1074.8200 1704.6800 ;
        RECT 1073.2200 1698.7600 1074.8200 1699.2400 ;
        RECT 1073.2200 1693.3200 1074.8200 1693.8000 ;
        RECT 1073.2200 1687.8800 1074.8200 1688.3600 ;
        RECT 1073.2200 1682.4400 1074.8200 1682.9200 ;
        RECT 1073.2200 1677.0000 1074.8200 1677.4800 ;
        RECT 1073.2200 1671.5600 1074.8200 1672.0400 ;
        RECT 1073.2200 1666.1200 1074.8200 1666.6000 ;
        RECT 1073.2200 1660.6800 1074.8200 1661.1600 ;
        RECT 1073.2200 1655.2400 1074.8200 1655.7200 ;
        RECT 1073.2200 1649.8000 1074.8200 1650.2800 ;
        RECT 1073.2200 1644.3600 1074.8200 1644.8400 ;
        RECT 1073.2200 1638.9200 1074.8200 1639.4000 ;
        RECT 1073.2200 1633.4800 1074.8200 1633.9600 ;
        RECT 1073.2200 1628.0400 1074.8200 1628.5200 ;
        RECT 1073.2200 1622.6000 1074.8200 1623.0800 ;
        RECT 1073.2200 1611.7200 1074.8200 1612.2000 ;
        RECT 1073.2200 1606.2800 1074.8200 1606.7600 ;
        RECT 1073.2200 1600.8400 1074.8200 1601.3200 ;
        RECT 1073.2200 1595.4000 1074.8200 1595.8800 ;
        RECT 1073.2200 1589.9600 1074.8200 1590.4400 ;
        RECT 1073.2200 1584.5200 1074.8200 1585.0000 ;
        RECT 1073.2200 1579.0800 1074.8200 1579.5600 ;
        RECT 1073.2200 1573.6400 1074.8200 1574.1200 ;
        RECT 1073.2200 1617.1600 1074.8200 1617.6400 ;
        RECT 1275.9200 1785.8000 1277.5200 1786.2800 ;
        RECT 1073.2200 1785.8000 1074.8200 1786.2800 ;
        RECT 1070.2600 2006.5200 1280.4800 2008.1200 ;
        RECT 1070.2600 1564.1300 1280.4800 1565.7300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 1561.3000 1074.8200 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 2009.5200 1074.8200 2011.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 1561.3000 1277.5200 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 2009.5200 1277.5200 2011.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1564.1300 1071.8600 1565.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1564.1300 1280.4800 1565.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 2006.5200 1071.8600 2008.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 2006.5200 1280.4800 2008.1200 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1073.2200 1102.0200 1074.8200 1551.8400 ;
        RECT 1275.9200 1102.0200 1277.5200 1551.8400 ;
        RECT 1080.3800 1104.8500 1081.9800 1548.8400 ;
        RECT 1125.3800 1104.8500 1126.9800 1548.8400 ;
        RECT 1170.3800 1104.8500 1171.9800 1548.8400 ;
        RECT 1215.3800 1104.8500 1216.9800 1548.8400 ;
        RECT 1260.3800 1104.8500 1261.9800 1548.8400 ;
      LAYER met3 ;
        RECT 1275.9200 1538.6800 1277.5200 1539.1600 ;
        RECT 1275.9200 1533.2400 1277.5200 1533.7200 ;
        RECT 1275.9200 1527.8000 1277.5200 1528.2800 ;
        RECT 1275.9200 1522.3600 1277.5200 1522.8400 ;
        RECT 1275.9200 1516.9200 1277.5200 1517.4000 ;
        RECT 1275.9200 1511.4800 1277.5200 1511.9600 ;
        RECT 1275.9200 1506.0400 1277.5200 1506.5200 ;
        RECT 1275.9200 1500.6000 1277.5200 1501.0800 ;
        RECT 1275.9200 1489.7200 1277.5200 1490.2000 ;
        RECT 1275.9200 1484.2800 1277.5200 1484.7600 ;
        RECT 1275.9200 1478.8400 1277.5200 1479.3200 ;
        RECT 1275.9200 1473.4000 1277.5200 1473.8800 ;
        RECT 1275.9200 1467.9600 1277.5200 1468.4400 ;
        RECT 1275.9200 1462.5200 1277.5200 1463.0000 ;
        RECT 1275.9200 1457.0800 1277.5200 1457.5600 ;
        RECT 1275.9200 1451.6400 1277.5200 1452.1200 ;
        RECT 1275.9200 1446.2000 1277.5200 1446.6800 ;
        RECT 1275.9200 1440.7600 1277.5200 1441.2400 ;
        RECT 1275.9200 1495.1600 1277.5200 1495.6400 ;
        RECT 1275.9200 1435.3200 1277.5200 1435.8000 ;
        RECT 1275.9200 1429.8800 1277.5200 1430.3600 ;
        RECT 1275.9200 1424.4400 1277.5200 1424.9200 ;
        RECT 1275.9200 1419.0000 1277.5200 1419.4800 ;
        RECT 1275.9200 1413.5600 1277.5200 1414.0400 ;
        RECT 1275.9200 1408.1200 1277.5200 1408.6000 ;
        RECT 1275.9200 1402.6800 1277.5200 1403.1600 ;
        RECT 1275.9200 1397.2400 1277.5200 1397.7200 ;
        RECT 1275.9200 1391.8000 1277.5200 1392.2800 ;
        RECT 1275.9200 1386.3600 1277.5200 1386.8400 ;
        RECT 1275.9200 1380.9200 1277.5200 1381.4000 ;
        RECT 1275.9200 1375.4800 1277.5200 1375.9600 ;
        RECT 1275.9200 1370.0400 1277.5200 1370.5200 ;
        RECT 1275.9200 1364.6000 1277.5200 1365.0800 ;
        RECT 1275.9200 1359.1600 1277.5200 1359.6400 ;
        RECT 1275.9200 1353.7200 1277.5200 1354.2000 ;
        RECT 1275.9200 1348.2800 1277.5200 1348.7600 ;
        RECT 1275.9200 1342.8400 1277.5200 1343.3200 ;
        RECT 1275.9200 1337.4000 1277.5200 1337.8800 ;
        RECT 1275.9200 1331.9600 1277.5200 1332.4400 ;
        RECT 1073.2200 1538.6800 1074.8200 1539.1600 ;
        RECT 1073.2200 1533.2400 1074.8200 1533.7200 ;
        RECT 1073.2200 1527.8000 1074.8200 1528.2800 ;
        RECT 1073.2200 1522.3600 1074.8200 1522.8400 ;
        RECT 1073.2200 1516.9200 1074.8200 1517.4000 ;
        RECT 1073.2200 1511.4800 1074.8200 1511.9600 ;
        RECT 1073.2200 1506.0400 1074.8200 1506.5200 ;
        RECT 1073.2200 1500.6000 1074.8200 1501.0800 ;
        RECT 1073.2200 1489.7200 1074.8200 1490.2000 ;
        RECT 1073.2200 1484.2800 1074.8200 1484.7600 ;
        RECT 1073.2200 1478.8400 1074.8200 1479.3200 ;
        RECT 1073.2200 1473.4000 1074.8200 1473.8800 ;
        RECT 1073.2200 1467.9600 1074.8200 1468.4400 ;
        RECT 1073.2200 1462.5200 1074.8200 1463.0000 ;
        RECT 1073.2200 1457.0800 1074.8200 1457.5600 ;
        RECT 1073.2200 1451.6400 1074.8200 1452.1200 ;
        RECT 1073.2200 1446.2000 1074.8200 1446.6800 ;
        RECT 1073.2200 1440.7600 1074.8200 1441.2400 ;
        RECT 1073.2200 1495.1600 1074.8200 1495.6400 ;
        RECT 1073.2200 1435.3200 1074.8200 1435.8000 ;
        RECT 1073.2200 1429.8800 1074.8200 1430.3600 ;
        RECT 1073.2200 1424.4400 1074.8200 1424.9200 ;
        RECT 1073.2200 1419.0000 1074.8200 1419.4800 ;
        RECT 1073.2200 1413.5600 1074.8200 1414.0400 ;
        RECT 1073.2200 1408.1200 1074.8200 1408.6000 ;
        RECT 1073.2200 1402.6800 1074.8200 1403.1600 ;
        RECT 1073.2200 1397.2400 1074.8200 1397.7200 ;
        RECT 1073.2200 1391.8000 1074.8200 1392.2800 ;
        RECT 1073.2200 1386.3600 1074.8200 1386.8400 ;
        RECT 1073.2200 1380.9200 1074.8200 1381.4000 ;
        RECT 1073.2200 1375.4800 1074.8200 1375.9600 ;
        RECT 1073.2200 1370.0400 1074.8200 1370.5200 ;
        RECT 1073.2200 1364.6000 1074.8200 1365.0800 ;
        RECT 1073.2200 1359.1600 1074.8200 1359.6400 ;
        RECT 1073.2200 1353.7200 1074.8200 1354.2000 ;
        RECT 1073.2200 1348.2800 1074.8200 1348.7600 ;
        RECT 1073.2200 1342.8400 1074.8200 1343.3200 ;
        RECT 1073.2200 1337.4000 1074.8200 1337.8800 ;
        RECT 1073.2200 1331.9600 1074.8200 1332.4400 ;
        RECT 1275.9200 1321.0800 1277.5200 1321.5600 ;
        RECT 1275.9200 1315.6400 1277.5200 1316.1200 ;
        RECT 1275.9200 1310.2000 1277.5200 1310.6800 ;
        RECT 1275.9200 1304.7600 1277.5200 1305.2400 ;
        RECT 1275.9200 1299.3200 1277.5200 1299.8000 ;
        RECT 1275.9200 1293.8800 1277.5200 1294.3600 ;
        RECT 1275.9200 1288.4400 1277.5200 1288.9200 ;
        RECT 1275.9200 1283.0000 1277.5200 1283.4800 ;
        RECT 1275.9200 1277.5600 1277.5200 1278.0400 ;
        RECT 1275.9200 1272.1200 1277.5200 1272.6000 ;
        RECT 1275.9200 1266.6800 1277.5200 1267.1600 ;
        RECT 1275.9200 1261.2400 1277.5200 1261.7200 ;
        RECT 1275.9200 1255.8000 1277.5200 1256.2800 ;
        RECT 1275.9200 1250.3600 1277.5200 1250.8400 ;
        RECT 1275.9200 1244.9200 1277.5200 1245.4000 ;
        RECT 1275.9200 1239.4800 1277.5200 1239.9600 ;
        RECT 1275.9200 1234.0400 1277.5200 1234.5200 ;
        RECT 1275.9200 1228.6000 1277.5200 1229.0800 ;
        RECT 1275.9200 1223.1600 1277.5200 1223.6400 ;
        RECT 1275.9200 1217.7200 1277.5200 1218.2000 ;
        RECT 1275.9200 1212.2800 1277.5200 1212.7600 ;
        RECT 1275.9200 1206.8400 1277.5200 1207.3200 ;
        RECT 1275.9200 1201.4000 1277.5200 1201.8800 ;
        RECT 1275.9200 1195.9600 1277.5200 1196.4400 ;
        RECT 1275.9200 1190.5200 1277.5200 1191.0000 ;
        RECT 1275.9200 1185.0800 1277.5200 1185.5600 ;
        RECT 1275.9200 1179.6400 1277.5200 1180.1200 ;
        RECT 1275.9200 1174.2000 1277.5200 1174.6800 ;
        RECT 1275.9200 1168.7600 1277.5200 1169.2400 ;
        RECT 1275.9200 1163.3200 1277.5200 1163.8000 ;
        RECT 1275.9200 1152.4400 1277.5200 1152.9200 ;
        RECT 1275.9200 1147.0000 1277.5200 1147.4800 ;
        RECT 1275.9200 1141.5600 1277.5200 1142.0400 ;
        RECT 1275.9200 1136.1200 1277.5200 1136.6000 ;
        RECT 1275.9200 1130.6800 1277.5200 1131.1600 ;
        RECT 1275.9200 1125.2400 1277.5200 1125.7200 ;
        RECT 1275.9200 1119.8000 1277.5200 1120.2800 ;
        RECT 1275.9200 1114.3600 1277.5200 1114.8400 ;
        RECT 1275.9200 1157.8800 1277.5200 1158.3600 ;
        RECT 1073.2200 1321.0800 1074.8200 1321.5600 ;
        RECT 1073.2200 1315.6400 1074.8200 1316.1200 ;
        RECT 1073.2200 1310.2000 1074.8200 1310.6800 ;
        RECT 1073.2200 1304.7600 1074.8200 1305.2400 ;
        RECT 1073.2200 1299.3200 1074.8200 1299.8000 ;
        RECT 1073.2200 1293.8800 1074.8200 1294.3600 ;
        RECT 1073.2200 1288.4400 1074.8200 1288.9200 ;
        RECT 1073.2200 1283.0000 1074.8200 1283.4800 ;
        RECT 1073.2200 1277.5600 1074.8200 1278.0400 ;
        RECT 1073.2200 1272.1200 1074.8200 1272.6000 ;
        RECT 1073.2200 1266.6800 1074.8200 1267.1600 ;
        RECT 1073.2200 1261.2400 1074.8200 1261.7200 ;
        RECT 1073.2200 1255.8000 1074.8200 1256.2800 ;
        RECT 1073.2200 1250.3600 1074.8200 1250.8400 ;
        RECT 1073.2200 1244.9200 1074.8200 1245.4000 ;
        RECT 1073.2200 1239.4800 1074.8200 1239.9600 ;
        RECT 1073.2200 1234.0400 1074.8200 1234.5200 ;
        RECT 1073.2200 1228.6000 1074.8200 1229.0800 ;
        RECT 1073.2200 1223.1600 1074.8200 1223.6400 ;
        RECT 1073.2200 1217.7200 1074.8200 1218.2000 ;
        RECT 1073.2200 1212.2800 1074.8200 1212.7600 ;
        RECT 1073.2200 1206.8400 1074.8200 1207.3200 ;
        RECT 1073.2200 1201.4000 1074.8200 1201.8800 ;
        RECT 1073.2200 1195.9600 1074.8200 1196.4400 ;
        RECT 1073.2200 1190.5200 1074.8200 1191.0000 ;
        RECT 1073.2200 1185.0800 1074.8200 1185.5600 ;
        RECT 1073.2200 1179.6400 1074.8200 1180.1200 ;
        RECT 1073.2200 1174.2000 1074.8200 1174.6800 ;
        RECT 1073.2200 1168.7600 1074.8200 1169.2400 ;
        RECT 1073.2200 1163.3200 1074.8200 1163.8000 ;
        RECT 1073.2200 1152.4400 1074.8200 1152.9200 ;
        RECT 1073.2200 1147.0000 1074.8200 1147.4800 ;
        RECT 1073.2200 1141.5600 1074.8200 1142.0400 ;
        RECT 1073.2200 1136.1200 1074.8200 1136.6000 ;
        RECT 1073.2200 1130.6800 1074.8200 1131.1600 ;
        RECT 1073.2200 1125.2400 1074.8200 1125.7200 ;
        RECT 1073.2200 1119.8000 1074.8200 1120.2800 ;
        RECT 1073.2200 1114.3600 1074.8200 1114.8400 ;
        RECT 1073.2200 1157.8800 1074.8200 1158.3600 ;
        RECT 1275.9200 1326.5200 1277.5200 1327.0000 ;
        RECT 1073.2200 1326.5200 1074.8200 1327.0000 ;
        RECT 1070.2600 1547.2400 1280.4800 1548.8400 ;
        RECT 1070.2600 1104.8500 1280.4800 1106.4500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 1102.0200 1074.8200 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 1550.2400 1074.8200 1551.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 1102.0200 1277.5200 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 1550.2400 1277.5200 1551.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1104.8500 1071.8600 1106.4500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1104.8500 1280.4800 1106.4500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1547.2400 1071.8600 1548.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1547.2400 1280.4800 1548.8400 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1073.2200 642.7400 1074.8200 1092.5600 ;
        RECT 1275.9200 642.7400 1277.5200 1092.5600 ;
        RECT 1080.3800 645.5700 1081.9800 1089.5600 ;
        RECT 1125.3800 645.5700 1126.9800 1089.5600 ;
        RECT 1170.3800 645.5700 1171.9800 1089.5600 ;
        RECT 1215.3800 645.5700 1216.9800 1089.5600 ;
        RECT 1260.3800 645.5700 1261.9800 1089.5600 ;
      LAYER met3 ;
        RECT 1275.9200 1079.4000 1277.5200 1079.8800 ;
        RECT 1275.9200 1073.9600 1277.5200 1074.4400 ;
        RECT 1275.9200 1068.5200 1277.5200 1069.0000 ;
        RECT 1275.9200 1063.0800 1277.5200 1063.5600 ;
        RECT 1275.9200 1057.6400 1277.5200 1058.1200 ;
        RECT 1275.9200 1052.2000 1277.5200 1052.6800 ;
        RECT 1275.9200 1046.7600 1277.5200 1047.2400 ;
        RECT 1275.9200 1041.3200 1277.5200 1041.8000 ;
        RECT 1275.9200 1030.4400 1277.5200 1030.9200 ;
        RECT 1275.9200 1025.0000 1277.5200 1025.4800 ;
        RECT 1275.9200 1019.5600 1277.5200 1020.0400 ;
        RECT 1275.9200 1014.1200 1277.5200 1014.6000 ;
        RECT 1275.9200 1008.6800 1277.5200 1009.1600 ;
        RECT 1275.9200 1003.2400 1277.5200 1003.7200 ;
        RECT 1275.9200 997.8000 1277.5200 998.2800 ;
        RECT 1275.9200 992.3600 1277.5200 992.8400 ;
        RECT 1275.9200 986.9200 1277.5200 987.4000 ;
        RECT 1275.9200 981.4800 1277.5200 981.9600 ;
        RECT 1275.9200 1035.8800 1277.5200 1036.3600 ;
        RECT 1275.9200 976.0400 1277.5200 976.5200 ;
        RECT 1275.9200 970.6000 1277.5200 971.0800 ;
        RECT 1275.9200 965.1600 1277.5200 965.6400 ;
        RECT 1275.9200 959.7200 1277.5200 960.2000 ;
        RECT 1275.9200 954.2800 1277.5200 954.7600 ;
        RECT 1275.9200 948.8400 1277.5200 949.3200 ;
        RECT 1275.9200 943.4000 1277.5200 943.8800 ;
        RECT 1275.9200 937.9600 1277.5200 938.4400 ;
        RECT 1275.9200 932.5200 1277.5200 933.0000 ;
        RECT 1275.9200 927.0800 1277.5200 927.5600 ;
        RECT 1275.9200 921.6400 1277.5200 922.1200 ;
        RECT 1275.9200 916.2000 1277.5200 916.6800 ;
        RECT 1275.9200 910.7600 1277.5200 911.2400 ;
        RECT 1275.9200 905.3200 1277.5200 905.8000 ;
        RECT 1275.9200 899.8800 1277.5200 900.3600 ;
        RECT 1275.9200 894.4400 1277.5200 894.9200 ;
        RECT 1275.9200 889.0000 1277.5200 889.4800 ;
        RECT 1275.9200 883.5600 1277.5200 884.0400 ;
        RECT 1275.9200 878.1200 1277.5200 878.6000 ;
        RECT 1275.9200 872.6800 1277.5200 873.1600 ;
        RECT 1073.2200 1079.4000 1074.8200 1079.8800 ;
        RECT 1073.2200 1073.9600 1074.8200 1074.4400 ;
        RECT 1073.2200 1068.5200 1074.8200 1069.0000 ;
        RECT 1073.2200 1063.0800 1074.8200 1063.5600 ;
        RECT 1073.2200 1057.6400 1074.8200 1058.1200 ;
        RECT 1073.2200 1052.2000 1074.8200 1052.6800 ;
        RECT 1073.2200 1046.7600 1074.8200 1047.2400 ;
        RECT 1073.2200 1041.3200 1074.8200 1041.8000 ;
        RECT 1073.2200 1030.4400 1074.8200 1030.9200 ;
        RECT 1073.2200 1025.0000 1074.8200 1025.4800 ;
        RECT 1073.2200 1019.5600 1074.8200 1020.0400 ;
        RECT 1073.2200 1014.1200 1074.8200 1014.6000 ;
        RECT 1073.2200 1008.6800 1074.8200 1009.1600 ;
        RECT 1073.2200 1003.2400 1074.8200 1003.7200 ;
        RECT 1073.2200 997.8000 1074.8200 998.2800 ;
        RECT 1073.2200 992.3600 1074.8200 992.8400 ;
        RECT 1073.2200 986.9200 1074.8200 987.4000 ;
        RECT 1073.2200 981.4800 1074.8200 981.9600 ;
        RECT 1073.2200 1035.8800 1074.8200 1036.3600 ;
        RECT 1073.2200 976.0400 1074.8200 976.5200 ;
        RECT 1073.2200 970.6000 1074.8200 971.0800 ;
        RECT 1073.2200 965.1600 1074.8200 965.6400 ;
        RECT 1073.2200 959.7200 1074.8200 960.2000 ;
        RECT 1073.2200 954.2800 1074.8200 954.7600 ;
        RECT 1073.2200 948.8400 1074.8200 949.3200 ;
        RECT 1073.2200 943.4000 1074.8200 943.8800 ;
        RECT 1073.2200 937.9600 1074.8200 938.4400 ;
        RECT 1073.2200 932.5200 1074.8200 933.0000 ;
        RECT 1073.2200 927.0800 1074.8200 927.5600 ;
        RECT 1073.2200 921.6400 1074.8200 922.1200 ;
        RECT 1073.2200 916.2000 1074.8200 916.6800 ;
        RECT 1073.2200 910.7600 1074.8200 911.2400 ;
        RECT 1073.2200 905.3200 1074.8200 905.8000 ;
        RECT 1073.2200 899.8800 1074.8200 900.3600 ;
        RECT 1073.2200 894.4400 1074.8200 894.9200 ;
        RECT 1073.2200 889.0000 1074.8200 889.4800 ;
        RECT 1073.2200 883.5600 1074.8200 884.0400 ;
        RECT 1073.2200 878.1200 1074.8200 878.6000 ;
        RECT 1073.2200 872.6800 1074.8200 873.1600 ;
        RECT 1275.9200 861.8000 1277.5200 862.2800 ;
        RECT 1275.9200 856.3600 1277.5200 856.8400 ;
        RECT 1275.9200 850.9200 1277.5200 851.4000 ;
        RECT 1275.9200 845.4800 1277.5200 845.9600 ;
        RECT 1275.9200 840.0400 1277.5200 840.5200 ;
        RECT 1275.9200 834.6000 1277.5200 835.0800 ;
        RECT 1275.9200 829.1600 1277.5200 829.6400 ;
        RECT 1275.9200 823.7200 1277.5200 824.2000 ;
        RECT 1275.9200 818.2800 1277.5200 818.7600 ;
        RECT 1275.9200 812.8400 1277.5200 813.3200 ;
        RECT 1275.9200 807.4000 1277.5200 807.8800 ;
        RECT 1275.9200 801.9600 1277.5200 802.4400 ;
        RECT 1275.9200 796.5200 1277.5200 797.0000 ;
        RECT 1275.9200 791.0800 1277.5200 791.5600 ;
        RECT 1275.9200 785.6400 1277.5200 786.1200 ;
        RECT 1275.9200 780.2000 1277.5200 780.6800 ;
        RECT 1275.9200 774.7600 1277.5200 775.2400 ;
        RECT 1275.9200 769.3200 1277.5200 769.8000 ;
        RECT 1275.9200 763.8800 1277.5200 764.3600 ;
        RECT 1275.9200 758.4400 1277.5200 758.9200 ;
        RECT 1275.9200 753.0000 1277.5200 753.4800 ;
        RECT 1275.9200 747.5600 1277.5200 748.0400 ;
        RECT 1275.9200 742.1200 1277.5200 742.6000 ;
        RECT 1275.9200 736.6800 1277.5200 737.1600 ;
        RECT 1275.9200 731.2400 1277.5200 731.7200 ;
        RECT 1275.9200 725.8000 1277.5200 726.2800 ;
        RECT 1275.9200 720.3600 1277.5200 720.8400 ;
        RECT 1275.9200 714.9200 1277.5200 715.4000 ;
        RECT 1275.9200 709.4800 1277.5200 709.9600 ;
        RECT 1275.9200 704.0400 1277.5200 704.5200 ;
        RECT 1275.9200 693.1600 1277.5200 693.6400 ;
        RECT 1275.9200 687.7200 1277.5200 688.2000 ;
        RECT 1275.9200 682.2800 1277.5200 682.7600 ;
        RECT 1275.9200 676.8400 1277.5200 677.3200 ;
        RECT 1275.9200 671.4000 1277.5200 671.8800 ;
        RECT 1275.9200 665.9600 1277.5200 666.4400 ;
        RECT 1275.9200 660.5200 1277.5200 661.0000 ;
        RECT 1275.9200 655.0800 1277.5200 655.5600 ;
        RECT 1275.9200 698.6000 1277.5200 699.0800 ;
        RECT 1073.2200 861.8000 1074.8200 862.2800 ;
        RECT 1073.2200 856.3600 1074.8200 856.8400 ;
        RECT 1073.2200 850.9200 1074.8200 851.4000 ;
        RECT 1073.2200 845.4800 1074.8200 845.9600 ;
        RECT 1073.2200 840.0400 1074.8200 840.5200 ;
        RECT 1073.2200 834.6000 1074.8200 835.0800 ;
        RECT 1073.2200 829.1600 1074.8200 829.6400 ;
        RECT 1073.2200 823.7200 1074.8200 824.2000 ;
        RECT 1073.2200 818.2800 1074.8200 818.7600 ;
        RECT 1073.2200 812.8400 1074.8200 813.3200 ;
        RECT 1073.2200 807.4000 1074.8200 807.8800 ;
        RECT 1073.2200 801.9600 1074.8200 802.4400 ;
        RECT 1073.2200 796.5200 1074.8200 797.0000 ;
        RECT 1073.2200 791.0800 1074.8200 791.5600 ;
        RECT 1073.2200 785.6400 1074.8200 786.1200 ;
        RECT 1073.2200 780.2000 1074.8200 780.6800 ;
        RECT 1073.2200 774.7600 1074.8200 775.2400 ;
        RECT 1073.2200 769.3200 1074.8200 769.8000 ;
        RECT 1073.2200 763.8800 1074.8200 764.3600 ;
        RECT 1073.2200 758.4400 1074.8200 758.9200 ;
        RECT 1073.2200 753.0000 1074.8200 753.4800 ;
        RECT 1073.2200 747.5600 1074.8200 748.0400 ;
        RECT 1073.2200 742.1200 1074.8200 742.6000 ;
        RECT 1073.2200 736.6800 1074.8200 737.1600 ;
        RECT 1073.2200 731.2400 1074.8200 731.7200 ;
        RECT 1073.2200 725.8000 1074.8200 726.2800 ;
        RECT 1073.2200 720.3600 1074.8200 720.8400 ;
        RECT 1073.2200 714.9200 1074.8200 715.4000 ;
        RECT 1073.2200 709.4800 1074.8200 709.9600 ;
        RECT 1073.2200 704.0400 1074.8200 704.5200 ;
        RECT 1073.2200 693.1600 1074.8200 693.6400 ;
        RECT 1073.2200 687.7200 1074.8200 688.2000 ;
        RECT 1073.2200 682.2800 1074.8200 682.7600 ;
        RECT 1073.2200 676.8400 1074.8200 677.3200 ;
        RECT 1073.2200 671.4000 1074.8200 671.8800 ;
        RECT 1073.2200 665.9600 1074.8200 666.4400 ;
        RECT 1073.2200 660.5200 1074.8200 661.0000 ;
        RECT 1073.2200 655.0800 1074.8200 655.5600 ;
        RECT 1073.2200 698.6000 1074.8200 699.0800 ;
        RECT 1275.9200 867.2400 1277.5200 867.7200 ;
        RECT 1073.2200 867.2400 1074.8200 867.7200 ;
        RECT 1070.2600 1087.9600 1280.4800 1089.5600 ;
        RECT 1070.2600 645.5700 1280.4800 647.1700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 642.7400 1074.8200 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 1090.9600 1074.8200 1092.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 642.7400 1277.5200 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 1090.9600 1277.5200 1092.5600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 645.5700 1071.8600 647.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 645.5700 1280.4800 647.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1087.9600 1071.8600 1089.5600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1087.9600 1280.4800 1089.5600 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1073.2200 183.4600 1074.8200 633.2800 ;
        RECT 1275.9200 183.4600 1277.5200 633.2800 ;
        RECT 1080.3800 186.2900 1081.9800 630.2800 ;
        RECT 1125.3800 186.2900 1126.9800 630.2800 ;
        RECT 1170.3800 186.2900 1171.9800 630.2800 ;
        RECT 1215.3800 186.2900 1216.9800 630.2800 ;
        RECT 1260.3800 186.2900 1261.9800 630.2800 ;
      LAYER met3 ;
        RECT 1275.9200 620.1200 1277.5200 620.6000 ;
        RECT 1275.9200 614.6800 1277.5200 615.1600 ;
        RECT 1275.9200 609.2400 1277.5200 609.7200 ;
        RECT 1275.9200 603.8000 1277.5200 604.2800 ;
        RECT 1275.9200 598.3600 1277.5200 598.8400 ;
        RECT 1275.9200 592.9200 1277.5200 593.4000 ;
        RECT 1275.9200 587.4800 1277.5200 587.9600 ;
        RECT 1275.9200 582.0400 1277.5200 582.5200 ;
        RECT 1275.9200 571.1600 1277.5200 571.6400 ;
        RECT 1275.9200 565.7200 1277.5200 566.2000 ;
        RECT 1275.9200 560.2800 1277.5200 560.7600 ;
        RECT 1275.9200 554.8400 1277.5200 555.3200 ;
        RECT 1275.9200 549.4000 1277.5200 549.8800 ;
        RECT 1275.9200 543.9600 1277.5200 544.4400 ;
        RECT 1275.9200 538.5200 1277.5200 539.0000 ;
        RECT 1275.9200 533.0800 1277.5200 533.5600 ;
        RECT 1275.9200 527.6400 1277.5200 528.1200 ;
        RECT 1275.9200 522.2000 1277.5200 522.6800 ;
        RECT 1275.9200 576.6000 1277.5200 577.0800 ;
        RECT 1275.9200 516.7600 1277.5200 517.2400 ;
        RECT 1275.9200 511.3200 1277.5200 511.8000 ;
        RECT 1275.9200 505.8800 1277.5200 506.3600 ;
        RECT 1275.9200 500.4400 1277.5200 500.9200 ;
        RECT 1275.9200 495.0000 1277.5200 495.4800 ;
        RECT 1275.9200 489.5600 1277.5200 490.0400 ;
        RECT 1275.9200 484.1200 1277.5200 484.6000 ;
        RECT 1275.9200 478.6800 1277.5200 479.1600 ;
        RECT 1275.9200 473.2400 1277.5200 473.7200 ;
        RECT 1275.9200 467.8000 1277.5200 468.2800 ;
        RECT 1275.9200 462.3600 1277.5200 462.8400 ;
        RECT 1275.9200 456.9200 1277.5200 457.4000 ;
        RECT 1275.9200 451.4800 1277.5200 451.9600 ;
        RECT 1275.9200 446.0400 1277.5200 446.5200 ;
        RECT 1275.9200 440.6000 1277.5200 441.0800 ;
        RECT 1275.9200 435.1600 1277.5200 435.6400 ;
        RECT 1275.9200 429.7200 1277.5200 430.2000 ;
        RECT 1275.9200 424.2800 1277.5200 424.7600 ;
        RECT 1275.9200 418.8400 1277.5200 419.3200 ;
        RECT 1275.9200 413.4000 1277.5200 413.8800 ;
        RECT 1073.2200 620.1200 1074.8200 620.6000 ;
        RECT 1073.2200 614.6800 1074.8200 615.1600 ;
        RECT 1073.2200 609.2400 1074.8200 609.7200 ;
        RECT 1073.2200 603.8000 1074.8200 604.2800 ;
        RECT 1073.2200 598.3600 1074.8200 598.8400 ;
        RECT 1073.2200 592.9200 1074.8200 593.4000 ;
        RECT 1073.2200 587.4800 1074.8200 587.9600 ;
        RECT 1073.2200 582.0400 1074.8200 582.5200 ;
        RECT 1073.2200 571.1600 1074.8200 571.6400 ;
        RECT 1073.2200 565.7200 1074.8200 566.2000 ;
        RECT 1073.2200 560.2800 1074.8200 560.7600 ;
        RECT 1073.2200 554.8400 1074.8200 555.3200 ;
        RECT 1073.2200 549.4000 1074.8200 549.8800 ;
        RECT 1073.2200 543.9600 1074.8200 544.4400 ;
        RECT 1073.2200 538.5200 1074.8200 539.0000 ;
        RECT 1073.2200 533.0800 1074.8200 533.5600 ;
        RECT 1073.2200 527.6400 1074.8200 528.1200 ;
        RECT 1073.2200 522.2000 1074.8200 522.6800 ;
        RECT 1073.2200 576.6000 1074.8200 577.0800 ;
        RECT 1073.2200 516.7600 1074.8200 517.2400 ;
        RECT 1073.2200 511.3200 1074.8200 511.8000 ;
        RECT 1073.2200 505.8800 1074.8200 506.3600 ;
        RECT 1073.2200 500.4400 1074.8200 500.9200 ;
        RECT 1073.2200 495.0000 1074.8200 495.4800 ;
        RECT 1073.2200 489.5600 1074.8200 490.0400 ;
        RECT 1073.2200 484.1200 1074.8200 484.6000 ;
        RECT 1073.2200 478.6800 1074.8200 479.1600 ;
        RECT 1073.2200 473.2400 1074.8200 473.7200 ;
        RECT 1073.2200 467.8000 1074.8200 468.2800 ;
        RECT 1073.2200 462.3600 1074.8200 462.8400 ;
        RECT 1073.2200 456.9200 1074.8200 457.4000 ;
        RECT 1073.2200 451.4800 1074.8200 451.9600 ;
        RECT 1073.2200 446.0400 1074.8200 446.5200 ;
        RECT 1073.2200 440.6000 1074.8200 441.0800 ;
        RECT 1073.2200 435.1600 1074.8200 435.6400 ;
        RECT 1073.2200 429.7200 1074.8200 430.2000 ;
        RECT 1073.2200 424.2800 1074.8200 424.7600 ;
        RECT 1073.2200 418.8400 1074.8200 419.3200 ;
        RECT 1073.2200 413.4000 1074.8200 413.8800 ;
        RECT 1275.9200 402.5200 1277.5200 403.0000 ;
        RECT 1275.9200 397.0800 1277.5200 397.5600 ;
        RECT 1275.9200 391.6400 1277.5200 392.1200 ;
        RECT 1275.9200 386.2000 1277.5200 386.6800 ;
        RECT 1275.9200 380.7600 1277.5200 381.2400 ;
        RECT 1275.9200 375.3200 1277.5200 375.8000 ;
        RECT 1275.9200 369.8800 1277.5200 370.3600 ;
        RECT 1275.9200 364.4400 1277.5200 364.9200 ;
        RECT 1275.9200 359.0000 1277.5200 359.4800 ;
        RECT 1275.9200 353.5600 1277.5200 354.0400 ;
        RECT 1275.9200 348.1200 1277.5200 348.6000 ;
        RECT 1275.9200 342.6800 1277.5200 343.1600 ;
        RECT 1275.9200 337.2400 1277.5200 337.7200 ;
        RECT 1275.9200 331.8000 1277.5200 332.2800 ;
        RECT 1275.9200 326.3600 1277.5200 326.8400 ;
        RECT 1275.9200 320.9200 1277.5200 321.4000 ;
        RECT 1275.9200 315.4800 1277.5200 315.9600 ;
        RECT 1275.9200 310.0400 1277.5200 310.5200 ;
        RECT 1275.9200 304.6000 1277.5200 305.0800 ;
        RECT 1275.9200 299.1600 1277.5200 299.6400 ;
        RECT 1275.9200 293.7200 1277.5200 294.2000 ;
        RECT 1275.9200 288.2800 1277.5200 288.7600 ;
        RECT 1275.9200 282.8400 1277.5200 283.3200 ;
        RECT 1275.9200 277.4000 1277.5200 277.8800 ;
        RECT 1275.9200 271.9600 1277.5200 272.4400 ;
        RECT 1275.9200 266.5200 1277.5200 267.0000 ;
        RECT 1275.9200 261.0800 1277.5200 261.5600 ;
        RECT 1275.9200 255.6400 1277.5200 256.1200 ;
        RECT 1275.9200 250.2000 1277.5200 250.6800 ;
        RECT 1275.9200 244.7600 1277.5200 245.2400 ;
        RECT 1275.9200 233.8800 1277.5200 234.3600 ;
        RECT 1275.9200 228.4400 1277.5200 228.9200 ;
        RECT 1275.9200 223.0000 1277.5200 223.4800 ;
        RECT 1275.9200 217.5600 1277.5200 218.0400 ;
        RECT 1275.9200 212.1200 1277.5200 212.6000 ;
        RECT 1275.9200 206.6800 1277.5200 207.1600 ;
        RECT 1275.9200 201.2400 1277.5200 201.7200 ;
        RECT 1275.9200 195.8000 1277.5200 196.2800 ;
        RECT 1275.9200 239.3200 1277.5200 239.8000 ;
        RECT 1073.2200 402.5200 1074.8200 403.0000 ;
        RECT 1073.2200 397.0800 1074.8200 397.5600 ;
        RECT 1073.2200 391.6400 1074.8200 392.1200 ;
        RECT 1073.2200 386.2000 1074.8200 386.6800 ;
        RECT 1073.2200 380.7600 1074.8200 381.2400 ;
        RECT 1073.2200 375.3200 1074.8200 375.8000 ;
        RECT 1073.2200 369.8800 1074.8200 370.3600 ;
        RECT 1073.2200 364.4400 1074.8200 364.9200 ;
        RECT 1073.2200 359.0000 1074.8200 359.4800 ;
        RECT 1073.2200 353.5600 1074.8200 354.0400 ;
        RECT 1073.2200 348.1200 1074.8200 348.6000 ;
        RECT 1073.2200 342.6800 1074.8200 343.1600 ;
        RECT 1073.2200 337.2400 1074.8200 337.7200 ;
        RECT 1073.2200 331.8000 1074.8200 332.2800 ;
        RECT 1073.2200 326.3600 1074.8200 326.8400 ;
        RECT 1073.2200 320.9200 1074.8200 321.4000 ;
        RECT 1073.2200 315.4800 1074.8200 315.9600 ;
        RECT 1073.2200 310.0400 1074.8200 310.5200 ;
        RECT 1073.2200 304.6000 1074.8200 305.0800 ;
        RECT 1073.2200 299.1600 1074.8200 299.6400 ;
        RECT 1073.2200 293.7200 1074.8200 294.2000 ;
        RECT 1073.2200 288.2800 1074.8200 288.7600 ;
        RECT 1073.2200 282.8400 1074.8200 283.3200 ;
        RECT 1073.2200 277.4000 1074.8200 277.8800 ;
        RECT 1073.2200 271.9600 1074.8200 272.4400 ;
        RECT 1073.2200 266.5200 1074.8200 267.0000 ;
        RECT 1073.2200 261.0800 1074.8200 261.5600 ;
        RECT 1073.2200 255.6400 1074.8200 256.1200 ;
        RECT 1073.2200 250.2000 1074.8200 250.6800 ;
        RECT 1073.2200 244.7600 1074.8200 245.2400 ;
        RECT 1073.2200 233.8800 1074.8200 234.3600 ;
        RECT 1073.2200 228.4400 1074.8200 228.9200 ;
        RECT 1073.2200 223.0000 1074.8200 223.4800 ;
        RECT 1073.2200 217.5600 1074.8200 218.0400 ;
        RECT 1073.2200 212.1200 1074.8200 212.6000 ;
        RECT 1073.2200 206.6800 1074.8200 207.1600 ;
        RECT 1073.2200 201.2400 1074.8200 201.7200 ;
        RECT 1073.2200 195.8000 1074.8200 196.2800 ;
        RECT 1073.2200 239.3200 1074.8200 239.8000 ;
        RECT 1275.9200 407.9600 1277.5200 408.4400 ;
        RECT 1073.2200 407.9600 1074.8200 408.4400 ;
        RECT 1070.2600 628.6800 1280.4800 630.2800 ;
        RECT 1070.2600 186.2900 1280.4800 187.8900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 183.4600 1074.8200 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.2200 631.6800 1074.8200 633.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 183.4600 1277.5200 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.9200 631.6800 1277.5200 633.2800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 186.2900 1071.8600 187.8900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 186.2900 1280.4800 187.8900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 628.6800 1071.8600 630.2800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 628.6800 1280.4800 630.2800 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1293.4000 2479.6000 1295.0000 2509.8600 ;
        RECT 1495.9000 2479.6000 1497.5000 2509.8600 ;
      LAYER met3 ;
        RECT 1495.9000 2500.1000 1497.5000 2500.5800 ;
        RECT 1293.4000 2500.1000 1295.0000 2500.5800 ;
        RECT 1495.9000 2489.2200 1497.5000 2489.7000 ;
        RECT 1293.4000 2489.2200 1295.0000 2489.7000 ;
        RECT 1495.9000 2494.6600 1497.5000 2495.1400 ;
        RECT 1293.4000 2494.6600 1295.0000 2495.1400 ;
        RECT 1290.3400 2505.5000 1500.5600 2507.1000 ;
        RECT 1290.3400 2481.1700 1500.5600 2482.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.4000 2479.6000 1295.0000 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.4000 2508.2600 1295.0000 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1495.9000 2479.6000 1497.5000 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1495.9000 2508.2600 1497.5000 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2481.1700 1291.9400 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2481.1700 1500.5600 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2505.5000 1291.9400 2507.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2505.5000 1500.5600 2507.1000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 186.0300 1482.0600 399.3300 ;
        RECT 1435.4600 186.0300 1437.0600 399.3300 ;
        RECT 1390.4600 186.0300 1392.0600 399.3300 ;
        RECT 1345.4600 186.0300 1347.0600 399.3300 ;
        RECT 1300.4600 186.0300 1302.0600 399.3300 ;
        RECT 1496.0000 183.2000 1497.6000 402.8400 ;
        RECT 1293.3000 183.2000 1294.9000 402.8400 ;
      LAYER met3 ;
        RECT 1480.4600 391.3800 1482.0600 391.8600 ;
        RECT 1496.0000 391.3800 1497.6000 391.8600 ;
        RECT 1496.0000 380.5000 1497.6000 380.9800 ;
        RECT 1496.0000 385.9400 1497.6000 386.4200 ;
        RECT 1480.4600 380.5000 1482.0600 380.9800 ;
        RECT 1480.4600 385.9400 1482.0600 386.4200 ;
        RECT 1496.0000 364.1800 1497.6000 364.6600 ;
        RECT 1496.0000 369.6200 1497.6000 370.1000 ;
        RECT 1480.4600 364.1800 1482.0600 364.6600 ;
        RECT 1480.4600 369.6200 1482.0600 370.1000 ;
        RECT 1496.0000 353.3000 1497.6000 353.7800 ;
        RECT 1496.0000 358.7400 1497.6000 359.2200 ;
        RECT 1480.4600 353.3000 1482.0600 353.7800 ;
        RECT 1480.4600 358.7400 1482.0600 359.2200 ;
        RECT 1480.4600 375.0600 1482.0600 375.5400 ;
        RECT 1496.0000 375.0600 1497.6000 375.5400 ;
        RECT 1435.4600 380.5000 1437.0600 380.9800 ;
        RECT 1435.4600 385.9400 1437.0600 386.4200 ;
        RECT 1435.4600 391.3800 1437.0600 391.8600 ;
        RECT 1435.4600 364.1800 1437.0600 364.6600 ;
        RECT 1435.4600 369.6200 1437.0600 370.1000 ;
        RECT 1435.4600 358.7400 1437.0600 359.2200 ;
        RECT 1435.4600 353.3000 1437.0600 353.7800 ;
        RECT 1435.4600 375.0600 1437.0600 375.5400 ;
        RECT 1496.0000 336.9800 1497.6000 337.4600 ;
        RECT 1496.0000 342.4200 1497.6000 342.9000 ;
        RECT 1480.4600 336.9800 1482.0600 337.4600 ;
        RECT 1480.4600 342.4200 1482.0600 342.9000 ;
        RECT 1496.0000 320.6600 1497.6000 321.1400 ;
        RECT 1496.0000 326.1000 1497.6000 326.5800 ;
        RECT 1496.0000 331.5400 1497.6000 332.0200 ;
        RECT 1480.4600 320.6600 1482.0600 321.1400 ;
        RECT 1480.4600 326.1000 1482.0600 326.5800 ;
        RECT 1480.4600 331.5400 1482.0600 332.0200 ;
        RECT 1496.0000 309.7800 1497.6000 310.2600 ;
        RECT 1496.0000 315.2200 1497.6000 315.7000 ;
        RECT 1480.4600 309.7800 1482.0600 310.2600 ;
        RECT 1480.4600 315.2200 1482.0600 315.7000 ;
        RECT 1496.0000 293.4600 1497.6000 293.9400 ;
        RECT 1496.0000 298.9000 1497.6000 299.3800 ;
        RECT 1496.0000 304.3400 1497.6000 304.8200 ;
        RECT 1480.4600 293.4600 1482.0600 293.9400 ;
        RECT 1480.4600 298.9000 1482.0600 299.3800 ;
        RECT 1480.4600 304.3400 1482.0600 304.8200 ;
        RECT 1435.4600 336.9800 1437.0600 337.4600 ;
        RECT 1435.4600 342.4200 1437.0600 342.9000 ;
        RECT 1435.4600 320.6600 1437.0600 321.1400 ;
        RECT 1435.4600 326.1000 1437.0600 326.5800 ;
        RECT 1435.4600 331.5400 1437.0600 332.0200 ;
        RECT 1435.4600 309.7800 1437.0600 310.2600 ;
        RECT 1435.4600 315.2200 1437.0600 315.7000 ;
        RECT 1435.4600 293.4600 1437.0600 293.9400 ;
        RECT 1435.4600 298.9000 1437.0600 299.3800 ;
        RECT 1435.4600 304.3400 1437.0600 304.8200 ;
        RECT 1435.4600 347.8600 1437.0600 348.3400 ;
        RECT 1480.4600 347.8600 1482.0600 348.3400 ;
        RECT 1496.0000 347.8600 1497.6000 348.3400 ;
        RECT 1390.4600 380.5000 1392.0600 380.9800 ;
        RECT 1390.4600 385.9400 1392.0600 386.4200 ;
        RECT 1390.4600 391.3800 1392.0600 391.8600 ;
        RECT 1345.4600 380.5000 1347.0600 380.9800 ;
        RECT 1345.4600 385.9400 1347.0600 386.4200 ;
        RECT 1345.4600 391.3800 1347.0600 391.8600 ;
        RECT 1390.4600 364.1800 1392.0600 364.6600 ;
        RECT 1390.4600 369.6200 1392.0600 370.1000 ;
        RECT 1390.4600 353.3000 1392.0600 353.7800 ;
        RECT 1390.4600 358.7400 1392.0600 359.2200 ;
        RECT 1345.4600 364.1800 1347.0600 364.6600 ;
        RECT 1345.4600 369.6200 1347.0600 370.1000 ;
        RECT 1345.4600 353.3000 1347.0600 353.7800 ;
        RECT 1345.4600 358.7400 1347.0600 359.2200 ;
        RECT 1345.4600 375.0600 1347.0600 375.5400 ;
        RECT 1390.4600 375.0600 1392.0600 375.5400 ;
        RECT 1293.3000 391.3800 1294.9000 391.8600 ;
        RECT 1300.4600 391.3800 1302.0600 391.8600 ;
        RECT 1300.4600 380.5000 1302.0600 380.9800 ;
        RECT 1300.4600 385.9400 1302.0600 386.4200 ;
        RECT 1293.3000 380.5000 1294.9000 380.9800 ;
        RECT 1293.3000 385.9400 1294.9000 386.4200 ;
        RECT 1300.4600 364.1800 1302.0600 364.6600 ;
        RECT 1300.4600 369.6200 1302.0600 370.1000 ;
        RECT 1293.3000 364.1800 1294.9000 364.6600 ;
        RECT 1293.3000 369.6200 1294.9000 370.1000 ;
        RECT 1300.4600 353.3000 1302.0600 353.7800 ;
        RECT 1300.4600 358.7400 1302.0600 359.2200 ;
        RECT 1293.3000 353.3000 1294.9000 353.7800 ;
        RECT 1293.3000 358.7400 1294.9000 359.2200 ;
        RECT 1293.3000 375.0600 1294.9000 375.5400 ;
        RECT 1300.4600 375.0600 1302.0600 375.5400 ;
        RECT 1390.4600 336.9800 1392.0600 337.4600 ;
        RECT 1390.4600 342.4200 1392.0600 342.9000 ;
        RECT 1390.4600 320.6600 1392.0600 321.1400 ;
        RECT 1390.4600 326.1000 1392.0600 326.5800 ;
        RECT 1390.4600 331.5400 1392.0600 332.0200 ;
        RECT 1345.4600 336.9800 1347.0600 337.4600 ;
        RECT 1345.4600 342.4200 1347.0600 342.9000 ;
        RECT 1345.4600 320.6600 1347.0600 321.1400 ;
        RECT 1345.4600 326.1000 1347.0600 326.5800 ;
        RECT 1345.4600 331.5400 1347.0600 332.0200 ;
        RECT 1390.4600 309.7800 1392.0600 310.2600 ;
        RECT 1390.4600 315.2200 1392.0600 315.7000 ;
        RECT 1390.4600 293.4600 1392.0600 293.9400 ;
        RECT 1390.4600 298.9000 1392.0600 299.3800 ;
        RECT 1390.4600 304.3400 1392.0600 304.8200 ;
        RECT 1345.4600 309.7800 1347.0600 310.2600 ;
        RECT 1345.4600 315.2200 1347.0600 315.7000 ;
        RECT 1345.4600 293.4600 1347.0600 293.9400 ;
        RECT 1345.4600 298.9000 1347.0600 299.3800 ;
        RECT 1345.4600 304.3400 1347.0600 304.8200 ;
        RECT 1300.4600 336.9800 1302.0600 337.4600 ;
        RECT 1300.4600 342.4200 1302.0600 342.9000 ;
        RECT 1293.3000 336.9800 1294.9000 337.4600 ;
        RECT 1293.3000 342.4200 1294.9000 342.9000 ;
        RECT 1300.4600 320.6600 1302.0600 321.1400 ;
        RECT 1300.4600 326.1000 1302.0600 326.5800 ;
        RECT 1300.4600 331.5400 1302.0600 332.0200 ;
        RECT 1293.3000 320.6600 1294.9000 321.1400 ;
        RECT 1293.3000 326.1000 1294.9000 326.5800 ;
        RECT 1293.3000 331.5400 1294.9000 332.0200 ;
        RECT 1300.4600 309.7800 1302.0600 310.2600 ;
        RECT 1300.4600 315.2200 1302.0600 315.7000 ;
        RECT 1293.3000 309.7800 1294.9000 310.2600 ;
        RECT 1293.3000 315.2200 1294.9000 315.7000 ;
        RECT 1300.4600 293.4600 1302.0600 293.9400 ;
        RECT 1300.4600 298.9000 1302.0600 299.3800 ;
        RECT 1300.4600 304.3400 1302.0600 304.8200 ;
        RECT 1293.3000 293.4600 1294.9000 293.9400 ;
        RECT 1293.3000 298.9000 1294.9000 299.3800 ;
        RECT 1293.3000 304.3400 1294.9000 304.8200 ;
        RECT 1293.3000 347.8600 1294.9000 348.3400 ;
        RECT 1300.4600 347.8600 1302.0600 348.3400 ;
        RECT 1345.4600 347.8600 1347.0600 348.3400 ;
        RECT 1390.4600 347.8600 1392.0600 348.3400 ;
        RECT 1496.0000 282.5800 1497.6000 283.0600 ;
        RECT 1496.0000 288.0200 1497.6000 288.5000 ;
        RECT 1480.4600 282.5800 1482.0600 283.0600 ;
        RECT 1480.4600 288.0200 1482.0600 288.5000 ;
        RECT 1496.0000 266.2600 1497.6000 266.7400 ;
        RECT 1496.0000 271.7000 1497.6000 272.1800 ;
        RECT 1496.0000 277.1400 1497.6000 277.6200 ;
        RECT 1480.4600 266.2600 1482.0600 266.7400 ;
        RECT 1480.4600 271.7000 1482.0600 272.1800 ;
        RECT 1480.4600 277.1400 1482.0600 277.6200 ;
        RECT 1496.0000 255.3800 1497.6000 255.8600 ;
        RECT 1496.0000 260.8200 1497.6000 261.3000 ;
        RECT 1480.4600 255.3800 1482.0600 255.8600 ;
        RECT 1480.4600 260.8200 1482.0600 261.3000 ;
        RECT 1496.0000 239.0600 1497.6000 239.5400 ;
        RECT 1496.0000 244.5000 1497.6000 244.9800 ;
        RECT 1496.0000 249.9400 1497.6000 250.4200 ;
        RECT 1480.4600 239.0600 1482.0600 239.5400 ;
        RECT 1480.4600 244.5000 1482.0600 244.9800 ;
        RECT 1480.4600 249.9400 1482.0600 250.4200 ;
        RECT 1435.4600 282.5800 1437.0600 283.0600 ;
        RECT 1435.4600 288.0200 1437.0600 288.5000 ;
        RECT 1435.4600 266.2600 1437.0600 266.7400 ;
        RECT 1435.4600 271.7000 1437.0600 272.1800 ;
        RECT 1435.4600 277.1400 1437.0600 277.6200 ;
        RECT 1435.4600 255.3800 1437.0600 255.8600 ;
        RECT 1435.4600 260.8200 1437.0600 261.3000 ;
        RECT 1435.4600 239.0600 1437.0600 239.5400 ;
        RECT 1435.4600 244.5000 1437.0600 244.9800 ;
        RECT 1435.4600 249.9400 1437.0600 250.4200 ;
        RECT 1496.0000 228.1800 1497.6000 228.6600 ;
        RECT 1496.0000 233.6200 1497.6000 234.1000 ;
        RECT 1480.4600 228.1800 1482.0600 228.6600 ;
        RECT 1480.4600 233.6200 1482.0600 234.1000 ;
        RECT 1496.0000 211.8600 1497.6000 212.3400 ;
        RECT 1496.0000 217.3000 1497.6000 217.7800 ;
        RECT 1496.0000 222.7400 1497.6000 223.2200 ;
        RECT 1480.4600 211.8600 1482.0600 212.3400 ;
        RECT 1480.4600 217.3000 1482.0600 217.7800 ;
        RECT 1480.4600 222.7400 1482.0600 223.2200 ;
        RECT 1496.0000 200.9800 1497.6000 201.4600 ;
        RECT 1496.0000 206.4200 1497.6000 206.9000 ;
        RECT 1480.4600 200.9800 1482.0600 201.4600 ;
        RECT 1480.4600 206.4200 1482.0600 206.9000 ;
        RECT 1480.4600 195.5400 1482.0600 196.0200 ;
        RECT 1496.0000 195.5400 1497.6000 196.0200 ;
        RECT 1435.4600 228.1800 1437.0600 228.6600 ;
        RECT 1435.4600 233.6200 1437.0600 234.1000 ;
        RECT 1435.4600 211.8600 1437.0600 212.3400 ;
        RECT 1435.4600 217.3000 1437.0600 217.7800 ;
        RECT 1435.4600 222.7400 1437.0600 223.2200 ;
        RECT 1435.4600 200.9800 1437.0600 201.4600 ;
        RECT 1435.4600 206.4200 1437.0600 206.9000 ;
        RECT 1435.4600 195.5400 1437.0600 196.0200 ;
        RECT 1390.4600 282.5800 1392.0600 283.0600 ;
        RECT 1390.4600 288.0200 1392.0600 288.5000 ;
        RECT 1390.4600 266.2600 1392.0600 266.7400 ;
        RECT 1390.4600 271.7000 1392.0600 272.1800 ;
        RECT 1390.4600 277.1400 1392.0600 277.6200 ;
        RECT 1345.4600 282.5800 1347.0600 283.0600 ;
        RECT 1345.4600 288.0200 1347.0600 288.5000 ;
        RECT 1345.4600 266.2600 1347.0600 266.7400 ;
        RECT 1345.4600 271.7000 1347.0600 272.1800 ;
        RECT 1345.4600 277.1400 1347.0600 277.6200 ;
        RECT 1390.4600 255.3800 1392.0600 255.8600 ;
        RECT 1390.4600 260.8200 1392.0600 261.3000 ;
        RECT 1390.4600 239.0600 1392.0600 239.5400 ;
        RECT 1390.4600 244.5000 1392.0600 244.9800 ;
        RECT 1390.4600 249.9400 1392.0600 250.4200 ;
        RECT 1345.4600 255.3800 1347.0600 255.8600 ;
        RECT 1345.4600 260.8200 1347.0600 261.3000 ;
        RECT 1345.4600 239.0600 1347.0600 239.5400 ;
        RECT 1345.4600 244.5000 1347.0600 244.9800 ;
        RECT 1345.4600 249.9400 1347.0600 250.4200 ;
        RECT 1300.4600 282.5800 1302.0600 283.0600 ;
        RECT 1300.4600 288.0200 1302.0600 288.5000 ;
        RECT 1293.3000 282.5800 1294.9000 283.0600 ;
        RECT 1293.3000 288.0200 1294.9000 288.5000 ;
        RECT 1300.4600 266.2600 1302.0600 266.7400 ;
        RECT 1300.4600 271.7000 1302.0600 272.1800 ;
        RECT 1300.4600 277.1400 1302.0600 277.6200 ;
        RECT 1293.3000 266.2600 1294.9000 266.7400 ;
        RECT 1293.3000 271.7000 1294.9000 272.1800 ;
        RECT 1293.3000 277.1400 1294.9000 277.6200 ;
        RECT 1300.4600 255.3800 1302.0600 255.8600 ;
        RECT 1300.4600 260.8200 1302.0600 261.3000 ;
        RECT 1293.3000 255.3800 1294.9000 255.8600 ;
        RECT 1293.3000 260.8200 1294.9000 261.3000 ;
        RECT 1300.4600 239.0600 1302.0600 239.5400 ;
        RECT 1300.4600 244.5000 1302.0600 244.9800 ;
        RECT 1300.4600 249.9400 1302.0600 250.4200 ;
        RECT 1293.3000 239.0600 1294.9000 239.5400 ;
        RECT 1293.3000 244.5000 1294.9000 244.9800 ;
        RECT 1293.3000 249.9400 1294.9000 250.4200 ;
        RECT 1390.4600 228.1800 1392.0600 228.6600 ;
        RECT 1390.4600 233.6200 1392.0600 234.1000 ;
        RECT 1390.4600 211.8600 1392.0600 212.3400 ;
        RECT 1390.4600 217.3000 1392.0600 217.7800 ;
        RECT 1390.4600 222.7400 1392.0600 223.2200 ;
        RECT 1345.4600 228.1800 1347.0600 228.6600 ;
        RECT 1345.4600 233.6200 1347.0600 234.1000 ;
        RECT 1345.4600 211.8600 1347.0600 212.3400 ;
        RECT 1345.4600 217.3000 1347.0600 217.7800 ;
        RECT 1345.4600 222.7400 1347.0600 223.2200 ;
        RECT 1390.4600 206.4200 1392.0600 206.9000 ;
        RECT 1390.4600 200.9800 1392.0600 201.4600 ;
        RECT 1390.4600 195.5400 1392.0600 196.0200 ;
        RECT 1345.4600 206.4200 1347.0600 206.9000 ;
        RECT 1345.4600 200.9800 1347.0600 201.4600 ;
        RECT 1345.4600 195.5400 1347.0600 196.0200 ;
        RECT 1300.4600 228.1800 1302.0600 228.6600 ;
        RECT 1300.4600 233.6200 1302.0600 234.1000 ;
        RECT 1293.3000 228.1800 1294.9000 228.6600 ;
        RECT 1293.3000 233.6200 1294.9000 234.1000 ;
        RECT 1300.4600 211.8600 1302.0600 212.3400 ;
        RECT 1300.4600 217.3000 1302.0600 217.7800 ;
        RECT 1300.4600 222.7400 1302.0600 223.2200 ;
        RECT 1293.3000 211.8600 1294.9000 212.3400 ;
        RECT 1293.3000 217.3000 1294.9000 217.7800 ;
        RECT 1293.3000 222.7400 1294.9000 223.2200 ;
        RECT 1300.4600 200.9800 1302.0600 201.4600 ;
        RECT 1300.4600 206.4200 1302.0600 206.9000 ;
        RECT 1293.3000 200.9800 1294.9000 201.4600 ;
        RECT 1293.3000 206.4200 1294.9000 206.9000 ;
        RECT 1293.3000 195.5400 1294.9000 196.0200 ;
        RECT 1300.4600 195.5400 1302.0600 196.0200 ;
        RECT 1290.3400 397.7300 1500.5600 399.3300 ;
        RECT 1290.3400 186.0300 1500.5600 187.6300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 183.2000 1294.9000 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 401.2400 1294.9000 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 183.2000 1497.6000 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 401.2400 1497.6000 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 186.0300 1291.9400 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 186.0300 1500.5600 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 397.7300 1291.9400 399.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 397.7300 1500.5600 399.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1293.4000 142.9400 1295.0000 173.2000 ;
        RECT 1495.9000 142.9400 1497.5000 173.2000 ;
      LAYER met3 ;
        RECT 1495.9000 163.4400 1497.5000 163.9200 ;
        RECT 1293.4000 163.4400 1295.0000 163.9200 ;
        RECT 1495.9000 152.5600 1497.5000 153.0400 ;
        RECT 1293.4000 152.5600 1295.0000 153.0400 ;
        RECT 1495.9000 158.0000 1497.5000 158.4800 ;
        RECT 1293.4000 158.0000 1295.0000 158.4800 ;
        RECT 1290.3400 168.8400 1500.5600 170.4400 ;
        RECT 1290.3400 144.5100 1500.5600 146.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.4000 142.9400 1295.0000 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.4000 171.6000 1295.0000 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1495.9000 142.9400 1497.5000 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1495.9000 171.6000 1497.5000 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 144.5100 1291.9400 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 144.5100 1500.5600 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 168.8400 1291.9400 170.4400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 168.8400 1500.5600 170.4400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 2252.7900 1482.0600 2466.0900 ;
        RECT 1435.4600 2252.7900 1437.0600 2466.0900 ;
        RECT 1390.4600 2252.7900 1392.0600 2466.0900 ;
        RECT 1345.4600 2252.7900 1347.0600 2466.0900 ;
        RECT 1300.4600 2252.7900 1302.0600 2466.0900 ;
        RECT 1496.0000 2249.9600 1497.6000 2469.6000 ;
        RECT 1293.3000 2249.9600 1294.9000 2469.6000 ;
      LAYER met3 ;
        RECT 1480.4600 2458.1400 1482.0600 2458.6200 ;
        RECT 1496.0000 2458.1400 1497.6000 2458.6200 ;
        RECT 1496.0000 2447.2600 1497.6000 2447.7400 ;
        RECT 1496.0000 2452.7000 1497.6000 2453.1800 ;
        RECT 1480.4600 2447.2600 1482.0600 2447.7400 ;
        RECT 1480.4600 2452.7000 1482.0600 2453.1800 ;
        RECT 1496.0000 2430.9400 1497.6000 2431.4200 ;
        RECT 1496.0000 2436.3800 1497.6000 2436.8600 ;
        RECT 1480.4600 2430.9400 1482.0600 2431.4200 ;
        RECT 1480.4600 2436.3800 1482.0600 2436.8600 ;
        RECT 1496.0000 2420.0600 1497.6000 2420.5400 ;
        RECT 1496.0000 2425.5000 1497.6000 2425.9800 ;
        RECT 1480.4600 2420.0600 1482.0600 2420.5400 ;
        RECT 1480.4600 2425.5000 1482.0600 2425.9800 ;
        RECT 1480.4600 2441.8200 1482.0600 2442.3000 ;
        RECT 1496.0000 2441.8200 1497.6000 2442.3000 ;
        RECT 1435.4600 2447.2600 1437.0600 2447.7400 ;
        RECT 1435.4600 2452.7000 1437.0600 2453.1800 ;
        RECT 1435.4600 2458.1400 1437.0600 2458.6200 ;
        RECT 1435.4600 2430.9400 1437.0600 2431.4200 ;
        RECT 1435.4600 2436.3800 1437.0600 2436.8600 ;
        RECT 1435.4600 2425.5000 1437.0600 2425.9800 ;
        RECT 1435.4600 2420.0600 1437.0600 2420.5400 ;
        RECT 1435.4600 2441.8200 1437.0600 2442.3000 ;
        RECT 1496.0000 2403.7400 1497.6000 2404.2200 ;
        RECT 1496.0000 2409.1800 1497.6000 2409.6600 ;
        RECT 1480.4600 2403.7400 1482.0600 2404.2200 ;
        RECT 1480.4600 2409.1800 1482.0600 2409.6600 ;
        RECT 1496.0000 2387.4200 1497.6000 2387.9000 ;
        RECT 1496.0000 2392.8600 1497.6000 2393.3400 ;
        RECT 1496.0000 2398.3000 1497.6000 2398.7800 ;
        RECT 1480.4600 2387.4200 1482.0600 2387.9000 ;
        RECT 1480.4600 2392.8600 1482.0600 2393.3400 ;
        RECT 1480.4600 2398.3000 1482.0600 2398.7800 ;
        RECT 1496.0000 2376.5400 1497.6000 2377.0200 ;
        RECT 1496.0000 2381.9800 1497.6000 2382.4600 ;
        RECT 1480.4600 2376.5400 1482.0600 2377.0200 ;
        RECT 1480.4600 2381.9800 1482.0600 2382.4600 ;
        RECT 1496.0000 2360.2200 1497.6000 2360.7000 ;
        RECT 1496.0000 2365.6600 1497.6000 2366.1400 ;
        RECT 1496.0000 2371.1000 1497.6000 2371.5800 ;
        RECT 1480.4600 2360.2200 1482.0600 2360.7000 ;
        RECT 1480.4600 2365.6600 1482.0600 2366.1400 ;
        RECT 1480.4600 2371.1000 1482.0600 2371.5800 ;
        RECT 1435.4600 2403.7400 1437.0600 2404.2200 ;
        RECT 1435.4600 2409.1800 1437.0600 2409.6600 ;
        RECT 1435.4600 2387.4200 1437.0600 2387.9000 ;
        RECT 1435.4600 2392.8600 1437.0600 2393.3400 ;
        RECT 1435.4600 2398.3000 1437.0600 2398.7800 ;
        RECT 1435.4600 2376.5400 1437.0600 2377.0200 ;
        RECT 1435.4600 2381.9800 1437.0600 2382.4600 ;
        RECT 1435.4600 2360.2200 1437.0600 2360.7000 ;
        RECT 1435.4600 2365.6600 1437.0600 2366.1400 ;
        RECT 1435.4600 2371.1000 1437.0600 2371.5800 ;
        RECT 1435.4600 2414.6200 1437.0600 2415.1000 ;
        RECT 1480.4600 2414.6200 1482.0600 2415.1000 ;
        RECT 1496.0000 2414.6200 1497.6000 2415.1000 ;
        RECT 1390.4600 2447.2600 1392.0600 2447.7400 ;
        RECT 1390.4600 2452.7000 1392.0600 2453.1800 ;
        RECT 1390.4600 2458.1400 1392.0600 2458.6200 ;
        RECT 1345.4600 2447.2600 1347.0600 2447.7400 ;
        RECT 1345.4600 2452.7000 1347.0600 2453.1800 ;
        RECT 1345.4600 2458.1400 1347.0600 2458.6200 ;
        RECT 1390.4600 2430.9400 1392.0600 2431.4200 ;
        RECT 1390.4600 2436.3800 1392.0600 2436.8600 ;
        RECT 1390.4600 2420.0600 1392.0600 2420.5400 ;
        RECT 1390.4600 2425.5000 1392.0600 2425.9800 ;
        RECT 1345.4600 2430.9400 1347.0600 2431.4200 ;
        RECT 1345.4600 2436.3800 1347.0600 2436.8600 ;
        RECT 1345.4600 2420.0600 1347.0600 2420.5400 ;
        RECT 1345.4600 2425.5000 1347.0600 2425.9800 ;
        RECT 1345.4600 2441.8200 1347.0600 2442.3000 ;
        RECT 1390.4600 2441.8200 1392.0600 2442.3000 ;
        RECT 1293.3000 2458.1400 1294.9000 2458.6200 ;
        RECT 1300.4600 2458.1400 1302.0600 2458.6200 ;
        RECT 1300.4600 2447.2600 1302.0600 2447.7400 ;
        RECT 1300.4600 2452.7000 1302.0600 2453.1800 ;
        RECT 1293.3000 2447.2600 1294.9000 2447.7400 ;
        RECT 1293.3000 2452.7000 1294.9000 2453.1800 ;
        RECT 1300.4600 2430.9400 1302.0600 2431.4200 ;
        RECT 1300.4600 2436.3800 1302.0600 2436.8600 ;
        RECT 1293.3000 2430.9400 1294.9000 2431.4200 ;
        RECT 1293.3000 2436.3800 1294.9000 2436.8600 ;
        RECT 1300.4600 2420.0600 1302.0600 2420.5400 ;
        RECT 1300.4600 2425.5000 1302.0600 2425.9800 ;
        RECT 1293.3000 2420.0600 1294.9000 2420.5400 ;
        RECT 1293.3000 2425.5000 1294.9000 2425.9800 ;
        RECT 1293.3000 2441.8200 1294.9000 2442.3000 ;
        RECT 1300.4600 2441.8200 1302.0600 2442.3000 ;
        RECT 1390.4600 2403.7400 1392.0600 2404.2200 ;
        RECT 1390.4600 2409.1800 1392.0600 2409.6600 ;
        RECT 1390.4600 2387.4200 1392.0600 2387.9000 ;
        RECT 1390.4600 2392.8600 1392.0600 2393.3400 ;
        RECT 1390.4600 2398.3000 1392.0600 2398.7800 ;
        RECT 1345.4600 2403.7400 1347.0600 2404.2200 ;
        RECT 1345.4600 2409.1800 1347.0600 2409.6600 ;
        RECT 1345.4600 2387.4200 1347.0600 2387.9000 ;
        RECT 1345.4600 2392.8600 1347.0600 2393.3400 ;
        RECT 1345.4600 2398.3000 1347.0600 2398.7800 ;
        RECT 1390.4600 2376.5400 1392.0600 2377.0200 ;
        RECT 1390.4600 2381.9800 1392.0600 2382.4600 ;
        RECT 1390.4600 2360.2200 1392.0600 2360.7000 ;
        RECT 1390.4600 2365.6600 1392.0600 2366.1400 ;
        RECT 1390.4600 2371.1000 1392.0600 2371.5800 ;
        RECT 1345.4600 2376.5400 1347.0600 2377.0200 ;
        RECT 1345.4600 2381.9800 1347.0600 2382.4600 ;
        RECT 1345.4600 2360.2200 1347.0600 2360.7000 ;
        RECT 1345.4600 2365.6600 1347.0600 2366.1400 ;
        RECT 1345.4600 2371.1000 1347.0600 2371.5800 ;
        RECT 1300.4600 2403.7400 1302.0600 2404.2200 ;
        RECT 1300.4600 2409.1800 1302.0600 2409.6600 ;
        RECT 1293.3000 2403.7400 1294.9000 2404.2200 ;
        RECT 1293.3000 2409.1800 1294.9000 2409.6600 ;
        RECT 1300.4600 2387.4200 1302.0600 2387.9000 ;
        RECT 1300.4600 2392.8600 1302.0600 2393.3400 ;
        RECT 1300.4600 2398.3000 1302.0600 2398.7800 ;
        RECT 1293.3000 2387.4200 1294.9000 2387.9000 ;
        RECT 1293.3000 2392.8600 1294.9000 2393.3400 ;
        RECT 1293.3000 2398.3000 1294.9000 2398.7800 ;
        RECT 1300.4600 2376.5400 1302.0600 2377.0200 ;
        RECT 1300.4600 2381.9800 1302.0600 2382.4600 ;
        RECT 1293.3000 2376.5400 1294.9000 2377.0200 ;
        RECT 1293.3000 2381.9800 1294.9000 2382.4600 ;
        RECT 1300.4600 2360.2200 1302.0600 2360.7000 ;
        RECT 1300.4600 2365.6600 1302.0600 2366.1400 ;
        RECT 1300.4600 2371.1000 1302.0600 2371.5800 ;
        RECT 1293.3000 2360.2200 1294.9000 2360.7000 ;
        RECT 1293.3000 2365.6600 1294.9000 2366.1400 ;
        RECT 1293.3000 2371.1000 1294.9000 2371.5800 ;
        RECT 1293.3000 2414.6200 1294.9000 2415.1000 ;
        RECT 1300.4600 2414.6200 1302.0600 2415.1000 ;
        RECT 1345.4600 2414.6200 1347.0600 2415.1000 ;
        RECT 1390.4600 2414.6200 1392.0600 2415.1000 ;
        RECT 1496.0000 2349.3400 1497.6000 2349.8200 ;
        RECT 1496.0000 2354.7800 1497.6000 2355.2600 ;
        RECT 1480.4600 2349.3400 1482.0600 2349.8200 ;
        RECT 1480.4600 2354.7800 1482.0600 2355.2600 ;
        RECT 1496.0000 2333.0200 1497.6000 2333.5000 ;
        RECT 1496.0000 2338.4600 1497.6000 2338.9400 ;
        RECT 1496.0000 2343.9000 1497.6000 2344.3800 ;
        RECT 1480.4600 2333.0200 1482.0600 2333.5000 ;
        RECT 1480.4600 2338.4600 1482.0600 2338.9400 ;
        RECT 1480.4600 2343.9000 1482.0600 2344.3800 ;
        RECT 1496.0000 2322.1400 1497.6000 2322.6200 ;
        RECT 1496.0000 2327.5800 1497.6000 2328.0600 ;
        RECT 1480.4600 2322.1400 1482.0600 2322.6200 ;
        RECT 1480.4600 2327.5800 1482.0600 2328.0600 ;
        RECT 1496.0000 2305.8200 1497.6000 2306.3000 ;
        RECT 1496.0000 2311.2600 1497.6000 2311.7400 ;
        RECT 1496.0000 2316.7000 1497.6000 2317.1800 ;
        RECT 1480.4600 2305.8200 1482.0600 2306.3000 ;
        RECT 1480.4600 2311.2600 1482.0600 2311.7400 ;
        RECT 1480.4600 2316.7000 1482.0600 2317.1800 ;
        RECT 1435.4600 2349.3400 1437.0600 2349.8200 ;
        RECT 1435.4600 2354.7800 1437.0600 2355.2600 ;
        RECT 1435.4600 2333.0200 1437.0600 2333.5000 ;
        RECT 1435.4600 2338.4600 1437.0600 2338.9400 ;
        RECT 1435.4600 2343.9000 1437.0600 2344.3800 ;
        RECT 1435.4600 2322.1400 1437.0600 2322.6200 ;
        RECT 1435.4600 2327.5800 1437.0600 2328.0600 ;
        RECT 1435.4600 2305.8200 1437.0600 2306.3000 ;
        RECT 1435.4600 2311.2600 1437.0600 2311.7400 ;
        RECT 1435.4600 2316.7000 1437.0600 2317.1800 ;
        RECT 1496.0000 2294.9400 1497.6000 2295.4200 ;
        RECT 1496.0000 2300.3800 1497.6000 2300.8600 ;
        RECT 1480.4600 2294.9400 1482.0600 2295.4200 ;
        RECT 1480.4600 2300.3800 1482.0600 2300.8600 ;
        RECT 1496.0000 2278.6200 1497.6000 2279.1000 ;
        RECT 1496.0000 2284.0600 1497.6000 2284.5400 ;
        RECT 1496.0000 2289.5000 1497.6000 2289.9800 ;
        RECT 1480.4600 2278.6200 1482.0600 2279.1000 ;
        RECT 1480.4600 2284.0600 1482.0600 2284.5400 ;
        RECT 1480.4600 2289.5000 1482.0600 2289.9800 ;
        RECT 1496.0000 2267.7400 1497.6000 2268.2200 ;
        RECT 1496.0000 2273.1800 1497.6000 2273.6600 ;
        RECT 1480.4600 2267.7400 1482.0600 2268.2200 ;
        RECT 1480.4600 2273.1800 1482.0600 2273.6600 ;
        RECT 1480.4600 2262.3000 1482.0600 2262.7800 ;
        RECT 1496.0000 2262.3000 1497.6000 2262.7800 ;
        RECT 1435.4600 2294.9400 1437.0600 2295.4200 ;
        RECT 1435.4600 2300.3800 1437.0600 2300.8600 ;
        RECT 1435.4600 2278.6200 1437.0600 2279.1000 ;
        RECT 1435.4600 2284.0600 1437.0600 2284.5400 ;
        RECT 1435.4600 2289.5000 1437.0600 2289.9800 ;
        RECT 1435.4600 2267.7400 1437.0600 2268.2200 ;
        RECT 1435.4600 2273.1800 1437.0600 2273.6600 ;
        RECT 1435.4600 2262.3000 1437.0600 2262.7800 ;
        RECT 1390.4600 2349.3400 1392.0600 2349.8200 ;
        RECT 1390.4600 2354.7800 1392.0600 2355.2600 ;
        RECT 1390.4600 2333.0200 1392.0600 2333.5000 ;
        RECT 1390.4600 2338.4600 1392.0600 2338.9400 ;
        RECT 1390.4600 2343.9000 1392.0600 2344.3800 ;
        RECT 1345.4600 2349.3400 1347.0600 2349.8200 ;
        RECT 1345.4600 2354.7800 1347.0600 2355.2600 ;
        RECT 1345.4600 2333.0200 1347.0600 2333.5000 ;
        RECT 1345.4600 2338.4600 1347.0600 2338.9400 ;
        RECT 1345.4600 2343.9000 1347.0600 2344.3800 ;
        RECT 1390.4600 2322.1400 1392.0600 2322.6200 ;
        RECT 1390.4600 2327.5800 1392.0600 2328.0600 ;
        RECT 1390.4600 2305.8200 1392.0600 2306.3000 ;
        RECT 1390.4600 2311.2600 1392.0600 2311.7400 ;
        RECT 1390.4600 2316.7000 1392.0600 2317.1800 ;
        RECT 1345.4600 2322.1400 1347.0600 2322.6200 ;
        RECT 1345.4600 2327.5800 1347.0600 2328.0600 ;
        RECT 1345.4600 2305.8200 1347.0600 2306.3000 ;
        RECT 1345.4600 2311.2600 1347.0600 2311.7400 ;
        RECT 1345.4600 2316.7000 1347.0600 2317.1800 ;
        RECT 1300.4600 2349.3400 1302.0600 2349.8200 ;
        RECT 1300.4600 2354.7800 1302.0600 2355.2600 ;
        RECT 1293.3000 2349.3400 1294.9000 2349.8200 ;
        RECT 1293.3000 2354.7800 1294.9000 2355.2600 ;
        RECT 1300.4600 2333.0200 1302.0600 2333.5000 ;
        RECT 1300.4600 2338.4600 1302.0600 2338.9400 ;
        RECT 1300.4600 2343.9000 1302.0600 2344.3800 ;
        RECT 1293.3000 2333.0200 1294.9000 2333.5000 ;
        RECT 1293.3000 2338.4600 1294.9000 2338.9400 ;
        RECT 1293.3000 2343.9000 1294.9000 2344.3800 ;
        RECT 1300.4600 2322.1400 1302.0600 2322.6200 ;
        RECT 1300.4600 2327.5800 1302.0600 2328.0600 ;
        RECT 1293.3000 2322.1400 1294.9000 2322.6200 ;
        RECT 1293.3000 2327.5800 1294.9000 2328.0600 ;
        RECT 1300.4600 2305.8200 1302.0600 2306.3000 ;
        RECT 1300.4600 2311.2600 1302.0600 2311.7400 ;
        RECT 1300.4600 2316.7000 1302.0600 2317.1800 ;
        RECT 1293.3000 2305.8200 1294.9000 2306.3000 ;
        RECT 1293.3000 2311.2600 1294.9000 2311.7400 ;
        RECT 1293.3000 2316.7000 1294.9000 2317.1800 ;
        RECT 1390.4600 2294.9400 1392.0600 2295.4200 ;
        RECT 1390.4600 2300.3800 1392.0600 2300.8600 ;
        RECT 1390.4600 2278.6200 1392.0600 2279.1000 ;
        RECT 1390.4600 2284.0600 1392.0600 2284.5400 ;
        RECT 1390.4600 2289.5000 1392.0600 2289.9800 ;
        RECT 1345.4600 2294.9400 1347.0600 2295.4200 ;
        RECT 1345.4600 2300.3800 1347.0600 2300.8600 ;
        RECT 1345.4600 2278.6200 1347.0600 2279.1000 ;
        RECT 1345.4600 2284.0600 1347.0600 2284.5400 ;
        RECT 1345.4600 2289.5000 1347.0600 2289.9800 ;
        RECT 1390.4600 2273.1800 1392.0600 2273.6600 ;
        RECT 1390.4600 2267.7400 1392.0600 2268.2200 ;
        RECT 1390.4600 2262.3000 1392.0600 2262.7800 ;
        RECT 1345.4600 2273.1800 1347.0600 2273.6600 ;
        RECT 1345.4600 2267.7400 1347.0600 2268.2200 ;
        RECT 1345.4600 2262.3000 1347.0600 2262.7800 ;
        RECT 1300.4600 2294.9400 1302.0600 2295.4200 ;
        RECT 1300.4600 2300.3800 1302.0600 2300.8600 ;
        RECT 1293.3000 2294.9400 1294.9000 2295.4200 ;
        RECT 1293.3000 2300.3800 1294.9000 2300.8600 ;
        RECT 1300.4600 2278.6200 1302.0600 2279.1000 ;
        RECT 1300.4600 2284.0600 1302.0600 2284.5400 ;
        RECT 1300.4600 2289.5000 1302.0600 2289.9800 ;
        RECT 1293.3000 2278.6200 1294.9000 2279.1000 ;
        RECT 1293.3000 2284.0600 1294.9000 2284.5400 ;
        RECT 1293.3000 2289.5000 1294.9000 2289.9800 ;
        RECT 1300.4600 2267.7400 1302.0600 2268.2200 ;
        RECT 1300.4600 2273.1800 1302.0600 2273.6600 ;
        RECT 1293.3000 2267.7400 1294.9000 2268.2200 ;
        RECT 1293.3000 2273.1800 1294.9000 2273.6600 ;
        RECT 1293.3000 2262.3000 1294.9000 2262.7800 ;
        RECT 1300.4600 2262.3000 1302.0600 2262.7800 ;
        RECT 1290.3400 2464.4900 1500.5600 2466.0900 ;
        RECT 1290.3400 2252.7900 1500.5600 2254.3900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 2249.9600 1294.9000 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 2468.0000 1294.9000 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 2249.9600 1497.6000 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 2468.0000 1497.6000 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2252.7900 1291.9400 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2252.7900 1500.5600 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2464.4900 1291.9400 2466.0900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2464.4900 1500.5600 2466.0900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 2023.1500 1482.0600 2236.4500 ;
        RECT 1435.4600 2023.1500 1437.0600 2236.4500 ;
        RECT 1390.4600 2023.1500 1392.0600 2236.4500 ;
        RECT 1345.4600 2023.1500 1347.0600 2236.4500 ;
        RECT 1300.4600 2023.1500 1302.0600 2236.4500 ;
        RECT 1496.0000 2020.3200 1497.6000 2239.9600 ;
        RECT 1293.3000 2020.3200 1294.9000 2239.9600 ;
      LAYER met3 ;
        RECT 1480.4600 2228.5000 1482.0600 2228.9800 ;
        RECT 1496.0000 2228.5000 1497.6000 2228.9800 ;
        RECT 1496.0000 2217.6200 1497.6000 2218.1000 ;
        RECT 1496.0000 2223.0600 1497.6000 2223.5400 ;
        RECT 1480.4600 2217.6200 1482.0600 2218.1000 ;
        RECT 1480.4600 2223.0600 1482.0600 2223.5400 ;
        RECT 1496.0000 2201.3000 1497.6000 2201.7800 ;
        RECT 1496.0000 2206.7400 1497.6000 2207.2200 ;
        RECT 1480.4600 2201.3000 1482.0600 2201.7800 ;
        RECT 1480.4600 2206.7400 1482.0600 2207.2200 ;
        RECT 1496.0000 2190.4200 1497.6000 2190.9000 ;
        RECT 1496.0000 2195.8600 1497.6000 2196.3400 ;
        RECT 1480.4600 2190.4200 1482.0600 2190.9000 ;
        RECT 1480.4600 2195.8600 1482.0600 2196.3400 ;
        RECT 1480.4600 2212.1800 1482.0600 2212.6600 ;
        RECT 1496.0000 2212.1800 1497.6000 2212.6600 ;
        RECT 1435.4600 2217.6200 1437.0600 2218.1000 ;
        RECT 1435.4600 2223.0600 1437.0600 2223.5400 ;
        RECT 1435.4600 2228.5000 1437.0600 2228.9800 ;
        RECT 1435.4600 2201.3000 1437.0600 2201.7800 ;
        RECT 1435.4600 2206.7400 1437.0600 2207.2200 ;
        RECT 1435.4600 2195.8600 1437.0600 2196.3400 ;
        RECT 1435.4600 2190.4200 1437.0600 2190.9000 ;
        RECT 1435.4600 2212.1800 1437.0600 2212.6600 ;
        RECT 1496.0000 2174.1000 1497.6000 2174.5800 ;
        RECT 1496.0000 2179.5400 1497.6000 2180.0200 ;
        RECT 1480.4600 2174.1000 1482.0600 2174.5800 ;
        RECT 1480.4600 2179.5400 1482.0600 2180.0200 ;
        RECT 1496.0000 2157.7800 1497.6000 2158.2600 ;
        RECT 1496.0000 2163.2200 1497.6000 2163.7000 ;
        RECT 1496.0000 2168.6600 1497.6000 2169.1400 ;
        RECT 1480.4600 2157.7800 1482.0600 2158.2600 ;
        RECT 1480.4600 2163.2200 1482.0600 2163.7000 ;
        RECT 1480.4600 2168.6600 1482.0600 2169.1400 ;
        RECT 1496.0000 2146.9000 1497.6000 2147.3800 ;
        RECT 1496.0000 2152.3400 1497.6000 2152.8200 ;
        RECT 1480.4600 2146.9000 1482.0600 2147.3800 ;
        RECT 1480.4600 2152.3400 1482.0600 2152.8200 ;
        RECT 1496.0000 2130.5800 1497.6000 2131.0600 ;
        RECT 1496.0000 2136.0200 1497.6000 2136.5000 ;
        RECT 1496.0000 2141.4600 1497.6000 2141.9400 ;
        RECT 1480.4600 2130.5800 1482.0600 2131.0600 ;
        RECT 1480.4600 2136.0200 1482.0600 2136.5000 ;
        RECT 1480.4600 2141.4600 1482.0600 2141.9400 ;
        RECT 1435.4600 2174.1000 1437.0600 2174.5800 ;
        RECT 1435.4600 2179.5400 1437.0600 2180.0200 ;
        RECT 1435.4600 2157.7800 1437.0600 2158.2600 ;
        RECT 1435.4600 2163.2200 1437.0600 2163.7000 ;
        RECT 1435.4600 2168.6600 1437.0600 2169.1400 ;
        RECT 1435.4600 2146.9000 1437.0600 2147.3800 ;
        RECT 1435.4600 2152.3400 1437.0600 2152.8200 ;
        RECT 1435.4600 2130.5800 1437.0600 2131.0600 ;
        RECT 1435.4600 2136.0200 1437.0600 2136.5000 ;
        RECT 1435.4600 2141.4600 1437.0600 2141.9400 ;
        RECT 1435.4600 2184.9800 1437.0600 2185.4600 ;
        RECT 1480.4600 2184.9800 1482.0600 2185.4600 ;
        RECT 1496.0000 2184.9800 1497.6000 2185.4600 ;
        RECT 1390.4600 2217.6200 1392.0600 2218.1000 ;
        RECT 1390.4600 2223.0600 1392.0600 2223.5400 ;
        RECT 1390.4600 2228.5000 1392.0600 2228.9800 ;
        RECT 1345.4600 2217.6200 1347.0600 2218.1000 ;
        RECT 1345.4600 2223.0600 1347.0600 2223.5400 ;
        RECT 1345.4600 2228.5000 1347.0600 2228.9800 ;
        RECT 1390.4600 2201.3000 1392.0600 2201.7800 ;
        RECT 1390.4600 2206.7400 1392.0600 2207.2200 ;
        RECT 1390.4600 2190.4200 1392.0600 2190.9000 ;
        RECT 1390.4600 2195.8600 1392.0600 2196.3400 ;
        RECT 1345.4600 2201.3000 1347.0600 2201.7800 ;
        RECT 1345.4600 2206.7400 1347.0600 2207.2200 ;
        RECT 1345.4600 2190.4200 1347.0600 2190.9000 ;
        RECT 1345.4600 2195.8600 1347.0600 2196.3400 ;
        RECT 1345.4600 2212.1800 1347.0600 2212.6600 ;
        RECT 1390.4600 2212.1800 1392.0600 2212.6600 ;
        RECT 1293.3000 2228.5000 1294.9000 2228.9800 ;
        RECT 1300.4600 2228.5000 1302.0600 2228.9800 ;
        RECT 1300.4600 2217.6200 1302.0600 2218.1000 ;
        RECT 1300.4600 2223.0600 1302.0600 2223.5400 ;
        RECT 1293.3000 2217.6200 1294.9000 2218.1000 ;
        RECT 1293.3000 2223.0600 1294.9000 2223.5400 ;
        RECT 1300.4600 2201.3000 1302.0600 2201.7800 ;
        RECT 1300.4600 2206.7400 1302.0600 2207.2200 ;
        RECT 1293.3000 2201.3000 1294.9000 2201.7800 ;
        RECT 1293.3000 2206.7400 1294.9000 2207.2200 ;
        RECT 1300.4600 2190.4200 1302.0600 2190.9000 ;
        RECT 1300.4600 2195.8600 1302.0600 2196.3400 ;
        RECT 1293.3000 2190.4200 1294.9000 2190.9000 ;
        RECT 1293.3000 2195.8600 1294.9000 2196.3400 ;
        RECT 1293.3000 2212.1800 1294.9000 2212.6600 ;
        RECT 1300.4600 2212.1800 1302.0600 2212.6600 ;
        RECT 1390.4600 2174.1000 1392.0600 2174.5800 ;
        RECT 1390.4600 2179.5400 1392.0600 2180.0200 ;
        RECT 1390.4600 2157.7800 1392.0600 2158.2600 ;
        RECT 1390.4600 2163.2200 1392.0600 2163.7000 ;
        RECT 1390.4600 2168.6600 1392.0600 2169.1400 ;
        RECT 1345.4600 2174.1000 1347.0600 2174.5800 ;
        RECT 1345.4600 2179.5400 1347.0600 2180.0200 ;
        RECT 1345.4600 2157.7800 1347.0600 2158.2600 ;
        RECT 1345.4600 2163.2200 1347.0600 2163.7000 ;
        RECT 1345.4600 2168.6600 1347.0600 2169.1400 ;
        RECT 1390.4600 2146.9000 1392.0600 2147.3800 ;
        RECT 1390.4600 2152.3400 1392.0600 2152.8200 ;
        RECT 1390.4600 2130.5800 1392.0600 2131.0600 ;
        RECT 1390.4600 2136.0200 1392.0600 2136.5000 ;
        RECT 1390.4600 2141.4600 1392.0600 2141.9400 ;
        RECT 1345.4600 2146.9000 1347.0600 2147.3800 ;
        RECT 1345.4600 2152.3400 1347.0600 2152.8200 ;
        RECT 1345.4600 2130.5800 1347.0600 2131.0600 ;
        RECT 1345.4600 2136.0200 1347.0600 2136.5000 ;
        RECT 1345.4600 2141.4600 1347.0600 2141.9400 ;
        RECT 1300.4600 2174.1000 1302.0600 2174.5800 ;
        RECT 1300.4600 2179.5400 1302.0600 2180.0200 ;
        RECT 1293.3000 2174.1000 1294.9000 2174.5800 ;
        RECT 1293.3000 2179.5400 1294.9000 2180.0200 ;
        RECT 1300.4600 2157.7800 1302.0600 2158.2600 ;
        RECT 1300.4600 2163.2200 1302.0600 2163.7000 ;
        RECT 1300.4600 2168.6600 1302.0600 2169.1400 ;
        RECT 1293.3000 2157.7800 1294.9000 2158.2600 ;
        RECT 1293.3000 2163.2200 1294.9000 2163.7000 ;
        RECT 1293.3000 2168.6600 1294.9000 2169.1400 ;
        RECT 1300.4600 2146.9000 1302.0600 2147.3800 ;
        RECT 1300.4600 2152.3400 1302.0600 2152.8200 ;
        RECT 1293.3000 2146.9000 1294.9000 2147.3800 ;
        RECT 1293.3000 2152.3400 1294.9000 2152.8200 ;
        RECT 1300.4600 2130.5800 1302.0600 2131.0600 ;
        RECT 1300.4600 2136.0200 1302.0600 2136.5000 ;
        RECT 1300.4600 2141.4600 1302.0600 2141.9400 ;
        RECT 1293.3000 2130.5800 1294.9000 2131.0600 ;
        RECT 1293.3000 2136.0200 1294.9000 2136.5000 ;
        RECT 1293.3000 2141.4600 1294.9000 2141.9400 ;
        RECT 1293.3000 2184.9800 1294.9000 2185.4600 ;
        RECT 1300.4600 2184.9800 1302.0600 2185.4600 ;
        RECT 1345.4600 2184.9800 1347.0600 2185.4600 ;
        RECT 1390.4600 2184.9800 1392.0600 2185.4600 ;
        RECT 1496.0000 2119.7000 1497.6000 2120.1800 ;
        RECT 1496.0000 2125.1400 1497.6000 2125.6200 ;
        RECT 1480.4600 2119.7000 1482.0600 2120.1800 ;
        RECT 1480.4600 2125.1400 1482.0600 2125.6200 ;
        RECT 1496.0000 2103.3800 1497.6000 2103.8600 ;
        RECT 1496.0000 2108.8200 1497.6000 2109.3000 ;
        RECT 1496.0000 2114.2600 1497.6000 2114.7400 ;
        RECT 1480.4600 2103.3800 1482.0600 2103.8600 ;
        RECT 1480.4600 2108.8200 1482.0600 2109.3000 ;
        RECT 1480.4600 2114.2600 1482.0600 2114.7400 ;
        RECT 1496.0000 2092.5000 1497.6000 2092.9800 ;
        RECT 1496.0000 2097.9400 1497.6000 2098.4200 ;
        RECT 1480.4600 2092.5000 1482.0600 2092.9800 ;
        RECT 1480.4600 2097.9400 1482.0600 2098.4200 ;
        RECT 1496.0000 2076.1800 1497.6000 2076.6600 ;
        RECT 1496.0000 2081.6200 1497.6000 2082.1000 ;
        RECT 1496.0000 2087.0600 1497.6000 2087.5400 ;
        RECT 1480.4600 2076.1800 1482.0600 2076.6600 ;
        RECT 1480.4600 2081.6200 1482.0600 2082.1000 ;
        RECT 1480.4600 2087.0600 1482.0600 2087.5400 ;
        RECT 1435.4600 2119.7000 1437.0600 2120.1800 ;
        RECT 1435.4600 2125.1400 1437.0600 2125.6200 ;
        RECT 1435.4600 2103.3800 1437.0600 2103.8600 ;
        RECT 1435.4600 2108.8200 1437.0600 2109.3000 ;
        RECT 1435.4600 2114.2600 1437.0600 2114.7400 ;
        RECT 1435.4600 2092.5000 1437.0600 2092.9800 ;
        RECT 1435.4600 2097.9400 1437.0600 2098.4200 ;
        RECT 1435.4600 2076.1800 1437.0600 2076.6600 ;
        RECT 1435.4600 2081.6200 1437.0600 2082.1000 ;
        RECT 1435.4600 2087.0600 1437.0600 2087.5400 ;
        RECT 1496.0000 2065.3000 1497.6000 2065.7800 ;
        RECT 1496.0000 2070.7400 1497.6000 2071.2200 ;
        RECT 1480.4600 2065.3000 1482.0600 2065.7800 ;
        RECT 1480.4600 2070.7400 1482.0600 2071.2200 ;
        RECT 1496.0000 2048.9800 1497.6000 2049.4600 ;
        RECT 1496.0000 2054.4200 1497.6000 2054.9000 ;
        RECT 1496.0000 2059.8600 1497.6000 2060.3400 ;
        RECT 1480.4600 2048.9800 1482.0600 2049.4600 ;
        RECT 1480.4600 2054.4200 1482.0600 2054.9000 ;
        RECT 1480.4600 2059.8600 1482.0600 2060.3400 ;
        RECT 1496.0000 2038.1000 1497.6000 2038.5800 ;
        RECT 1496.0000 2043.5400 1497.6000 2044.0200 ;
        RECT 1480.4600 2038.1000 1482.0600 2038.5800 ;
        RECT 1480.4600 2043.5400 1482.0600 2044.0200 ;
        RECT 1480.4600 2032.6600 1482.0600 2033.1400 ;
        RECT 1496.0000 2032.6600 1497.6000 2033.1400 ;
        RECT 1435.4600 2065.3000 1437.0600 2065.7800 ;
        RECT 1435.4600 2070.7400 1437.0600 2071.2200 ;
        RECT 1435.4600 2048.9800 1437.0600 2049.4600 ;
        RECT 1435.4600 2054.4200 1437.0600 2054.9000 ;
        RECT 1435.4600 2059.8600 1437.0600 2060.3400 ;
        RECT 1435.4600 2038.1000 1437.0600 2038.5800 ;
        RECT 1435.4600 2043.5400 1437.0600 2044.0200 ;
        RECT 1435.4600 2032.6600 1437.0600 2033.1400 ;
        RECT 1390.4600 2119.7000 1392.0600 2120.1800 ;
        RECT 1390.4600 2125.1400 1392.0600 2125.6200 ;
        RECT 1390.4600 2103.3800 1392.0600 2103.8600 ;
        RECT 1390.4600 2108.8200 1392.0600 2109.3000 ;
        RECT 1390.4600 2114.2600 1392.0600 2114.7400 ;
        RECT 1345.4600 2119.7000 1347.0600 2120.1800 ;
        RECT 1345.4600 2125.1400 1347.0600 2125.6200 ;
        RECT 1345.4600 2103.3800 1347.0600 2103.8600 ;
        RECT 1345.4600 2108.8200 1347.0600 2109.3000 ;
        RECT 1345.4600 2114.2600 1347.0600 2114.7400 ;
        RECT 1390.4600 2092.5000 1392.0600 2092.9800 ;
        RECT 1390.4600 2097.9400 1392.0600 2098.4200 ;
        RECT 1390.4600 2076.1800 1392.0600 2076.6600 ;
        RECT 1390.4600 2081.6200 1392.0600 2082.1000 ;
        RECT 1390.4600 2087.0600 1392.0600 2087.5400 ;
        RECT 1345.4600 2092.5000 1347.0600 2092.9800 ;
        RECT 1345.4600 2097.9400 1347.0600 2098.4200 ;
        RECT 1345.4600 2076.1800 1347.0600 2076.6600 ;
        RECT 1345.4600 2081.6200 1347.0600 2082.1000 ;
        RECT 1345.4600 2087.0600 1347.0600 2087.5400 ;
        RECT 1300.4600 2119.7000 1302.0600 2120.1800 ;
        RECT 1300.4600 2125.1400 1302.0600 2125.6200 ;
        RECT 1293.3000 2119.7000 1294.9000 2120.1800 ;
        RECT 1293.3000 2125.1400 1294.9000 2125.6200 ;
        RECT 1300.4600 2103.3800 1302.0600 2103.8600 ;
        RECT 1300.4600 2108.8200 1302.0600 2109.3000 ;
        RECT 1300.4600 2114.2600 1302.0600 2114.7400 ;
        RECT 1293.3000 2103.3800 1294.9000 2103.8600 ;
        RECT 1293.3000 2108.8200 1294.9000 2109.3000 ;
        RECT 1293.3000 2114.2600 1294.9000 2114.7400 ;
        RECT 1300.4600 2092.5000 1302.0600 2092.9800 ;
        RECT 1300.4600 2097.9400 1302.0600 2098.4200 ;
        RECT 1293.3000 2092.5000 1294.9000 2092.9800 ;
        RECT 1293.3000 2097.9400 1294.9000 2098.4200 ;
        RECT 1300.4600 2076.1800 1302.0600 2076.6600 ;
        RECT 1300.4600 2081.6200 1302.0600 2082.1000 ;
        RECT 1300.4600 2087.0600 1302.0600 2087.5400 ;
        RECT 1293.3000 2076.1800 1294.9000 2076.6600 ;
        RECT 1293.3000 2081.6200 1294.9000 2082.1000 ;
        RECT 1293.3000 2087.0600 1294.9000 2087.5400 ;
        RECT 1390.4600 2065.3000 1392.0600 2065.7800 ;
        RECT 1390.4600 2070.7400 1392.0600 2071.2200 ;
        RECT 1390.4600 2048.9800 1392.0600 2049.4600 ;
        RECT 1390.4600 2054.4200 1392.0600 2054.9000 ;
        RECT 1390.4600 2059.8600 1392.0600 2060.3400 ;
        RECT 1345.4600 2065.3000 1347.0600 2065.7800 ;
        RECT 1345.4600 2070.7400 1347.0600 2071.2200 ;
        RECT 1345.4600 2048.9800 1347.0600 2049.4600 ;
        RECT 1345.4600 2054.4200 1347.0600 2054.9000 ;
        RECT 1345.4600 2059.8600 1347.0600 2060.3400 ;
        RECT 1390.4600 2043.5400 1392.0600 2044.0200 ;
        RECT 1390.4600 2038.1000 1392.0600 2038.5800 ;
        RECT 1390.4600 2032.6600 1392.0600 2033.1400 ;
        RECT 1345.4600 2043.5400 1347.0600 2044.0200 ;
        RECT 1345.4600 2038.1000 1347.0600 2038.5800 ;
        RECT 1345.4600 2032.6600 1347.0600 2033.1400 ;
        RECT 1300.4600 2065.3000 1302.0600 2065.7800 ;
        RECT 1300.4600 2070.7400 1302.0600 2071.2200 ;
        RECT 1293.3000 2065.3000 1294.9000 2065.7800 ;
        RECT 1293.3000 2070.7400 1294.9000 2071.2200 ;
        RECT 1300.4600 2048.9800 1302.0600 2049.4600 ;
        RECT 1300.4600 2054.4200 1302.0600 2054.9000 ;
        RECT 1300.4600 2059.8600 1302.0600 2060.3400 ;
        RECT 1293.3000 2048.9800 1294.9000 2049.4600 ;
        RECT 1293.3000 2054.4200 1294.9000 2054.9000 ;
        RECT 1293.3000 2059.8600 1294.9000 2060.3400 ;
        RECT 1300.4600 2038.1000 1302.0600 2038.5800 ;
        RECT 1300.4600 2043.5400 1302.0600 2044.0200 ;
        RECT 1293.3000 2038.1000 1294.9000 2038.5800 ;
        RECT 1293.3000 2043.5400 1294.9000 2044.0200 ;
        RECT 1293.3000 2032.6600 1294.9000 2033.1400 ;
        RECT 1300.4600 2032.6600 1302.0600 2033.1400 ;
        RECT 1290.3400 2234.8500 1500.5600 2236.4500 ;
        RECT 1290.3400 2023.1500 1500.5600 2024.7500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 2020.3200 1294.9000 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 2238.3600 1294.9000 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 2020.3200 1497.6000 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 2238.3600 1497.6000 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2023.1500 1291.9400 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2023.1500 1500.5600 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2234.8500 1291.9400 2236.4500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2234.8500 1500.5600 2236.4500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 1793.5100 1482.0600 2006.8100 ;
        RECT 1435.4600 1793.5100 1437.0600 2006.8100 ;
        RECT 1390.4600 1793.5100 1392.0600 2006.8100 ;
        RECT 1345.4600 1793.5100 1347.0600 2006.8100 ;
        RECT 1300.4600 1793.5100 1302.0600 2006.8100 ;
        RECT 1496.0000 1790.6800 1497.6000 2010.3200 ;
        RECT 1293.3000 1790.6800 1294.9000 2010.3200 ;
      LAYER met3 ;
        RECT 1480.4600 1998.8600 1482.0600 1999.3400 ;
        RECT 1496.0000 1998.8600 1497.6000 1999.3400 ;
        RECT 1496.0000 1987.9800 1497.6000 1988.4600 ;
        RECT 1496.0000 1993.4200 1497.6000 1993.9000 ;
        RECT 1480.4600 1987.9800 1482.0600 1988.4600 ;
        RECT 1480.4600 1993.4200 1482.0600 1993.9000 ;
        RECT 1496.0000 1971.6600 1497.6000 1972.1400 ;
        RECT 1496.0000 1977.1000 1497.6000 1977.5800 ;
        RECT 1480.4600 1971.6600 1482.0600 1972.1400 ;
        RECT 1480.4600 1977.1000 1482.0600 1977.5800 ;
        RECT 1496.0000 1960.7800 1497.6000 1961.2600 ;
        RECT 1496.0000 1966.2200 1497.6000 1966.7000 ;
        RECT 1480.4600 1960.7800 1482.0600 1961.2600 ;
        RECT 1480.4600 1966.2200 1482.0600 1966.7000 ;
        RECT 1480.4600 1982.5400 1482.0600 1983.0200 ;
        RECT 1496.0000 1982.5400 1497.6000 1983.0200 ;
        RECT 1435.4600 1987.9800 1437.0600 1988.4600 ;
        RECT 1435.4600 1993.4200 1437.0600 1993.9000 ;
        RECT 1435.4600 1998.8600 1437.0600 1999.3400 ;
        RECT 1435.4600 1971.6600 1437.0600 1972.1400 ;
        RECT 1435.4600 1977.1000 1437.0600 1977.5800 ;
        RECT 1435.4600 1966.2200 1437.0600 1966.7000 ;
        RECT 1435.4600 1960.7800 1437.0600 1961.2600 ;
        RECT 1435.4600 1982.5400 1437.0600 1983.0200 ;
        RECT 1496.0000 1944.4600 1497.6000 1944.9400 ;
        RECT 1496.0000 1949.9000 1497.6000 1950.3800 ;
        RECT 1480.4600 1944.4600 1482.0600 1944.9400 ;
        RECT 1480.4600 1949.9000 1482.0600 1950.3800 ;
        RECT 1496.0000 1928.1400 1497.6000 1928.6200 ;
        RECT 1496.0000 1933.5800 1497.6000 1934.0600 ;
        RECT 1496.0000 1939.0200 1497.6000 1939.5000 ;
        RECT 1480.4600 1928.1400 1482.0600 1928.6200 ;
        RECT 1480.4600 1933.5800 1482.0600 1934.0600 ;
        RECT 1480.4600 1939.0200 1482.0600 1939.5000 ;
        RECT 1496.0000 1917.2600 1497.6000 1917.7400 ;
        RECT 1496.0000 1922.7000 1497.6000 1923.1800 ;
        RECT 1480.4600 1917.2600 1482.0600 1917.7400 ;
        RECT 1480.4600 1922.7000 1482.0600 1923.1800 ;
        RECT 1496.0000 1900.9400 1497.6000 1901.4200 ;
        RECT 1496.0000 1906.3800 1497.6000 1906.8600 ;
        RECT 1496.0000 1911.8200 1497.6000 1912.3000 ;
        RECT 1480.4600 1900.9400 1482.0600 1901.4200 ;
        RECT 1480.4600 1906.3800 1482.0600 1906.8600 ;
        RECT 1480.4600 1911.8200 1482.0600 1912.3000 ;
        RECT 1435.4600 1944.4600 1437.0600 1944.9400 ;
        RECT 1435.4600 1949.9000 1437.0600 1950.3800 ;
        RECT 1435.4600 1928.1400 1437.0600 1928.6200 ;
        RECT 1435.4600 1933.5800 1437.0600 1934.0600 ;
        RECT 1435.4600 1939.0200 1437.0600 1939.5000 ;
        RECT 1435.4600 1917.2600 1437.0600 1917.7400 ;
        RECT 1435.4600 1922.7000 1437.0600 1923.1800 ;
        RECT 1435.4600 1900.9400 1437.0600 1901.4200 ;
        RECT 1435.4600 1906.3800 1437.0600 1906.8600 ;
        RECT 1435.4600 1911.8200 1437.0600 1912.3000 ;
        RECT 1435.4600 1955.3400 1437.0600 1955.8200 ;
        RECT 1480.4600 1955.3400 1482.0600 1955.8200 ;
        RECT 1496.0000 1955.3400 1497.6000 1955.8200 ;
        RECT 1390.4600 1987.9800 1392.0600 1988.4600 ;
        RECT 1390.4600 1993.4200 1392.0600 1993.9000 ;
        RECT 1390.4600 1998.8600 1392.0600 1999.3400 ;
        RECT 1345.4600 1987.9800 1347.0600 1988.4600 ;
        RECT 1345.4600 1993.4200 1347.0600 1993.9000 ;
        RECT 1345.4600 1998.8600 1347.0600 1999.3400 ;
        RECT 1390.4600 1971.6600 1392.0600 1972.1400 ;
        RECT 1390.4600 1977.1000 1392.0600 1977.5800 ;
        RECT 1390.4600 1960.7800 1392.0600 1961.2600 ;
        RECT 1390.4600 1966.2200 1392.0600 1966.7000 ;
        RECT 1345.4600 1971.6600 1347.0600 1972.1400 ;
        RECT 1345.4600 1977.1000 1347.0600 1977.5800 ;
        RECT 1345.4600 1960.7800 1347.0600 1961.2600 ;
        RECT 1345.4600 1966.2200 1347.0600 1966.7000 ;
        RECT 1345.4600 1982.5400 1347.0600 1983.0200 ;
        RECT 1390.4600 1982.5400 1392.0600 1983.0200 ;
        RECT 1293.3000 1998.8600 1294.9000 1999.3400 ;
        RECT 1300.4600 1998.8600 1302.0600 1999.3400 ;
        RECT 1300.4600 1987.9800 1302.0600 1988.4600 ;
        RECT 1300.4600 1993.4200 1302.0600 1993.9000 ;
        RECT 1293.3000 1987.9800 1294.9000 1988.4600 ;
        RECT 1293.3000 1993.4200 1294.9000 1993.9000 ;
        RECT 1300.4600 1971.6600 1302.0600 1972.1400 ;
        RECT 1300.4600 1977.1000 1302.0600 1977.5800 ;
        RECT 1293.3000 1971.6600 1294.9000 1972.1400 ;
        RECT 1293.3000 1977.1000 1294.9000 1977.5800 ;
        RECT 1300.4600 1960.7800 1302.0600 1961.2600 ;
        RECT 1300.4600 1966.2200 1302.0600 1966.7000 ;
        RECT 1293.3000 1960.7800 1294.9000 1961.2600 ;
        RECT 1293.3000 1966.2200 1294.9000 1966.7000 ;
        RECT 1293.3000 1982.5400 1294.9000 1983.0200 ;
        RECT 1300.4600 1982.5400 1302.0600 1983.0200 ;
        RECT 1390.4600 1944.4600 1392.0600 1944.9400 ;
        RECT 1390.4600 1949.9000 1392.0600 1950.3800 ;
        RECT 1390.4600 1928.1400 1392.0600 1928.6200 ;
        RECT 1390.4600 1933.5800 1392.0600 1934.0600 ;
        RECT 1390.4600 1939.0200 1392.0600 1939.5000 ;
        RECT 1345.4600 1944.4600 1347.0600 1944.9400 ;
        RECT 1345.4600 1949.9000 1347.0600 1950.3800 ;
        RECT 1345.4600 1928.1400 1347.0600 1928.6200 ;
        RECT 1345.4600 1933.5800 1347.0600 1934.0600 ;
        RECT 1345.4600 1939.0200 1347.0600 1939.5000 ;
        RECT 1390.4600 1917.2600 1392.0600 1917.7400 ;
        RECT 1390.4600 1922.7000 1392.0600 1923.1800 ;
        RECT 1390.4600 1900.9400 1392.0600 1901.4200 ;
        RECT 1390.4600 1906.3800 1392.0600 1906.8600 ;
        RECT 1390.4600 1911.8200 1392.0600 1912.3000 ;
        RECT 1345.4600 1917.2600 1347.0600 1917.7400 ;
        RECT 1345.4600 1922.7000 1347.0600 1923.1800 ;
        RECT 1345.4600 1900.9400 1347.0600 1901.4200 ;
        RECT 1345.4600 1906.3800 1347.0600 1906.8600 ;
        RECT 1345.4600 1911.8200 1347.0600 1912.3000 ;
        RECT 1300.4600 1944.4600 1302.0600 1944.9400 ;
        RECT 1300.4600 1949.9000 1302.0600 1950.3800 ;
        RECT 1293.3000 1944.4600 1294.9000 1944.9400 ;
        RECT 1293.3000 1949.9000 1294.9000 1950.3800 ;
        RECT 1300.4600 1928.1400 1302.0600 1928.6200 ;
        RECT 1300.4600 1933.5800 1302.0600 1934.0600 ;
        RECT 1300.4600 1939.0200 1302.0600 1939.5000 ;
        RECT 1293.3000 1928.1400 1294.9000 1928.6200 ;
        RECT 1293.3000 1933.5800 1294.9000 1934.0600 ;
        RECT 1293.3000 1939.0200 1294.9000 1939.5000 ;
        RECT 1300.4600 1917.2600 1302.0600 1917.7400 ;
        RECT 1300.4600 1922.7000 1302.0600 1923.1800 ;
        RECT 1293.3000 1917.2600 1294.9000 1917.7400 ;
        RECT 1293.3000 1922.7000 1294.9000 1923.1800 ;
        RECT 1300.4600 1900.9400 1302.0600 1901.4200 ;
        RECT 1300.4600 1906.3800 1302.0600 1906.8600 ;
        RECT 1300.4600 1911.8200 1302.0600 1912.3000 ;
        RECT 1293.3000 1900.9400 1294.9000 1901.4200 ;
        RECT 1293.3000 1906.3800 1294.9000 1906.8600 ;
        RECT 1293.3000 1911.8200 1294.9000 1912.3000 ;
        RECT 1293.3000 1955.3400 1294.9000 1955.8200 ;
        RECT 1300.4600 1955.3400 1302.0600 1955.8200 ;
        RECT 1345.4600 1955.3400 1347.0600 1955.8200 ;
        RECT 1390.4600 1955.3400 1392.0600 1955.8200 ;
        RECT 1496.0000 1890.0600 1497.6000 1890.5400 ;
        RECT 1496.0000 1895.5000 1497.6000 1895.9800 ;
        RECT 1480.4600 1890.0600 1482.0600 1890.5400 ;
        RECT 1480.4600 1895.5000 1482.0600 1895.9800 ;
        RECT 1496.0000 1873.7400 1497.6000 1874.2200 ;
        RECT 1496.0000 1879.1800 1497.6000 1879.6600 ;
        RECT 1496.0000 1884.6200 1497.6000 1885.1000 ;
        RECT 1480.4600 1873.7400 1482.0600 1874.2200 ;
        RECT 1480.4600 1879.1800 1482.0600 1879.6600 ;
        RECT 1480.4600 1884.6200 1482.0600 1885.1000 ;
        RECT 1496.0000 1862.8600 1497.6000 1863.3400 ;
        RECT 1496.0000 1868.3000 1497.6000 1868.7800 ;
        RECT 1480.4600 1862.8600 1482.0600 1863.3400 ;
        RECT 1480.4600 1868.3000 1482.0600 1868.7800 ;
        RECT 1496.0000 1846.5400 1497.6000 1847.0200 ;
        RECT 1496.0000 1851.9800 1497.6000 1852.4600 ;
        RECT 1496.0000 1857.4200 1497.6000 1857.9000 ;
        RECT 1480.4600 1846.5400 1482.0600 1847.0200 ;
        RECT 1480.4600 1851.9800 1482.0600 1852.4600 ;
        RECT 1480.4600 1857.4200 1482.0600 1857.9000 ;
        RECT 1435.4600 1890.0600 1437.0600 1890.5400 ;
        RECT 1435.4600 1895.5000 1437.0600 1895.9800 ;
        RECT 1435.4600 1873.7400 1437.0600 1874.2200 ;
        RECT 1435.4600 1879.1800 1437.0600 1879.6600 ;
        RECT 1435.4600 1884.6200 1437.0600 1885.1000 ;
        RECT 1435.4600 1862.8600 1437.0600 1863.3400 ;
        RECT 1435.4600 1868.3000 1437.0600 1868.7800 ;
        RECT 1435.4600 1846.5400 1437.0600 1847.0200 ;
        RECT 1435.4600 1851.9800 1437.0600 1852.4600 ;
        RECT 1435.4600 1857.4200 1437.0600 1857.9000 ;
        RECT 1496.0000 1835.6600 1497.6000 1836.1400 ;
        RECT 1496.0000 1841.1000 1497.6000 1841.5800 ;
        RECT 1480.4600 1835.6600 1482.0600 1836.1400 ;
        RECT 1480.4600 1841.1000 1482.0600 1841.5800 ;
        RECT 1496.0000 1819.3400 1497.6000 1819.8200 ;
        RECT 1496.0000 1824.7800 1497.6000 1825.2600 ;
        RECT 1496.0000 1830.2200 1497.6000 1830.7000 ;
        RECT 1480.4600 1819.3400 1482.0600 1819.8200 ;
        RECT 1480.4600 1824.7800 1482.0600 1825.2600 ;
        RECT 1480.4600 1830.2200 1482.0600 1830.7000 ;
        RECT 1496.0000 1808.4600 1497.6000 1808.9400 ;
        RECT 1496.0000 1813.9000 1497.6000 1814.3800 ;
        RECT 1480.4600 1808.4600 1482.0600 1808.9400 ;
        RECT 1480.4600 1813.9000 1482.0600 1814.3800 ;
        RECT 1480.4600 1803.0200 1482.0600 1803.5000 ;
        RECT 1496.0000 1803.0200 1497.6000 1803.5000 ;
        RECT 1435.4600 1835.6600 1437.0600 1836.1400 ;
        RECT 1435.4600 1841.1000 1437.0600 1841.5800 ;
        RECT 1435.4600 1819.3400 1437.0600 1819.8200 ;
        RECT 1435.4600 1824.7800 1437.0600 1825.2600 ;
        RECT 1435.4600 1830.2200 1437.0600 1830.7000 ;
        RECT 1435.4600 1808.4600 1437.0600 1808.9400 ;
        RECT 1435.4600 1813.9000 1437.0600 1814.3800 ;
        RECT 1435.4600 1803.0200 1437.0600 1803.5000 ;
        RECT 1390.4600 1890.0600 1392.0600 1890.5400 ;
        RECT 1390.4600 1895.5000 1392.0600 1895.9800 ;
        RECT 1390.4600 1873.7400 1392.0600 1874.2200 ;
        RECT 1390.4600 1879.1800 1392.0600 1879.6600 ;
        RECT 1390.4600 1884.6200 1392.0600 1885.1000 ;
        RECT 1345.4600 1890.0600 1347.0600 1890.5400 ;
        RECT 1345.4600 1895.5000 1347.0600 1895.9800 ;
        RECT 1345.4600 1873.7400 1347.0600 1874.2200 ;
        RECT 1345.4600 1879.1800 1347.0600 1879.6600 ;
        RECT 1345.4600 1884.6200 1347.0600 1885.1000 ;
        RECT 1390.4600 1862.8600 1392.0600 1863.3400 ;
        RECT 1390.4600 1868.3000 1392.0600 1868.7800 ;
        RECT 1390.4600 1846.5400 1392.0600 1847.0200 ;
        RECT 1390.4600 1851.9800 1392.0600 1852.4600 ;
        RECT 1390.4600 1857.4200 1392.0600 1857.9000 ;
        RECT 1345.4600 1862.8600 1347.0600 1863.3400 ;
        RECT 1345.4600 1868.3000 1347.0600 1868.7800 ;
        RECT 1345.4600 1846.5400 1347.0600 1847.0200 ;
        RECT 1345.4600 1851.9800 1347.0600 1852.4600 ;
        RECT 1345.4600 1857.4200 1347.0600 1857.9000 ;
        RECT 1300.4600 1890.0600 1302.0600 1890.5400 ;
        RECT 1300.4600 1895.5000 1302.0600 1895.9800 ;
        RECT 1293.3000 1890.0600 1294.9000 1890.5400 ;
        RECT 1293.3000 1895.5000 1294.9000 1895.9800 ;
        RECT 1300.4600 1873.7400 1302.0600 1874.2200 ;
        RECT 1300.4600 1879.1800 1302.0600 1879.6600 ;
        RECT 1300.4600 1884.6200 1302.0600 1885.1000 ;
        RECT 1293.3000 1873.7400 1294.9000 1874.2200 ;
        RECT 1293.3000 1879.1800 1294.9000 1879.6600 ;
        RECT 1293.3000 1884.6200 1294.9000 1885.1000 ;
        RECT 1300.4600 1862.8600 1302.0600 1863.3400 ;
        RECT 1300.4600 1868.3000 1302.0600 1868.7800 ;
        RECT 1293.3000 1862.8600 1294.9000 1863.3400 ;
        RECT 1293.3000 1868.3000 1294.9000 1868.7800 ;
        RECT 1300.4600 1846.5400 1302.0600 1847.0200 ;
        RECT 1300.4600 1851.9800 1302.0600 1852.4600 ;
        RECT 1300.4600 1857.4200 1302.0600 1857.9000 ;
        RECT 1293.3000 1846.5400 1294.9000 1847.0200 ;
        RECT 1293.3000 1851.9800 1294.9000 1852.4600 ;
        RECT 1293.3000 1857.4200 1294.9000 1857.9000 ;
        RECT 1390.4600 1835.6600 1392.0600 1836.1400 ;
        RECT 1390.4600 1841.1000 1392.0600 1841.5800 ;
        RECT 1390.4600 1819.3400 1392.0600 1819.8200 ;
        RECT 1390.4600 1824.7800 1392.0600 1825.2600 ;
        RECT 1390.4600 1830.2200 1392.0600 1830.7000 ;
        RECT 1345.4600 1835.6600 1347.0600 1836.1400 ;
        RECT 1345.4600 1841.1000 1347.0600 1841.5800 ;
        RECT 1345.4600 1819.3400 1347.0600 1819.8200 ;
        RECT 1345.4600 1824.7800 1347.0600 1825.2600 ;
        RECT 1345.4600 1830.2200 1347.0600 1830.7000 ;
        RECT 1390.4600 1813.9000 1392.0600 1814.3800 ;
        RECT 1390.4600 1808.4600 1392.0600 1808.9400 ;
        RECT 1390.4600 1803.0200 1392.0600 1803.5000 ;
        RECT 1345.4600 1813.9000 1347.0600 1814.3800 ;
        RECT 1345.4600 1808.4600 1347.0600 1808.9400 ;
        RECT 1345.4600 1803.0200 1347.0600 1803.5000 ;
        RECT 1300.4600 1835.6600 1302.0600 1836.1400 ;
        RECT 1300.4600 1841.1000 1302.0600 1841.5800 ;
        RECT 1293.3000 1835.6600 1294.9000 1836.1400 ;
        RECT 1293.3000 1841.1000 1294.9000 1841.5800 ;
        RECT 1300.4600 1819.3400 1302.0600 1819.8200 ;
        RECT 1300.4600 1824.7800 1302.0600 1825.2600 ;
        RECT 1300.4600 1830.2200 1302.0600 1830.7000 ;
        RECT 1293.3000 1819.3400 1294.9000 1819.8200 ;
        RECT 1293.3000 1824.7800 1294.9000 1825.2600 ;
        RECT 1293.3000 1830.2200 1294.9000 1830.7000 ;
        RECT 1300.4600 1808.4600 1302.0600 1808.9400 ;
        RECT 1300.4600 1813.9000 1302.0600 1814.3800 ;
        RECT 1293.3000 1808.4600 1294.9000 1808.9400 ;
        RECT 1293.3000 1813.9000 1294.9000 1814.3800 ;
        RECT 1293.3000 1803.0200 1294.9000 1803.5000 ;
        RECT 1300.4600 1803.0200 1302.0600 1803.5000 ;
        RECT 1290.3400 2005.2100 1500.5600 2006.8100 ;
        RECT 1290.3400 1793.5100 1500.5600 1795.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1790.6800 1294.9000 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 2008.7200 1294.9000 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1790.6800 1497.6000 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 2008.7200 1497.6000 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1793.5100 1291.9400 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1793.5100 1500.5600 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2005.2100 1291.9400 2006.8100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2005.2100 1500.5600 2006.8100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 1563.8700 1482.0600 1777.1700 ;
        RECT 1435.4600 1563.8700 1437.0600 1777.1700 ;
        RECT 1390.4600 1563.8700 1392.0600 1777.1700 ;
        RECT 1345.4600 1563.8700 1347.0600 1777.1700 ;
        RECT 1300.4600 1563.8700 1302.0600 1777.1700 ;
        RECT 1496.0000 1561.0400 1497.6000 1780.6800 ;
        RECT 1293.3000 1561.0400 1294.9000 1780.6800 ;
      LAYER met3 ;
        RECT 1480.4600 1769.2200 1482.0600 1769.7000 ;
        RECT 1496.0000 1769.2200 1497.6000 1769.7000 ;
        RECT 1496.0000 1758.3400 1497.6000 1758.8200 ;
        RECT 1496.0000 1763.7800 1497.6000 1764.2600 ;
        RECT 1480.4600 1758.3400 1482.0600 1758.8200 ;
        RECT 1480.4600 1763.7800 1482.0600 1764.2600 ;
        RECT 1496.0000 1742.0200 1497.6000 1742.5000 ;
        RECT 1496.0000 1747.4600 1497.6000 1747.9400 ;
        RECT 1480.4600 1742.0200 1482.0600 1742.5000 ;
        RECT 1480.4600 1747.4600 1482.0600 1747.9400 ;
        RECT 1496.0000 1731.1400 1497.6000 1731.6200 ;
        RECT 1496.0000 1736.5800 1497.6000 1737.0600 ;
        RECT 1480.4600 1731.1400 1482.0600 1731.6200 ;
        RECT 1480.4600 1736.5800 1482.0600 1737.0600 ;
        RECT 1480.4600 1752.9000 1482.0600 1753.3800 ;
        RECT 1496.0000 1752.9000 1497.6000 1753.3800 ;
        RECT 1435.4600 1758.3400 1437.0600 1758.8200 ;
        RECT 1435.4600 1763.7800 1437.0600 1764.2600 ;
        RECT 1435.4600 1769.2200 1437.0600 1769.7000 ;
        RECT 1435.4600 1742.0200 1437.0600 1742.5000 ;
        RECT 1435.4600 1747.4600 1437.0600 1747.9400 ;
        RECT 1435.4600 1736.5800 1437.0600 1737.0600 ;
        RECT 1435.4600 1731.1400 1437.0600 1731.6200 ;
        RECT 1435.4600 1752.9000 1437.0600 1753.3800 ;
        RECT 1496.0000 1714.8200 1497.6000 1715.3000 ;
        RECT 1496.0000 1720.2600 1497.6000 1720.7400 ;
        RECT 1480.4600 1714.8200 1482.0600 1715.3000 ;
        RECT 1480.4600 1720.2600 1482.0600 1720.7400 ;
        RECT 1496.0000 1698.5000 1497.6000 1698.9800 ;
        RECT 1496.0000 1703.9400 1497.6000 1704.4200 ;
        RECT 1496.0000 1709.3800 1497.6000 1709.8600 ;
        RECT 1480.4600 1698.5000 1482.0600 1698.9800 ;
        RECT 1480.4600 1703.9400 1482.0600 1704.4200 ;
        RECT 1480.4600 1709.3800 1482.0600 1709.8600 ;
        RECT 1496.0000 1687.6200 1497.6000 1688.1000 ;
        RECT 1496.0000 1693.0600 1497.6000 1693.5400 ;
        RECT 1480.4600 1687.6200 1482.0600 1688.1000 ;
        RECT 1480.4600 1693.0600 1482.0600 1693.5400 ;
        RECT 1496.0000 1671.3000 1497.6000 1671.7800 ;
        RECT 1496.0000 1676.7400 1497.6000 1677.2200 ;
        RECT 1496.0000 1682.1800 1497.6000 1682.6600 ;
        RECT 1480.4600 1671.3000 1482.0600 1671.7800 ;
        RECT 1480.4600 1676.7400 1482.0600 1677.2200 ;
        RECT 1480.4600 1682.1800 1482.0600 1682.6600 ;
        RECT 1435.4600 1714.8200 1437.0600 1715.3000 ;
        RECT 1435.4600 1720.2600 1437.0600 1720.7400 ;
        RECT 1435.4600 1698.5000 1437.0600 1698.9800 ;
        RECT 1435.4600 1703.9400 1437.0600 1704.4200 ;
        RECT 1435.4600 1709.3800 1437.0600 1709.8600 ;
        RECT 1435.4600 1687.6200 1437.0600 1688.1000 ;
        RECT 1435.4600 1693.0600 1437.0600 1693.5400 ;
        RECT 1435.4600 1671.3000 1437.0600 1671.7800 ;
        RECT 1435.4600 1676.7400 1437.0600 1677.2200 ;
        RECT 1435.4600 1682.1800 1437.0600 1682.6600 ;
        RECT 1435.4600 1725.7000 1437.0600 1726.1800 ;
        RECT 1480.4600 1725.7000 1482.0600 1726.1800 ;
        RECT 1496.0000 1725.7000 1497.6000 1726.1800 ;
        RECT 1390.4600 1758.3400 1392.0600 1758.8200 ;
        RECT 1390.4600 1763.7800 1392.0600 1764.2600 ;
        RECT 1390.4600 1769.2200 1392.0600 1769.7000 ;
        RECT 1345.4600 1758.3400 1347.0600 1758.8200 ;
        RECT 1345.4600 1763.7800 1347.0600 1764.2600 ;
        RECT 1345.4600 1769.2200 1347.0600 1769.7000 ;
        RECT 1390.4600 1742.0200 1392.0600 1742.5000 ;
        RECT 1390.4600 1747.4600 1392.0600 1747.9400 ;
        RECT 1390.4600 1731.1400 1392.0600 1731.6200 ;
        RECT 1390.4600 1736.5800 1392.0600 1737.0600 ;
        RECT 1345.4600 1742.0200 1347.0600 1742.5000 ;
        RECT 1345.4600 1747.4600 1347.0600 1747.9400 ;
        RECT 1345.4600 1731.1400 1347.0600 1731.6200 ;
        RECT 1345.4600 1736.5800 1347.0600 1737.0600 ;
        RECT 1345.4600 1752.9000 1347.0600 1753.3800 ;
        RECT 1390.4600 1752.9000 1392.0600 1753.3800 ;
        RECT 1293.3000 1769.2200 1294.9000 1769.7000 ;
        RECT 1300.4600 1769.2200 1302.0600 1769.7000 ;
        RECT 1300.4600 1758.3400 1302.0600 1758.8200 ;
        RECT 1300.4600 1763.7800 1302.0600 1764.2600 ;
        RECT 1293.3000 1758.3400 1294.9000 1758.8200 ;
        RECT 1293.3000 1763.7800 1294.9000 1764.2600 ;
        RECT 1300.4600 1742.0200 1302.0600 1742.5000 ;
        RECT 1300.4600 1747.4600 1302.0600 1747.9400 ;
        RECT 1293.3000 1742.0200 1294.9000 1742.5000 ;
        RECT 1293.3000 1747.4600 1294.9000 1747.9400 ;
        RECT 1300.4600 1731.1400 1302.0600 1731.6200 ;
        RECT 1300.4600 1736.5800 1302.0600 1737.0600 ;
        RECT 1293.3000 1731.1400 1294.9000 1731.6200 ;
        RECT 1293.3000 1736.5800 1294.9000 1737.0600 ;
        RECT 1293.3000 1752.9000 1294.9000 1753.3800 ;
        RECT 1300.4600 1752.9000 1302.0600 1753.3800 ;
        RECT 1390.4600 1714.8200 1392.0600 1715.3000 ;
        RECT 1390.4600 1720.2600 1392.0600 1720.7400 ;
        RECT 1390.4600 1698.5000 1392.0600 1698.9800 ;
        RECT 1390.4600 1703.9400 1392.0600 1704.4200 ;
        RECT 1390.4600 1709.3800 1392.0600 1709.8600 ;
        RECT 1345.4600 1714.8200 1347.0600 1715.3000 ;
        RECT 1345.4600 1720.2600 1347.0600 1720.7400 ;
        RECT 1345.4600 1698.5000 1347.0600 1698.9800 ;
        RECT 1345.4600 1703.9400 1347.0600 1704.4200 ;
        RECT 1345.4600 1709.3800 1347.0600 1709.8600 ;
        RECT 1390.4600 1687.6200 1392.0600 1688.1000 ;
        RECT 1390.4600 1693.0600 1392.0600 1693.5400 ;
        RECT 1390.4600 1671.3000 1392.0600 1671.7800 ;
        RECT 1390.4600 1676.7400 1392.0600 1677.2200 ;
        RECT 1390.4600 1682.1800 1392.0600 1682.6600 ;
        RECT 1345.4600 1687.6200 1347.0600 1688.1000 ;
        RECT 1345.4600 1693.0600 1347.0600 1693.5400 ;
        RECT 1345.4600 1671.3000 1347.0600 1671.7800 ;
        RECT 1345.4600 1676.7400 1347.0600 1677.2200 ;
        RECT 1345.4600 1682.1800 1347.0600 1682.6600 ;
        RECT 1300.4600 1714.8200 1302.0600 1715.3000 ;
        RECT 1300.4600 1720.2600 1302.0600 1720.7400 ;
        RECT 1293.3000 1714.8200 1294.9000 1715.3000 ;
        RECT 1293.3000 1720.2600 1294.9000 1720.7400 ;
        RECT 1300.4600 1698.5000 1302.0600 1698.9800 ;
        RECT 1300.4600 1703.9400 1302.0600 1704.4200 ;
        RECT 1300.4600 1709.3800 1302.0600 1709.8600 ;
        RECT 1293.3000 1698.5000 1294.9000 1698.9800 ;
        RECT 1293.3000 1703.9400 1294.9000 1704.4200 ;
        RECT 1293.3000 1709.3800 1294.9000 1709.8600 ;
        RECT 1300.4600 1687.6200 1302.0600 1688.1000 ;
        RECT 1300.4600 1693.0600 1302.0600 1693.5400 ;
        RECT 1293.3000 1687.6200 1294.9000 1688.1000 ;
        RECT 1293.3000 1693.0600 1294.9000 1693.5400 ;
        RECT 1300.4600 1671.3000 1302.0600 1671.7800 ;
        RECT 1300.4600 1676.7400 1302.0600 1677.2200 ;
        RECT 1300.4600 1682.1800 1302.0600 1682.6600 ;
        RECT 1293.3000 1671.3000 1294.9000 1671.7800 ;
        RECT 1293.3000 1676.7400 1294.9000 1677.2200 ;
        RECT 1293.3000 1682.1800 1294.9000 1682.6600 ;
        RECT 1293.3000 1725.7000 1294.9000 1726.1800 ;
        RECT 1300.4600 1725.7000 1302.0600 1726.1800 ;
        RECT 1345.4600 1725.7000 1347.0600 1726.1800 ;
        RECT 1390.4600 1725.7000 1392.0600 1726.1800 ;
        RECT 1496.0000 1660.4200 1497.6000 1660.9000 ;
        RECT 1496.0000 1665.8600 1497.6000 1666.3400 ;
        RECT 1480.4600 1660.4200 1482.0600 1660.9000 ;
        RECT 1480.4600 1665.8600 1482.0600 1666.3400 ;
        RECT 1496.0000 1644.1000 1497.6000 1644.5800 ;
        RECT 1496.0000 1649.5400 1497.6000 1650.0200 ;
        RECT 1496.0000 1654.9800 1497.6000 1655.4600 ;
        RECT 1480.4600 1644.1000 1482.0600 1644.5800 ;
        RECT 1480.4600 1649.5400 1482.0600 1650.0200 ;
        RECT 1480.4600 1654.9800 1482.0600 1655.4600 ;
        RECT 1496.0000 1633.2200 1497.6000 1633.7000 ;
        RECT 1496.0000 1638.6600 1497.6000 1639.1400 ;
        RECT 1480.4600 1633.2200 1482.0600 1633.7000 ;
        RECT 1480.4600 1638.6600 1482.0600 1639.1400 ;
        RECT 1496.0000 1616.9000 1497.6000 1617.3800 ;
        RECT 1496.0000 1622.3400 1497.6000 1622.8200 ;
        RECT 1496.0000 1627.7800 1497.6000 1628.2600 ;
        RECT 1480.4600 1616.9000 1482.0600 1617.3800 ;
        RECT 1480.4600 1622.3400 1482.0600 1622.8200 ;
        RECT 1480.4600 1627.7800 1482.0600 1628.2600 ;
        RECT 1435.4600 1660.4200 1437.0600 1660.9000 ;
        RECT 1435.4600 1665.8600 1437.0600 1666.3400 ;
        RECT 1435.4600 1644.1000 1437.0600 1644.5800 ;
        RECT 1435.4600 1649.5400 1437.0600 1650.0200 ;
        RECT 1435.4600 1654.9800 1437.0600 1655.4600 ;
        RECT 1435.4600 1633.2200 1437.0600 1633.7000 ;
        RECT 1435.4600 1638.6600 1437.0600 1639.1400 ;
        RECT 1435.4600 1616.9000 1437.0600 1617.3800 ;
        RECT 1435.4600 1622.3400 1437.0600 1622.8200 ;
        RECT 1435.4600 1627.7800 1437.0600 1628.2600 ;
        RECT 1496.0000 1606.0200 1497.6000 1606.5000 ;
        RECT 1496.0000 1611.4600 1497.6000 1611.9400 ;
        RECT 1480.4600 1606.0200 1482.0600 1606.5000 ;
        RECT 1480.4600 1611.4600 1482.0600 1611.9400 ;
        RECT 1496.0000 1589.7000 1497.6000 1590.1800 ;
        RECT 1496.0000 1595.1400 1497.6000 1595.6200 ;
        RECT 1496.0000 1600.5800 1497.6000 1601.0600 ;
        RECT 1480.4600 1589.7000 1482.0600 1590.1800 ;
        RECT 1480.4600 1595.1400 1482.0600 1595.6200 ;
        RECT 1480.4600 1600.5800 1482.0600 1601.0600 ;
        RECT 1496.0000 1578.8200 1497.6000 1579.3000 ;
        RECT 1496.0000 1584.2600 1497.6000 1584.7400 ;
        RECT 1480.4600 1578.8200 1482.0600 1579.3000 ;
        RECT 1480.4600 1584.2600 1482.0600 1584.7400 ;
        RECT 1480.4600 1573.3800 1482.0600 1573.8600 ;
        RECT 1496.0000 1573.3800 1497.6000 1573.8600 ;
        RECT 1435.4600 1606.0200 1437.0600 1606.5000 ;
        RECT 1435.4600 1611.4600 1437.0600 1611.9400 ;
        RECT 1435.4600 1589.7000 1437.0600 1590.1800 ;
        RECT 1435.4600 1595.1400 1437.0600 1595.6200 ;
        RECT 1435.4600 1600.5800 1437.0600 1601.0600 ;
        RECT 1435.4600 1578.8200 1437.0600 1579.3000 ;
        RECT 1435.4600 1584.2600 1437.0600 1584.7400 ;
        RECT 1435.4600 1573.3800 1437.0600 1573.8600 ;
        RECT 1390.4600 1660.4200 1392.0600 1660.9000 ;
        RECT 1390.4600 1665.8600 1392.0600 1666.3400 ;
        RECT 1390.4600 1644.1000 1392.0600 1644.5800 ;
        RECT 1390.4600 1649.5400 1392.0600 1650.0200 ;
        RECT 1390.4600 1654.9800 1392.0600 1655.4600 ;
        RECT 1345.4600 1660.4200 1347.0600 1660.9000 ;
        RECT 1345.4600 1665.8600 1347.0600 1666.3400 ;
        RECT 1345.4600 1644.1000 1347.0600 1644.5800 ;
        RECT 1345.4600 1649.5400 1347.0600 1650.0200 ;
        RECT 1345.4600 1654.9800 1347.0600 1655.4600 ;
        RECT 1390.4600 1633.2200 1392.0600 1633.7000 ;
        RECT 1390.4600 1638.6600 1392.0600 1639.1400 ;
        RECT 1390.4600 1616.9000 1392.0600 1617.3800 ;
        RECT 1390.4600 1622.3400 1392.0600 1622.8200 ;
        RECT 1390.4600 1627.7800 1392.0600 1628.2600 ;
        RECT 1345.4600 1633.2200 1347.0600 1633.7000 ;
        RECT 1345.4600 1638.6600 1347.0600 1639.1400 ;
        RECT 1345.4600 1616.9000 1347.0600 1617.3800 ;
        RECT 1345.4600 1622.3400 1347.0600 1622.8200 ;
        RECT 1345.4600 1627.7800 1347.0600 1628.2600 ;
        RECT 1300.4600 1660.4200 1302.0600 1660.9000 ;
        RECT 1300.4600 1665.8600 1302.0600 1666.3400 ;
        RECT 1293.3000 1660.4200 1294.9000 1660.9000 ;
        RECT 1293.3000 1665.8600 1294.9000 1666.3400 ;
        RECT 1300.4600 1644.1000 1302.0600 1644.5800 ;
        RECT 1300.4600 1649.5400 1302.0600 1650.0200 ;
        RECT 1300.4600 1654.9800 1302.0600 1655.4600 ;
        RECT 1293.3000 1644.1000 1294.9000 1644.5800 ;
        RECT 1293.3000 1649.5400 1294.9000 1650.0200 ;
        RECT 1293.3000 1654.9800 1294.9000 1655.4600 ;
        RECT 1300.4600 1633.2200 1302.0600 1633.7000 ;
        RECT 1300.4600 1638.6600 1302.0600 1639.1400 ;
        RECT 1293.3000 1633.2200 1294.9000 1633.7000 ;
        RECT 1293.3000 1638.6600 1294.9000 1639.1400 ;
        RECT 1300.4600 1616.9000 1302.0600 1617.3800 ;
        RECT 1300.4600 1622.3400 1302.0600 1622.8200 ;
        RECT 1300.4600 1627.7800 1302.0600 1628.2600 ;
        RECT 1293.3000 1616.9000 1294.9000 1617.3800 ;
        RECT 1293.3000 1622.3400 1294.9000 1622.8200 ;
        RECT 1293.3000 1627.7800 1294.9000 1628.2600 ;
        RECT 1390.4600 1606.0200 1392.0600 1606.5000 ;
        RECT 1390.4600 1611.4600 1392.0600 1611.9400 ;
        RECT 1390.4600 1589.7000 1392.0600 1590.1800 ;
        RECT 1390.4600 1595.1400 1392.0600 1595.6200 ;
        RECT 1390.4600 1600.5800 1392.0600 1601.0600 ;
        RECT 1345.4600 1606.0200 1347.0600 1606.5000 ;
        RECT 1345.4600 1611.4600 1347.0600 1611.9400 ;
        RECT 1345.4600 1589.7000 1347.0600 1590.1800 ;
        RECT 1345.4600 1595.1400 1347.0600 1595.6200 ;
        RECT 1345.4600 1600.5800 1347.0600 1601.0600 ;
        RECT 1390.4600 1584.2600 1392.0600 1584.7400 ;
        RECT 1390.4600 1578.8200 1392.0600 1579.3000 ;
        RECT 1390.4600 1573.3800 1392.0600 1573.8600 ;
        RECT 1345.4600 1584.2600 1347.0600 1584.7400 ;
        RECT 1345.4600 1578.8200 1347.0600 1579.3000 ;
        RECT 1345.4600 1573.3800 1347.0600 1573.8600 ;
        RECT 1300.4600 1606.0200 1302.0600 1606.5000 ;
        RECT 1300.4600 1611.4600 1302.0600 1611.9400 ;
        RECT 1293.3000 1606.0200 1294.9000 1606.5000 ;
        RECT 1293.3000 1611.4600 1294.9000 1611.9400 ;
        RECT 1300.4600 1589.7000 1302.0600 1590.1800 ;
        RECT 1300.4600 1595.1400 1302.0600 1595.6200 ;
        RECT 1300.4600 1600.5800 1302.0600 1601.0600 ;
        RECT 1293.3000 1589.7000 1294.9000 1590.1800 ;
        RECT 1293.3000 1595.1400 1294.9000 1595.6200 ;
        RECT 1293.3000 1600.5800 1294.9000 1601.0600 ;
        RECT 1300.4600 1578.8200 1302.0600 1579.3000 ;
        RECT 1300.4600 1584.2600 1302.0600 1584.7400 ;
        RECT 1293.3000 1578.8200 1294.9000 1579.3000 ;
        RECT 1293.3000 1584.2600 1294.9000 1584.7400 ;
        RECT 1293.3000 1573.3800 1294.9000 1573.8600 ;
        RECT 1300.4600 1573.3800 1302.0600 1573.8600 ;
        RECT 1290.3400 1775.5700 1500.5600 1777.1700 ;
        RECT 1290.3400 1563.8700 1500.5600 1565.4700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1561.0400 1294.9000 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1779.0800 1294.9000 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1561.0400 1497.6000 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1779.0800 1497.6000 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1563.8700 1291.9400 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1563.8700 1500.5600 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1775.5700 1291.9400 1777.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1775.5700 1500.5600 1777.1700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 1334.2300 1482.0600 1547.5300 ;
        RECT 1435.4600 1334.2300 1437.0600 1547.5300 ;
        RECT 1390.4600 1334.2300 1392.0600 1547.5300 ;
        RECT 1345.4600 1334.2300 1347.0600 1547.5300 ;
        RECT 1300.4600 1334.2300 1302.0600 1547.5300 ;
        RECT 1496.0000 1331.4000 1497.6000 1551.0400 ;
        RECT 1293.3000 1331.4000 1294.9000 1551.0400 ;
      LAYER met3 ;
        RECT 1480.4600 1539.5800 1482.0600 1540.0600 ;
        RECT 1496.0000 1539.5800 1497.6000 1540.0600 ;
        RECT 1496.0000 1528.7000 1497.6000 1529.1800 ;
        RECT 1496.0000 1534.1400 1497.6000 1534.6200 ;
        RECT 1480.4600 1528.7000 1482.0600 1529.1800 ;
        RECT 1480.4600 1534.1400 1482.0600 1534.6200 ;
        RECT 1496.0000 1512.3800 1497.6000 1512.8600 ;
        RECT 1496.0000 1517.8200 1497.6000 1518.3000 ;
        RECT 1480.4600 1512.3800 1482.0600 1512.8600 ;
        RECT 1480.4600 1517.8200 1482.0600 1518.3000 ;
        RECT 1496.0000 1501.5000 1497.6000 1501.9800 ;
        RECT 1496.0000 1506.9400 1497.6000 1507.4200 ;
        RECT 1480.4600 1501.5000 1482.0600 1501.9800 ;
        RECT 1480.4600 1506.9400 1482.0600 1507.4200 ;
        RECT 1480.4600 1523.2600 1482.0600 1523.7400 ;
        RECT 1496.0000 1523.2600 1497.6000 1523.7400 ;
        RECT 1435.4600 1528.7000 1437.0600 1529.1800 ;
        RECT 1435.4600 1534.1400 1437.0600 1534.6200 ;
        RECT 1435.4600 1539.5800 1437.0600 1540.0600 ;
        RECT 1435.4600 1512.3800 1437.0600 1512.8600 ;
        RECT 1435.4600 1517.8200 1437.0600 1518.3000 ;
        RECT 1435.4600 1506.9400 1437.0600 1507.4200 ;
        RECT 1435.4600 1501.5000 1437.0600 1501.9800 ;
        RECT 1435.4600 1523.2600 1437.0600 1523.7400 ;
        RECT 1496.0000 1485.1800 1497.6000 1485.6600 ;
        RECT 1496.0000 1490.6200 1497.6000 1491.1000 ;
        RECT 1480.4600 1485.1800 1482.0600 1485.6600 ;
        RECT 1480.4600 1490.6200 1482.0600 1491.1000 ;
        RECT 1496.0000 1468.8600 1497.6000 1469.3400 ;
        RECT 1496.0000 1474.3000 1497.6000 1474.7800 ;
        RECT 1496.0000 1479.7400 1497.6000 1480.2200 ;
        RECT 1480.4600 1468.8600 1482.0600 1469.3400 ;
        RECT 1480.4600 1474.3000 1482.0600 1474.7800 ;
        RECT 1480.4600 1479.7400 1482.0600 1480.2200 ;
        RECT 1496.0000 1457.9800 1497.6000 1458.4600 ;
        RECT 1496.0000 1463.4200 1497.6000 1463.9000 ;
        RECT 1480.4600 1457.9800 1482.0600 1458.4600 ;
        RECT 1480.4600 1463.4200 1482.0600 1463.9000 ;
        RECT 1496.0000 1441.6600 1497.6000 1442.1400 ;
        RECT 1496.0000 1447.1000 1497.6000 1447.5800 ;
        RECT 1496.0000 1452.5400 1497.6000 1453.0200 ;
        RECT 1480.4600 1441.6600 1482.0600 1442.1400 ;
        RECT 1480.4600 1447.1000 1482.0600 1447.5800 ;
        RECT 1480.4600 1452.5400 1482.0600 1453.0200 ;
        RECT 1435.4600 1485.1800 1437.0600 1485.6600 ;
        RECT 1435.4600 1490.6200 1437.0600 1491.1000 ;
        RECT 1435.4600 1468.8600 1437.0600 1469.3400 ;
        RECT 1435.4600 1474.3000 1437.0600 1474.7800 ;
        RECT 1435.4600 1479.7400 1437.0600 1480.2200 ;
        RECT 1435.4600 1457.9800 1437.0600 1458.4600 ;
        RECT 1435.4600 1463.4200 1437.0600 1463.9000 ;
        RECT 1435.4600 1441.6600 1437.0600 1442.1400 ;
        RECT 1435.4600 1447.1000 1437.0600 1447.5800 ;
        RECT 1435.4600 1452.5400 1437.0600 1453.0200 ;
        RECT 1435.4600 1496.0600 1437.0600 1496.5400 ;
        RECT 1480.4600 1496.0600 1482.0600 1496.5400 ;
        RECT 1496.0000 1496.0600 1497.6000 1496.5400 ;
        RECT 1390.4600 1528.7000 1392.0600 1529.1800 ;
        RECT 1390.4600 1534.1400 1392.0600 1534.6200 ;
        RECT 1390.4600 1539.5800 1392.0600 1540.0600 ;
        RECT 1345.4600 1528.7000 1347.0600 1529.1800 ;
        RECT 1345.4600 1534.1400 1347.0600 1534.6200 ;
        RECT 1345.4600 1539.5800 1347.0600 1540.0600 ;
        RECT 1390.4600 1512.3800 1392.0600 1512.8600 ;
        RECT 1390.4600 1517.8200 1392.0600 1518.3000 ;
        RECT 1390.4600 1501.5000 1392.0600 1501.9800 ;
        RECT 1390.4600 1506.9400 1392.0600 1507.4200 ;
        RECT 1345.4600 1512.3800 1347.0600 1512.8600 ;
        RECT 1345.4600 1517.8200 1347.0600 1518.3000 ;
        RECT 1345.4600 1501.5000 1347.0600 1501.9800 ;
        RECT 1345.4600 1506.9400 1347.0600 1507.4200 ;
        RECT 1345.4600 1523.2600 1347.0600 1523.7400 ;
        RECT 1390.4600 1523.2600 1392.0600 1523.7400 ;
        RECT 1293.3000 1539.5800 1294.9000 1540.0600 ;
        RECT 1300.4600 1539.5800 1302.0600 1540.0600 ;
        RECT 1300.4600 1528.7000 1302.0600 1529.1800 ;
        RECT 1300.4600 1534.1400 1302.0600 1534.6200 ;
        RECT 1293.3000 1528.7000 1294.9000 1529.1800 ;
        RECT 1293.3000 1534.1400 1294.9000 1534.6200 ;
        RECT 1300.4600 1512.3800 1302.0600 1512.8600 ;
        RECT 1300.4600 1517.8200 1302.0600 1518.3000 ;
        RECT 1293.3000 1512.3800 1294.9000 1512.8600 ;
        RECT 1293.3000 1517.8200 1294.9000 1518.3000 ;
        RECT 1300.4600 1501.5000 1302.0600 1501.9800 ;
        RECT 1300.4600 1506.9400 1302.0600 1507.4200 ;
        RECT 1293.3000 1501.5000 1294.9000 1501.9800 ;
        RECT 1293.3000 1506.9400 1294.9000 1507.4200 ;
        RECT 1293.3000 1523.2600 1294.9000 1523.7400 ;
        RECT 1300.4600 1523.2600 1302.0600 1523.7400 ;
        RECT 1390.4600 1485.1800 1392.0600 1485.6600 ;
        RECT 1390.4600 1490.6200 1392.0600 1491.1000 ;
        RECT 1390.4600 1468.8600 1392.0600 1469.3400 ;
        RECT 1390.4600 1474.3000 1392.0600 1474.7800 ;
        RECT 1390.4600 1479.7400 1392.0600 1480.2200 ;
        RECT 1345.4600 1485.1800 1347.0600 1485.6600 ;
        RECT 1345.4600 1490.6200 1347.0600 1491.1000 ;
        RECT 1345.4600 1468.8600 1347.0600 1469.3400 ;
        RECT 1345.4600 1474.3000 1347.0600 1474.7800 ;
        RECT 1345.4600 1479.7400 1347.0600 1480.2200 ;
        RECT 1390.4600 1457.9800 1392.0600 1458.4600 ;
        RECT 1390.4600 1463.4200 1392.0600 1463.9000 ;
        RECT 1390.4600 1441.6600 1392.0600 1442.1400 ;
        RECT 1390.4600 1447.1000 1392.0600 1447.5800 ;
        RECT 1390.4600 1452.5400 1392.0600 1453.0200 ;
        RECT 1345.4600 1457.9800 1347.0600 1458.4600 ;
        RECT 1345.4600 1463.4200 1347.0600 1463.9000 ;
        RECT 1345.4600 1441.6600 1347.0600 1442.1400 ;
        RECT 1345.4600 1447.1000 1347.0600 1447.5800 ;
        RECT 1345.4600 1452.5400 1347.0600 1453.0200 ;
        RECT 1300.4600 1485.1800 1302.0600 1485.6600 ;
        RECT 1300.4600 1490.6200 1302.0600 1491.1000 ;
        RECT 1293.3000 1485.1800 1294.9000 1485.6600 ;
        RECT 1293.3000 1490.6200 1294.9000 1491.1000 ;
        RECT 1300.4600 1468.8600 1302.0600 1469.3400 ;
        RECT 1300.4600 1474.3000 1302.0600 1474.7800 ;
        RECT 1300.4600 1479.7400 1302.0600 1480.2200 ;
        RECT 1293.3000 1468.8600 1294.9000 1469.3400 ;
        RECT 1293.3000 1474.3000 1294.9000 1474.7800 ;
        RECT 1293.3000 1479.7400 1294.9000 1480.2200 ;
        RECT 1300.4600 1457.9800 1302.0600 1458.4600 ;
        RECT 1300.4600 1463.4200 1302.0600 1463.9000 ;
        RECT 1293.3000 1457.9800 1294.9000 1458.4600 ;
        RECT 1293.3000 1463.4200 1294.9000 1463.9000 ;
        RECT 1300.4600 1441.6600 1302.0600 1442.1400 ;
        RECT 1300.4600 1447.1000 1302.0600 1447.5800 ;
        RECT 1300.4600 1452.5400 1302.0600 1453.0200 ;
        RECT 1293.3000 1441.6600 1294.9000 1442.1400 ;
        RECT 1293.3000 1447.1000 1294.9000 1447.5800 ;
        RECT 1293.3000 1452.5400 1294.9000 1453.0200 ;
        RECT 1293.3000 1496.0600 1294.9000 1496.5400 ;
        RECT 1300.4600 1496.0600 1302.0600 1496.5400 ;
        RECT 1345.4600 1496.0600 1347.0600 1496.5400 ;
        RECT 1390.4600 1496.0600 1392.0600 1496.5400 ;
        RECT 1496.0000 1430.7800 1497.6000 1431.2600 ;
        RECT 1496.0000 1436.2200 1497.6000 1436.7000 ;
        RECT 1480.4600 1430.7800 1482.0600 1431.2600 ;
        RECT 1480.4600 1436.2200 1482.0600 1436.7000 ;
        RECT 1496.0000 1414.4600 1497.6000 1414.9400 ;
        RECT 1496.0000 1419.9000 1497.6000 1420.3800 ;
        RECT 1496.0000 1425.3400 1497.6000 1425.8200 ;
        RECT 1480.4600 1414.4600 1482.0600 1414.9400 ;
        RECT 1480.4600 1419.9000 1482.0600 1420.3800 ;
        RECT 1480.4600 1425.3400 1482.0600 1425.8200 ;
        RECT 1496.0000 1403.5800 1497.6000 1404.0600 ;
        RECT 1496.0000 1409.0200 1497.6000 1409.5000 ;
        RECT 1480.4600 1403.5800 1482.0600 1404.0600 ;
        RECT 1480.4600 1409.0200 1482.0600 1409.5000 ;
        RECT 1496.0000 1387.2600 1497.6000 1387.7400 ;
        RECT 1496.0000 1392.7000 1497.6000 1393.1800 ;
        RECT 1496.0000 1398.1400 1497.6000 1398.6200 ;
        RECT 1480.4600 1387.2600 1482.0600 1387.7400 ;
        RECT 1480.4600 1392.7000 1482.0600 1393.1800 ;
        RECT 1480.4600 1398.1400 1482.0600 1398.6200 ;
        RECT 1435.4600 1430.7800 1437.0600 1431.2600 ;
        RECT 1435.4600 1436.2200 1437.0600 1436.7000 ;
        RECT 1435.4600 1414.4600 1437.0600 1414.9400 ;
        RECT 1435.4600 1419.9000 1437.0600 1420.3800 ;
        RECT 1435.4600 1425.3400 1437.0600 1425.8200 ;
        RECT 1435.4600 1403.5800 1437.0600 1404.0600 ;
        RECT 1435.4600 1409.0200 1437.0600 1409.5000 ;
        RECT 1435.4600 1387.2600 1437.0600 1387.7400 ;
        RECT 1435.4600 1392.7000 1437.0600 1393.1800 ;
        RECT 1435.4600 1398.1400 1437.0600 1398.6200 ;
        RECT 1496.0000 1376.3800 1497.6000 1376.8600 ;
        RECT 1496.0000 1381.8200 1497.6000 1382.3000 ;
        RECT 1480.4600 1376.3800 1482.0600 1376.8600 ;
        RECT 1480.4600 1381.8200 1482.0600 1382.3000 ;
        RECT 1496.0000 1360.0600 1497.6000 1360.5400 ;
        RECT 1496.0000 1365.5000 1497.6000 1365.9800 ;
        RECT 1496.0000 1370.9400 1497.6000 1371.4200 ;
        RECT 1480.4600 1360.0600 1482.0600 1360.5400 ;
        RECT 1480.4600 1365.5000 1482.0600 1365.9800 ;
        RECT 1480.4600 1370.9400 1482.0600 1371.4200 ;
        RECT 1496.0000 1349.1800 1497.6000 1349.6600 ;
        RECT 1496.0000 1354.6200 1497.6000 1355.1000 ;
        RECT 1480.4600 1349.1800 1482.0600 1349.6600 ;
        RECT 1480.4600 1354.6200 1482.0600 1355.1000 ;
        RECT 1480.4600 1343.7400 1482.0600 1344.2200 ;
        RECT 1496.0000 1343.7400 1497.6000 1344.2200 ;
        RECT 1435.4600 1376.3800 1437.0600 1376.8600 ;
        RECT 1435.4600 1381.8200 1437.0600 1382.3000 ;
        RECT 1435.4600 1360.0600 1437.0600 1360.5400 ;
        RECT 1435.4600 1365.5000 1437.0600 1365.9800 ;
        RECT 1435.4600 1370.9400 1437.0600 1371.4200 ;
        RECT 1435.4600 1349.1800 1437.0600 1349.6600 ;
        RECT 1435.4600 1354.6200 1437.0600 1355.1000 ;
        RECT 1435.4600 1343.7400 1437.0600 1344.2200 ;
        RECT 1390.4600 1430.7800 1392.0600 1431.2600 ;
        RECT 1390.4600 1436.2200 1392.0600 1436.7000 ;
        RECT 1390.4600 1414.4600 1392.0600 1414.9400 ;
        RECT 1390.4600 1419.9000 1392.0600 1420.3800 ;
        RECT 1390.4600 1425.3400 1392.0600 1425.8200 ;
        RECT 1345.4600 1430.7800 1347.0600 1431.2600 ;
        RECT 1345.4600 1436.2200 1347.0600 1436.7000 ;
        RECT 1345.4600 1414.4600 1347.0600 1414.9400 ;
        RECT 1345.4600 1419.9000 1347.0600 1420.3800 ;
        RECT 1345.4600 1425.3400 1347.0600 1425.8200 ;
        RECT 1390.4600 1403.5800 1392.0600 1404.0600 ;
        RECT 1390.4600 1409.0200 1392.0600 1409.5000 ;
        RECT 1390.4600 1387.2600 1392.0600 1387.7400 ;
        RECT 1390.4600 1392.7000 1392.0600 1393.1800 ;
        RECT 1390.4600 1398.1400 1392.0600 1398.6200 ;
        RECT 1345.4600 1403.5800 1347.0600 1404.0600 ;
        RECT 1345.4600 1409.0200 1347.0600 1409.5000 ;
        RECT 1345.4600 1387.2600 1347.0600 1387.7400 ;
        RECT 1345.4600 1392.7000 1347.0600 1393.1800 ;
        RECT 1345.4600 1398.1400 1347.0600 1398.6200 ;
        RECT 1300.4600 1430.7800 1302.0600 1431.2600 ;
        RECT 1300.4600 1436.2200 1302.0600 1436.7000 ;
        RECT 1293.3000 1430.7800 1294.9000 1431.2600 ;
        RECT 1293.3000 1436.2200 1294.9000 1436.7000 ;
        RECT 1300.4600 1414.4600 1302.0600 1414.9400 ;
        RECT 1300.4600 1419.9000 1302.0600 1420.3800 ;
        RECT 1300.4600 1425.3400 1302.0600 1425.8200 ;
        RECT 1293.3000 1414.4600 1294.9000 1414.9400 ;
        RECT 1293.3000 1419.9000 1294.9000 1420.3800 ;
        RECT 1293.3000 1425.3400 1294.9000 1425.8200 ;
        RECT 1300.4600 1403.5800 1302.0600 1404.0600 ;
        RECT 1300.4600 1409.0200 1302.0600 1409.5000 ;
        RECT 1293.3000 1403.5800 1294.9000 1404.0600 ;
        RECT 1293.3000 1409.0200 1294.9000 1409.5000 ;
        RECT 1300.4600 1387.2600 1302.0600 1387.7400 ;
        RECT 1300.4600 1392.7000 1302.0600 1393.1800 ;
        RECT 1300.4600 1398.1400 1302.0600 1398.6200 ;
        RECT 1293.3000 1387.2600 1294.9000 1387.7400 ;
        RECT 1293.3000 1392.7000 1294.9000 1393.1800 ;
        RECT 1293.3000 1398.1400 1294.9000 1398.6200 ;
        RECT 1390.4600 1376.3800 1392.0600 1376.8600 ;
        RECT 1390.4600 1381.8200 1392.0600 1382.3000 ;
        RECT 1390.4600 1360.0600 1392.0600 1360.5400 ;
        RECT 1390.4600 1365.5000 1392.0600 1365.9800 ;
        RECT 1390.4600 1370.9400 1392.0600 1371.4200 ;
        RECT 1345.4600 1376.3800 1347.0600 1376.8600 ;
        RECT 1345.4600 1381.8200 1347.0600 1382.3000 ;
        RECT 1345.4600 1360.0600 1347.0600 1360.5400 ;
        RECT 1345.4600 1365.5000 1347.0600 1365.9800 ;
        RECT 1345.4600 1370.9400 1347.0600 1371.4200 ;
        RECT 1390.4600 1354.6200 1392.0600 1355.1000 ;
        RECT 1390.4600 1349.1800 1392.0600 1349.6600 ;
        RECT 1390.4600 1343.7400 1392.0600 1344.2200 ;
        RECT 1345.4600 1354.6200 1347.0600 1355.1000 ;
        RECT 1345.4600 1349.1800 1347.0600 1349.6600 ;
        RECT 1345.4600 1343.7400 1347.0600 1344.2200 ;
        RECT 1300.4600 1376.3800 1302.0600 1376.8600 ;
        RECT 1300.4600 1381.8200 1302.0600 1382.3000 ;
        RECT 1293.3000 1376.3800 1294.9000 1376.8600 ;
        RECT 1293.3000 1381.8200 1294.9000 1382.3000 ;
        RECT 1300.4600 1360.0600 1302.0600 1360.5400 ;
        RECT 1300.4600 1365.5000 1302.0600 1365.9800 ;
        RECT 1300.4600 1370.9400 1302.0600 1371.4200 ;
        RECT 1293.3000 1360.0600 1294.9000 1360.5400 ;
        RECT 1293.3000 1365.5000 1294.9000 1365.9800 ;
        RECT 1293.3000 1370.9400 1294.9000 1371.4200 ;
        RECT 1300.4600 1349.1800 1302.0600 1349.6600 ;
        RECT 1300.4600 1354.6200 1302.0600 1355.1000 ;
        RECT 1293.3000 1349.1800 1294.9000 1349.6600 ;
        RECT 1293.3000 1354.6200 1294.9000 1355.1000 ;
        RECT 1293.3000 1343.7400 1294.9000 1344.2200 ;
        RECT 1300.4600 1343.7400 1302.0600 1344.2200 ;
        RECT 1290.3400 1545.9300 1500.5600 1547.5300 ;
        RECT 1290.3400 1334.2300 1500.5600 1335.8300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1331.4000 1294.9000 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1549.4400 1294.9000 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1331.4000 1497.6000 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1549.4400 1497.6000 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1334.2300 1291.9400 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1334.2300 1500.5600 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1545.9300 1291.9400 1547.5300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1545.9300 1500.5600 1547.5300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 1104.5900 1482.0600 1317.8900 ;
        RECT 1435.4600 1104.5900 1437.0600 1317.8900 ;
        RECT 1390.4600 1104.5900 1392.0600 1317.8900 ;
        RECT 1345.4600 1104.5900 1347.0600 1317.8900 ;
        RECT 1300.4600 1104.5900 1302.0600 1317.8900 ;
        RECT 1496.0000 1101.7600 1497.6000 1321.4000 ;
        RECT 1293.3000 1101.7600 1294.9000 1321.4000 ;
      LAYER met3 ;
        RECT 1480.4600 1309.9400 1482.0600 1310.4200 ;
        RECT 1496.0000 1309.9400 1497.6000 1310.4200 ;
        RECT 1496.0000 1299.0600 1497.6000 1299.5400 ;
        RECT 1496.0000 1304.5000 1497.6000 1304.9800 ;
        RECT 1480.4600 1299.0600 1482.0600 1299.5400 ;
        RECT 1480.4600 1304.5000 1482.0600 1304.9800 ;
        RECT 1496.0000 1282.7400 1497.6000 1283.2200 ;
        RECT 1496.0000 1288.1800 1497.6000 1288.6600 ;
        RECT 1480.4600 1282.7400 1482.0600 1283.2200 ;
        RECT 1480.4600 1288.1800 1482.0600 1288.6600 ;
        RECT 1496.0000 1271.8600 1497.6000 1272.3400 ;
        RECT 1496.0000 1277.3000 1497.6000 1277.7800 ;
        RECT 1480.4600 1271.8600 1482.0600 1272.3400 ;
        RECT 1480.4600 1277.3000 1482.0600 1277.7800 ;
        RECT 1480.4600 1293.6200 1482.0600 1294.1000 ;
        RECT 1496.0000 1293.6200 1497.6000 1294.1000 ;
        RECT 1435.4600 1299.0600 1437.0600 1299.5400 ;
        RECT 1435.4600 1304.5000 1437.0600 1304.9800 ;
        RECT 1435.4600 1309.9400 1437.0600 1310.4200 ;
        RECT 1435.4600 1282.7400 1437.0600 1283.2200 ;
        RECT 1435.4600 1288.1800 1437.0600 1288.6600 ;
        RECT 1435.4600 1277.3000 1437.0600 1277.7800 ;
        RECT 1435.4600 1271.8600 1437.0600 1272.3400 ;
        RECT 1435.4600 1293.6200 1437.0600 1294.1000 ;
        RECT 1496.0000 1255.5400 1497.6000 1256.0200 ;
        RECT 1496.0000 1260.9800 1497.6000 1261.4600 ;
        RECT 1480.4600 1255.5400 1482.0600 1256.0200 ;
        RECT 1480.4600 1260.9800 1482.0600 1261.4600 ;
        RECT 1496.0000 1239.2200 1497.6000 1239.7000 ;
        RECT 1496.0000 1244.6600 1497.6000 1245.1400 ;
        RECT 1496.0000 1250.1000 1497.6000 1250.5800 ;
        RECT 1480.4600 1239.2200 1482.0600 1239.7000 ;
        RECT 1480.4600 1244.6600 1482.0600 1245.1400 ;
        RECT 1480.4600 1250.1000 1482.0600 1250.5800 ;
        RECT 1496.0000 1228.3400 1497.6000 1228.8200 ;
        RECT 1496.0000 1233.7800 1497.6000 1234.2600 ;
        RECT 1480.4600 1228.3400 1482.0600 1228.8200 ;
        RECT 1480.4600 1233.7800 1482.0600 1234.2600 ;
        RECT 1496.0000 1212.0200 1497.6000 1212.5000 ;
        RECT 1496.0000 1217.4600 1497.6000 1217.9400 ;
        RECT 1496.0000 1222.9000 1497.6000 1223.3800 ;
        RECT 1480.4600 1212.0200 1482.0600 1212.5000 ;
        RECT 1480.4600 1217.4600 1482.0600 1217.9400 ;
        RECT 1480.4600 1222.9000 1482.0600 1223.3800 ;
        RECT 1435.4600 1255.5400 1437.0600 1256.0200 ;
        RECT 1435.4600 1260.9800 1437.0600 1261.4600 ;
        RECT 1435.4600 1239.2200 1437.0600 1239.7000 ;
        RECT 1435.4600 1244.6600 1437.0600 1245.1400 ;
        RECT 1435.4600 1250.1000 1437.0600 1250.5800 ;
        RECT 1435.4600 1228.3400 1437.0600 1228.8200 ;
        RECT 1435.4600 1233.7800 1437.0600 1234.2600 ;
        RECT 1435.4600 1212.0200 1437.0600 1212.5000 ;
        RECT 1435.4600 1217.4600 1437.0600 1217.9400 ;
        RECT 1435.4600 1222.9000 1437.0600 1223.3800 ;
        RECT 1435.4600 1266.4200 1437.0600 1266.9000 ;
        RECT 1480.4600 1266.4200 1482.0600 1266.9000 ;
        RECT 1496.0000 1266.4200 1497.6000 1266.9000 ;
        RECT 1390.4600 1299.0600 1392.0600 1299.5400 ;
        RECT 1390.4600 1304.5000 1392.0600 1304.9800 ;
        RECT 1390.4600 1309.9400 1392.0600 1310.4200 ;
        RECT 1345.4600 1299.0600 1347.0600 1299.5400 ;
        RECT 1345.4600 1304.5000 1347.0600 1304.9800 ;
        RECT 1345.4600 1309.9400 1347.0600 1310.4200 ;
        RECT 1390.4600 1282.7400 1392.0600 1283.2200 ;
        RECT 1390.4600 1288.1800 1392.0600 1288.6600 ;
        RECT 1390.4600 1271.8600 1392.0600 1272.3400 ;
        RECT 1390.4600 1277.3000 1392.0600 1277.7800 ;
        RECT 1345.4600 1282.7400 1347.0600 1283.2200 ;
        RECT 1345.4600 1288.1800 1347.0600 1288.6600 ;
        RECT 1345.4600 1271.8600 1347.0600 1272.3400 ;
        RECT 1345.4600 1277.3000 1347.0600 1277.7800 ;
        RECT 1345.4600 1293.6200 1347.0600 1294.1000 ;
        RECT 1390.4600 1293.6200 1392.0600 1294.1000 ;
        RECT 1293.3000 1309.9400 1294.9000 1310.4200 ;
        RECT 1300.4600 1309.9400 1302.0600 1310.4200 ;
        RECT 1300.4600 1299.0600 1302.0600 1299.5400 ;
        RECT 1300.4600 1304.5000 1302.0600 1304.9800 ;
        RECT 1293.3000 1299.0600 1294.9000 1299.5400 ;
        RECT 1293.3000 1304.5000 1294.9000 1304.9800 ;
        RECT 1300.4600 1282.7400 1302.0600 1283.2200 ;
        RECT 1300.4600 1288.1800 1302.0600 1288.6600 ;
        RECT 1293.3000 1282.7400 1294.9000 1283.2200 ;
        RECT 1293.3000 1288.1800 1294.9000 1288.6600 ;
        RECT 1300.4600 1271.8600 1302.0600 1272.3400 ;
        RECT 1300.4600 1277.3000 1302.0600 1277.7800 ;
        RECT 1293.3000 1271.8600 1294.9000 1272.3400 ;
        RECT 1293.3000 1277.3000 1294.9000 1277.7800 ;
        RECT 1293.3000 1293.6200 1294.9000 1294.1000 ;
        RECT 1300.4600 1293.6200 1302.0600 1294.1000 ;
        RECT 1390.4600 1255.5400 1392.0600 1256.0200 ;
        RECT 1390.4600 1260.9800 1392.0600 1261.4600 ;
        RECT 1390.4600 1239.2200 1392.0600 1239.7000 ;
        RECT 1390.4600 1244.6600 1392.0600 1245.1400 ;
        RECT 1390.4600 1250.1000 1392.0600 1250.5800 ;
        RECT 1345.4600 1255.5400 1347.0600 1256.0200 ;
        RECT 1345.4600 1260.9800 1347.0600 1261.4600 ;
        RECT 1345.4600 1239.2200 1347.0600 1239.7000 ;
        RECT 1345.4600 1244.6600 1347.0600 1245.1400 ;
        RECT 1345.4600 1250.1000 1347.0600 1250.5800 ;
        RECT 1390.4600 1228.3400 1392.0600 1228.8200 ;
        RECT 1390.4600 1233.7800 1392.0600 1234.2600 ;
        RECT 1390.4600 1212.0200 1392.0600 1212.5000 ;
        RECT 1390.4600 1217.4600 1392.0600 1217.9400 ;
        RECT 1390.4600 1222.9000 1392.0600 1223.3800 ;
        RECT 1345.4600 1228.3400 1347.0600 1228.8200 ;
        RECT 1345.4600 1233.7800 1347.0600 1234.2600 ;
        RECT 1345.4600 1212.0200 1347.0600 1212.5000 ;
        RECT 1345.4600 1217.4600 1347.0600 1217.9400 ;
        RECT 1345.4600 1222.9000 1347.0600 1223.3800 ;
        RECT 1300.4600 1255.5400 1302.0600 1256.0200 ;
        RECT 1300.4600 1260.9800 1302.0600 1261.4600 ;
        RECT 1293.3000 1255.5400 1294.9000 1256.0200 ;
        RECT 1293.3000 1260.9800 1294.9000 1261.4600 ;
        RECT 1300.4600 1239.2200 1302.0600 1239.7000 ;
        RECT 1300.4600 1244.6600 1302.0600 1245.1400 ;
        RECT 1300.4600 1250.1000 1302.0600 1250.5800 ;
        RECT 1293.3000 1239.2200 1294.9000 1239.7000 ;
        RECT 1293.3000 1244.6600 1294.9000 1245.1400 ;
        RECT 1293.3000 1250.1000 1294.9000 1250.5800 ;
        RECT 1300.4600 1228.3400 1302.0600 1228.8200 ;
        RECT 1300.4600 1233.7800 1302.0600 1234.2600 ;
        RECT 1293.3000 1228.3400 1294.9000 1228.8200 ;
        RECT 1293.3000 1233.7800 1294.9000 1234.2600 ;
        RECT 1300.4600 1212.0200 1302.0600 1212.5000 ;
        RECT 1300.4600 1217.4600 1302.0600 1217.9400 ;
        RECT 1300.4600 1222.9000 1302.0600 1223.3800 ;
        RECT 1293.3000 1212.0200 1294.9000 1212.5000 ;
        RECT 1293.3000 1217.4600 1294.9000 1217.9400 ;
        RECT 1293.3000 1222.9000 1294.9000 1223.3800 ;
        RECT 1293.3000 1266.4200 1294.9000 1266.9000 ;
        RECT 1300.4600 1266.4200 1302.0600 1266.9000 ;
        RECT 1345.4600 1266.4200 1347.0600 1266.9000 ;
        RECT 1390.4600 1266.4200 1392.0600 1266.9000 ;
        RECT 1496.0000 1201.1400 1497.6000 1201.6200 ;
        RECT 1496.0000 1206.5800 1497.6000 1207.0600 ;
        RECT 1480.4600 1201.1400 1482.0600 1201.6200 ;
        RECT 1480.4600 1206.5800 1482.0600 1207.0600 ;
        RECT 1496.0000 1184.8200 1497.6000 1185.3000 ;
        RECT 1496.0000 1190.2600 1497.6000 1190.7400 ;
        RECT 1496.0000 1195.7000 1497.6000 1196.1800 ;
        RECT 1480.4600 1184.8200 1482.0600 1185.3000 ;
        RECT 1480.4600 1190.2600 1482.0600 1190.7400 ;
        RECT 1480.4600 1195.7000 1482.0600 1196.1800 ;
        RECT 1496.0000 1173.9400 1497.6000 1174.4200 ;
        RECT 1496.0000 1179.3800 1497.6000 1179.8600 ;
        RECT 1480.4600 1173.9400 1482.0600 1174.4200 ;
        RECT 1480.4600 1179.3800 1482.0600 1179.8600 ;
        RECT 1496.0000 1157.6200 1497.6000 1158.1000 ;
        RECT 1496.0000 1163.0600 1497.6000 1163.5400 ;
        RECT 1496.0000 1168.5000 1497.6000 1168.9800 ;
        RECT 1480.4600 1157.6200 1482.0600 1158.1000 ;
        RECT 1480.4600 1163.0600 1482.0600 1163.5400 ;
        RECT 1480.4600 1168.5000 1482.0600 1168.9800 ;
        RECT 1435.4600 1201.1400 1437.0600 1201.6200 ;
        RECT 1435.4600 1206.5800 1437.0600 1207.0600 ;
        RECT 1435.4600 1184.8200 1437.0600 1185.3000 ;
        RECT 1435.4600 1190.2600 1437.0600 1190.7400 ;
        RECT 1435.4600 1195.7000 1437.0600 1196.1800 ;
        RECT 1435.4600 1173.9400 1437.0600 1174.4200 ;
        RECT 1435.4600 1179.3800 1437.0600 1179.8600 ;
        RECT 1435.4600 1157.6200 1437.0600 1158.1000 ;
        RECT 1435.4600 1163.0600 1437.0600 1163.5400 ;
        RECT 1435.4600 1168.5000 1437.0600 1168.9800 ;
        RECT 1496.0000 1146.7400 1497.6000 1147.2200 ;
        RECT 1496.0000 1152.1800 1497.6000 1152.6600 ;
        RECT 1480.4600 1146.7400 1482.0600 1147.2200 ;
        RECT 1480.4600 1152.1800 1482.0600 1152.6600 ;
        RECT 1496.0000 1130.4200 1497.6000 1130.9000 ;
        RECT 1496.0000 1135.8600 1497.6000 1136.3400 ;
        RECT 1496.0000 1141.3000 1497.6000 1141.7800 ;
        RECT 1480.4600 1130.4200 1482.0600 1130.9000 ;
        RECT 1480.4600 1135.8600 1482.0600 1136.3400 ;
        RECT 1480.4600 1141.3000 1482.0600 1141.7800 ;
        RECT 1496.0000 1119.5400 1497.6000 1120.0200 ;
        RECT 1496.0000 1124.9800 1497.6000 1125.4600 ;
        RECT 1480.4600 1119.5400 1482.0600 1120.0200 ;
        RECT 1480.4600 1124.9800 1482.0600 1125.4600 ;
        RECT 1480.4600 1114.1000 1482.0600 1114.5800 ;
        RECT 1496.0000 1114.1000 1497.6000 1114.5800 ;
        RECT 1435.4600 1146.7400 1437.0600 1147.2200 ;
        RECT 1435.4600 1152.1800 1437.0600 1152.6600 ;
        RECT 1435.4600 1130.4200 1437.0600 1130.9000 ;
        RECT 1435.4600 1135.8600 1437.0600 1136.3400 ;
        RECT 1435.4600 1141.3000 1437.0600 1141.7800 ;
        RECT 1435.4600 1119.5400 1437.0600 1120.0200 ;
        RECT 1435.4600 1124.9800 1437.0600 1125.4600 ;
        RECT 1435.4600 1114.1000 1437.0600 1114.5800 ;
        RECT 1390.4600 1201.1400 1392.0600 1201.6200 ;
        RECT 1390.4600 1206.5800 1392.0600 1207.0600 ;
        RECT 1390.4600 1184.8200 1392.0600 1185.3000 ;
        RECT 1390.4600 1190.2600 1392.0600 1190.7400 ;
        RECT 1390.4600 1195.7000 1392.0600 1196.1800 ;
        RECT 1345.4600 1201.1400 1347.0600 1201.6200 ;
        RECT 1345.4600 1206.5800 1347.0600 1207.0600 ;
        RECT 1345.4600 1184.8200 1347.0600 1185.3000 ;
        RECT 1345.4600 1190.2600 1347.0600 1190.7400 ;
        RECT 1345.4600 1195.7000 1347.0600 1196.1800 ;
        RECT 1390.4600 1173.9400 1392.0600 1174.4200 ;
        RECT 1390.4600 1179.3800 1392.0600 1179.8600 ;
        RECT 1390.4600 1157.6200 1392.0600 1158.1000 ;
        RECT 1390.4600 1163.0600 1392.0600 1163.5400 ;
        RECT 1390.4600 1168.5000 1392.0600 1168.9800 ;
        RECT 1345.4600 1173.9400 1347.0600 1174.4200 ;
        RECT 1345.4600 1179.3800 1347.0600 1179.8600 ;
        RECT 1345.4600 1157.6200 1347.0600 1158.1000 ;
        RECT 1345.4600 1163.0600 1347.0600 1163.5400 ;
        RECT 1345.4600 1168.5000 1347.0600 1168.9800 ;
        RECT 1300.4600 1201.1400 1302.0600 1201.6200 ;
        RECT 1300.4600 1206.5800 1302.0600 1207.0600 ;
        RECT 1293.3000 1201.1400 1294.9000 1201.6200 ;
        RECT 1293.3000 1206.5800 1294.9000 1207.0600 ;
        RECT 1300.4600 1184.8200 1302.0600 1185.3000 ;
        RECT 1300.4600 1190.2600 1302.0600 1190.7400 ;
        RECT 1300.4600 1195.7000 1302.0600 1196.1800 ;
        RECT 1293.3000 1184.8200 1294.9000 1185.3000 ;
        RECT 1293.3000 1190.2600 1294.9000 1190.7400 ;
        RECT 1293.3000 1195.7000 1294.9000 1196.1800 ;
        RECT 1300.4600 1173.9400 1302.0600 1174.4200 ;
        RECT 1300.4600 1179.3800 1302.0600 1179.8600 ;
        RECT 1293.3000 1173.9400 1294.9000 1174.4200 ;
        RECT 1293.3000 1179.3800 1294.9000 1179.8600 ;
        RECT 1300.4600 1157.6200 1302.0600 1158.1000 ;
        RECT 1300.4600 1163.0600 1302.0600 1163.5400 ;
        RECT 1300.4600 1168.5000 1302.0600 1168.9800 ;
        RECT 1293.3000 1157.6200 1294.9000 1158.1000 ;
        RECT 1293.3000 1163.0600 1294.9000 1163.5400 ;
        RECT 1293.3000 1168.5000 1294.9000 1168.9800 ;
        RECT 1390.4600 1146.7400 1392.0600 1147.2200 ;
        RECT 1390.4600 1152.1800 1392.0600 1152.6600 ;
        RECT 1390.4600 1130.4200 1392.0600 1130.9000 ;
        RECT 1390.4600 1135.8600 1392.0600 1136.3400 ;
        RECT 1390.4600 1141.3000 1392.0600 1141.7800 ;
        RECT 1345.4600 1146.7400 1347.0600 1147.2200 ;
        RECT 1345.4600 1152.1800 1347.0600 1152.6600 ;
        RECT 1345.4600 1130.4200 1347.0600 1130.9000 ;
        RECT 1345.4600 1135.8600 1347.0600 1136.3400 ;
        RECT 1345.4600 1141.3000 1347.0600 1141.7800 ;
        RECT 1390.4600 1124.9800 1392.0600 1125.4600 ;
        RECT 1390.4600 1119.5400 1392.0600 1120.0200 ;
        RECT 1390.4600 1114.1000 1392.0600 1114.5800 ;
        RECT 1345.4600 1124.9800 1347.0600 1125.4600 ;
        RECT 1345.4600 1119.5400 1347.0600 1120.0200 ;
        RECT 1345.4600 1114.1000 1347.0600 1114.5800 ;
        RECT 1300.4600 1146.7400 1302.0600 1147.2200 ;
        RECT 1300.4600 1152.1800 1302.0600 1152.6600 ;
        RECT 1293.3000 1146.7400 1294.9000 1147.2200 ;
        RECT 1293.3000 1152.1800 1294.9000 1152.6600 ;
        RECT 1300.4600 1130.4200 1302.0600 1130.9000 ;
        RECT 1300.4600 1135.8600 1302.0600 1136.3400 ;
        RECT 1300.4600 1141.3000 1302.0600 1141.7800 ;
        RECT 1293.3000 1130.4200 1294.9000 1130.9000 ;
        RECT 1293.3000 1135.8600 1294.9000 1136.3400 ;
        RECT 1293.3000 1141.3000 1294.9000 1141.7800 ;
        RECT 1300.4600 1119.5400 1302.0600 1120.0200 ;
        RECT 1300.4600 1124.9800 1302.0600 1125.4600 ;
        RECT 1293.3000 1119.5400 1294.9000 1120.0200 ;
        RECT 1293.3000 1124.9800 1294.9000 1125.4600 ;
        RECT 1293.3000 1114.1000 1294.9000 1114.5800 ;
        RECT 1300.4600 1114.1000 1302.0600 1114.5800 ;
        RECT 1290.3400 1316.2900 1500.5600 1317.8900 ;
        RECT 1290.3400 1104.5900 1500.5600 1106.1900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1101.7600 1294.9000 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1319.8000 1294.9000 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1101.7600 1497.6000 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1319.8000 1497.6000 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1104.5900 1291.9400 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1104.5900 1500.5600 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1316.2900 1291.9400 1317.8900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1316.2900 1500.5600 1317.8900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 874.9500 1482.0600 1088.2500 ;
        RECT 1435.4600 874.9500 1437.0600 1088.2500 ;
        RECT 1390.4600 874.9500 1392.0600 1088.2500 ;
        RECT 1345.4600 874.9500 1347.0600 1088.2500 ;
        RECT 1300.4600 874.9500 1302.0600 1088.2500 ;
        RECT 1496.0000 872.1200 1497.6000 1091.7600 ;
        RECT 1293.3000 872.1200 1294.9000 1091.7600 ;
      LAYER met3 ;
        RECT 1480.4600 1080.3000 1482.0600 1080.7800 ;
        RECT 1496.0000 1080.3000 1497.6000 1080.7800 ;
        RECT 1496.0000 1069.4200 1497.6000 1069.9000 ;
        RECT 1496.0000 1074.8600 1497.6000 1075.3400 ;
        RECT 1480.4600 1069.4200 1482.0600 1069.9000 ;
        RECT 1480.4600 1074.8600 1482.0600 1075.3400 ;
        RECT 1496.0000 1053.1000 1497.6000 1053.5800 ;
        RECT 1496.0000 1058.5400 1497.6000 1059.0200 ;
        RECT 1480.4600 1053.1000 1482.0600 1053.5800 ;
        RECT 1480.4600 1058.5400 1482.0600 1059.0200 ;
        RECT 1496.0000 1042.2200 1497.6000 1042.7000 ;
        RECT 1496.0000 1047.6600 1497.6000 1048.1400 ;
        RECT 1480.4600 1042.2200 1482.0600 1042.7000 ;
        RECT 1480.4600 1047.6600 1482.0600 1048.1400 ;
        RECT 1480.4600 1063.9800 1482.0600 1064.4600 ;
        RECT 1496.0000 1063.9800 1497.6000 1064.4600 ;
        RECT 1435.4600 1069.4200 1437.0600 1069.9000 ;
        RECT 1435.4600 1074.8600 1437.0600 1075.3400 ;
        RECT 1435.4600 1080.3000 1437.0600 1080.7800 ;
        RECT 1435.4600 1053.1000 1437.0600 1053.5800 ;
        RECT 1435.4600 1058.5400 1437.0600 1059.0200 ;
        RECT 1435.4600 1047.6600 1437.0600 1048.1400 ;
        RECT 1435.4600 1042.2200 1437.0600 1042.7000 ;
        RECT 1435.4600 1063.9800 1437.0600 1064.4600 ;
        RECT 1496.0000 1025.9000 1497.6000 1026.3800 ;
        RECT 1496.0000 1031.3400 1497.6000 1031.8200 ;
        RECT 1480.4600 1025.9000 1482.0600 1026.3800 ;
        RECT 1480.4600 1031.3400 1482.0600 1031.8200 ;
        RECT 1496.0000 1009.5800 1497.6000 1010.0600 ;
        RECT 1496.0000 1015.0200 1497.6000 1015.5000 ;
        RECT 1496.0000 1020.4600 1497.6000 1020.9400 ;
        RECT 1480.4600 1009.5800 1482.0600 1010.0600 ;
        RECT 1480.4600 1015.0200 1482.0600 1015.5000 ;
        RECT 1480.4600 1020.4600 1482.0600 1020.9400 ;
        RECT 1496.0000 998.7000 1497.6000 999.1800 ;
        RECT 1496.0000 1004.1400 1497.6000 1004.6200 ;
        RECT 1480.4600 998.7000 1482.0600 999.1800 ;
        RECT 1480.4600 1004.1400 1482.0600 1004.6200 ;
        RECT 1496.0000 982.3800 1497.6000 982.8600 ;
        RECT 1496.0000 987.8200 1497.6000 988.3000 ;
        RECT 1496.0000 993.2600 1497.6000 993.7400 ;
        RECT 1480.4600 982.3800 1482.0600 982.8600 ;
        RECT 1480.4600 987.8200 1482.0600 988.3000 ;
        RECT 1480.4600 993.2600 1482.0600 993.7400 ;
        RECT 1435.4600 1025.9000 1437.0600 1026.3800 ;
        RECT 1435.4600 1031.3400 1437.0600 1031.8200 ;
        RECT 1435.4600 1009.5800 1437.0600 1010.0600 ;
        RECT 1435.4600 1015.0200 1437.0600 1015.5000 ;
        RECT 1435.4600 1020.4600 1437.0600 1020.9400 ;
        RECT 1435.4600 998.7000 1437.0600 999.1800 ;
        RECT 1435.4600 1004.1400 1437.0600 1004.6200 ;
        RECT 1435.4600 982.3800 1437.0600 982.8600 ;
        RECT 1435.4600 987.8200 1437.0600 988.3000 ;
        RECT 1435.4600 993.2600 1437.0600 993.7400 ;
        RECT 1435.4600 1036.7800 1437.0600 1037.2600 ;
        RECT 1480.4600 1036.7800 1482.0600 1037.2600 ;
        RECT 1496.0000 1036.7800 1497.6000 1037.2600 ;
        RECT 1390.4600 1069.4200 1392.0600 1069.9000 ;
        RECT 1390.4600 1074.8600 1392.0600 1075.3400 ;
        RECT 1390.4600 1080.3000 1392.0600 1080.7800 ;
        RECT 1345.4600 1069.4200 1347.0600 1069.9000 ;
        RECT 1345.4600 1074.8600 1347.0600 1075.3400 ;
        RECT 1345.4600 1080.3000 1347.0600 1080.7800 ;
        RECT 1390.4600 1053.1000 1392.0600 1053.5800 ;
        RECT 1390.4600 1058.5400 1392.0600 1059.0200 ;
        RECT 1390.4600 1042.2200 1392.0600 1042.7000 ;
        RECT 1390.4600 1047.6600 1392.0600 1048.1400 ;
        RECT 1345.4600 1053.1000 1347.0600 1053.5800 ;
        RECT 1345.4600 1058.5400 1347.0600 1059.0200 ;
        RECT 1345.4600 1042.2200 1347.0600 1042.7000 ;
        RECT 1345.4600 1047.6600 1347.0600 1048.1400 ;
        RECT 1345.4600 1063.9800 1347.0600 1064.4600 ;
        RECT 1390.4600 1063.9800 1392.0600 1064.4600 ;
        RECT 1293.3000 1080.3000 1294.9000 1080.7800 ;
        RECT 1300.4600 1080.3000 1302.0600 1080.7800 ;
        RECT 1300.4600 1069.4200 1302.0600 1069.9000 ;
        RECT 1300.4600 1074.8600 1302.0600 1075.3400 ;
        RECT 1293.3000 1069.4200 1294.9000 1069.9000 ;
        RECT 1293.3000 1074.8600 1294.9000 1075.3400 ;
        RECT 1300.4600 1053.1000 1302.0600 1053.5800 ;
        RECT 1300.4600 1058.5400 1302.0600 1059.0200 ;
        RECT 1293.3000 1053.1000 1294.9000 1053.5800 ;
        RECT 1293.3000 1058.5400 1294.9000 1059.0200 ;
        RECT 1300.4600 1042.2200 1302.0600 1042.7000 ;
        RECT 1300.4600 1047.6600 1302.0600 1048.1400 ;
        RECT 1293.3000 1042.2200 1294.9000 1042.7000 ;
        RECT 1293.3000 1047.6600 1294.9000 1048.1400 ;
        RECT 1293.3000 1063.9800 1294.9000 1064.4600 ;
        RECT 1300.4600 1063.9800 1302.0600 1064.4600 ;
        RECT 1390.4600 1025.9000 1392.0600 1026.3800 ;
        RECT 1390.4600 1031.3400 1392.0600 1031.8200 ;
        RECT 1390.4600 1009.5800 1392.0600 1010.0600 ;
        RECT 1390.4600 1015.0200 1392.0600 1015.5000 ;
        RECT 1390.4600 1020.4600 1392.0600 1020.9400 ;
        RECT 1345.4600 1025.9000 1347.0600 1026.3800 ;
        RECT 1345.4600 1031.3400 1347.0600 1031.8200 ;
        RECT 1345.4600 1009.5800 1347.0600 1010.0600 ;
        RECT 1345.4600 1015.0200 1347.0600 1015.5000 ;
        RECT 1345.4600 1020.4600 1347.0600 1020.9400 ;
        RECT 1390.4600 998.7000 1392.0600 999.1800 ;
        RECT 1390.4600 1004.1400 1392.0600 1004.6200 ;
        RECT 1390.4600 982.3800 1392.0600 982.8600 ;
        RECT 1390.4600 987.8200 1392.0600 988.3000 ;
        RECT 1390.4600 993.2600 1392.0600 993.7400 ;
        RECT 1345.4600 998.7000 1347.0600 999.1800 ;
        RECT 1345.4600 1004.1400 1347.0600 1004.6200 ;
        RECT 1345.4600 982.3800 1347.0600 982.8600 ;
        RECT 1345.4600 987.8200 1347.0600 988.3000 ;
        RECT 1345.4600 993.2600 1347.0600 993.7400 ;
        RECT 1300.4600 1025.9000 1302.0600 1026.3800 ;
        RECT 1300.4600 1031.3400 1302.0600 1031.8200 ;
        RECT 1293.3000 1025.9000 1294.9000 1026.3800 ;
        RECT 1293.3000 1031.3400 1294.9000 1031.8200 ;
        RECT 1300.4600 1009.5800 1302.0600 1010.0600 ;
        RECT 1300.4600 1015.0200 1302.0600 1015.5000 ;
        RECT 1300.4600 1020.4600 1302.0600 1020.9400 ;
        RECT 1293.3000 1009.5800 1294.9000 1010.0600 ;
        RECT 1293.3000 1015.0200 1294.9000 1015.5000 ;
        RECT 1293.3000 1020.4600 1294.9000 1020.9400 ;
        RECT 1300.4600 998.7000 1302.0600 999.1800 ;
        RECT 1300.4600 1004.1400 1302.0600 1004.6200 ;
        RECT 1293.3000 998.7000 1294.9000 999.1800 ;
        RECT 1293.3000 1004.1400 1294.9000 1004.6200 ;
        RECT 1300.4600 982.3800 1302.0600 982.8600 ;
        RECT 1300.4600 987.8200 1302.0600 988.3000 ;
        RECT 1300.4600 993.2600 1302.0600 993.7400 ;
        RECT 1293.3000 982.3800 1294.9000 982.8600 ;
        RECT 1293.3000 987.8200 1294.9000 988.3000 ;
        RECT 1293.3000 993.2600 1294.9000 993.7400 ;
        RECT 1293.3000 1036.7800 1294.9000 1037.2600 ;
        RECT 1300.4600 1036.7800 1302.0600 1037.2600 ;
        RECT 1345.4600 1036.7800 1347.0600 1037.2600 ;
        RECT 1390.4600 1036.7800 1392.0600 1037.2600 ;
        RECT 1496.0000 971.5000 1497.6000 971.9800 ;
        RECT 1496.0000 976.9400 1497.6000 977.4200 ;
        RECT 1480.4600 971.5000 1482.0600 971.9800 ;
        RECT 1480.4600 976.9400 1482.0600 977.4200 ;
        RECT 1496.0000 955.1800 1497.6000 955.6600 ;
        RECT 1496.0000 960.6200 1497.6000 961.1000 ;
        RECT 1496.0000 966.0600 1497.6000 966.5400 ;
        RECT 1480.4600 955.1800 1482.0600 955.6600 ;
        RECT 1480.4600 960.6200 1482.0600 961.1000 ;
        RECT 1480.4600 966.0600 1482.0600 966.5400 ;
        RECT 1496.0000 944.3000 1497.6000 944.7800 ;
        RECT 1496.0000 949.7400 1497.6000 950.2200 ;
        RECT 1480.4600 944.3000 1482.0600 944.7800 ;
        RECT 1480.4600 949.7400 1482.0600 950.2200 ;
        RECT 1496.0000 927.9800 1497.6000 928.4600 ;
        RECT 1496.0000 933.4200 1497.6000 933.9000 ;
        RECT 1496.0000 938.8600 1497.6000 939.3400 ;
        RECT 1480.4600 927.9800 1482.0600 928.4600 ;
        RECT 1480.4600 933.4200 1482.0600 933.9000 ;
        RECT 1480.4600 938.8600 1482.0600 939.3400 ;
        RECT 1435.4600 971.5000 1437.0600 971.9800 ;
        RECT 1435.4600 976.9400 1437.0600 977.4200 ;
        RECT 1435.4600 955.1800 1437.0600 955.6600 ;
        RECT 1435.4600 960.6200 1437.0600 961.1000 ;
        RECT 1435.4600 966.0600 1437.0600 966.5400 ;
        RECT 1435.4600 944.3000 1437.0600 944.7800 ;
        RECT 1435.4600 949.7400 1437.0600 950.2200 ;
        RECT 1435.4600 927.9800 1437.0600 928.4600 ;
        RECT 1435.4600 933.4200 1437.0600 933.9000 ;
        RECT 1435.4600 938.8600 1437.0600 939.3400 ;
        RECT 1496.0000 917.1000 1497.6000 917.5800 ;
        RECT 1496.0000 922.5400 1497.6000 923.0200 ;
        RECT 1480.4600 917.1000 1482.0600 917.5800 ;
        RECT 1480.4600 922.5400 1482.0600 923.0200 ;
        RECT 1496.0000 900.7800 1497.6000 901.2600 ;
        RECT 1496.0000 906.2200 1497.6000 906.7000 ;
        RECT 1496.0000 911.6600 1497.6000 912.1400 ;
        RECT 1480.4600 900.7800 1482.0600 901.2600 ;
        RECT 1480.4600 906.2200 1482.0600 906.7000 ;
        RECT 1480.4600 911.6600 1482.0600 912.1400 ;
        RECT 1496.0000 889.9000 1497.6000 890.3800 ;
        RECT 1496.0000 895.3400 1497.6000 895.8200 ;
        RECT 1480.4600 889.9000 1482.0600 890.3800 ;
        RECT 1480.4600 895.3400 1482.0600 895.8200 ;
        RECT 1480.4600 884.4600 1482.0600 884.9400 ;
        RECT 1496.0000 884.4600 1497.6000 884.9400 ;
        RECT 1435.4600 917.1000 1437.0600 917.5800 ;
        RECT 1435.4600 922.5400 1437.0600 923.0200 ;
        RECT 1435.4600 900.7800 1437.0600 901.2600 ;
        RECT 1435.4600 906.2200 1437.0600 906.7000 ;
        RECT 1435.4600 911.6600 1437.0600 912.1400 ;
        RECT 1435.4600 889.9000 1437.0600 890.3800 ;
        RECT 1435.4600 895.3400 1437.0600 895.8200 ;
        RECT 1435.4600 884.4600 1437.0600 884.9400 ;
        RECT 1390.4600 971.5000 1392.0600 971.9800 ;
        RECT 1390.4600 976.9400 1392.0600 977.4200 ;
        RECT 1390.4600 955.1800 1392.0600 955.6600 ;
        RECT 1390.4600 960.6200 1392.0600 961.1000 ;
        RECT 1390.4600 966.0600 1392.0600 966.5400 ;
        RECT 1345.4600 971.5000 1347.0600 971.9800 ;
        RECT 1345.4600 976.9400 1347.0600 977.4200 ;
        RECT 1345.4600 955.1800 1347.0600 955.6600 ;
        RECT 1345.4600 960.6200 1347.0600 961.1000 ;
        RECT 1345.4600 966.0600 1347.0600 966.5400 ;
        RECT 1390.4600 944.3000 1392.0600 944.7800 ;
        RECT 1390.4600 949.7400 1392.0600 950.2200 ;
        RECT 1390.4600 927.9800 1392.0600 928.4600 ;
        RECT 1390.4600 933.4200 1392.0600 933.9000 ;
        RECT 1390.4600 938.8600 1392.0600 939.3400 ;
        RECT 1345.4600 944.3000 1347.0600 944.7800 ;
        RECT 1345.4600 949.7400 1347.0600 950.2200 ;
        RECT 1345.4600 927.9800 1347.0600 928.4600 ;
        RECT 1345.4600 933.4200 1347.0600 933.9000 ;
        RECT 1345.4600 938.8600 1347.0600 939.3400 ;
        RECT 1300.4600 971.5000 1302.0600 971.9800 ;
        RECT 1300.4600 976.9400 1302.0600 977.4200 ;
        RECT 1293.3000 971.5000 1294.9000 971.9800 ;
        RECT 1293.3000 976.9400 1294.9000 977.4200 ;
        RECT 1300.4600 955.1800 1302.0600 955.6600 ;
        RECT 1300.4600 960.6200 1302.0600 961.1000 ;
        RECT 1300.4600 966.0600 1302.0600 966.5400 ;
        RECT 1293.3000 955.1800 1294.9000 955.6600 ;
        RECT 1293.3000 960.6200 1294.9000 961.1000 ;
        RECT 1293.3000 966.0600 1294.9000 966.5400 ;
        RECT 1300.4600 944.3000 1302.0600 944.7800 ;
        RECT 1300.4600 949.7400 1302.0600 950.2200 ;
        RECT 1293.3000 944.3000 1294.9000 944.7800 ;
        RECT 1293.3000 949.7400 1294.9000 950.2200 ;
        RECT 1300.4600 927.9800 1302.0600 928.4600 ;
        RECT 1300.4600 933.4200 1302.0600 933.9000 ;
        RECT 1300.4600 938.8600 1302.0600 939.3400 ;
        RECT 1293.3000 927.9800 1294.9000 928.4600 ;
        RECT 1293.3000 933.4200 1294.9000 933.9000 ;
        RECT 1293.3000 938.8600 1294.9000 939.3400 ;
        RECT 1390.4600 917.1000 1392.0600 917.5800 ;
        RECT 1390.4600 922.5400 1392.0600 923.0200 ;
        RECT 1390.4600 900.7800 1392.0600 901.2600 ;
        RECT 1390.4600 906.2200 1392.0600 906.7000 ;
        RECT 1390.4600 911.6600 1392.0600 912.1400 ;
        RECT 1345.4600 917.1000 1347.0600 917.5800 ;
        RECT 1345.4600 922.5400 1347.0600 923.0200 ;
        RECT 1345.4600 900.7800 1347.0600 901.2600 ;
        RECT 1345.4600 906.2200 1347.0600 906.7000 ;
        RECT 1345.4600 911.6600 1347.0600 912.1400 ;
        RECT 1390.4600 895.3400 1392.0600 895.8200 ;
        RECT 1390.4600 889.9000 1392.0600 890.3800 ;
        RECT 1390.4600 884.4600 1392.0600 884.9400 ;
        RECT 1345.4600 895.3400 1347.0600 895.8200 ;
        RECT 1345.4600 889.9000 1347.0600 890.3800 ;
        RECT 1345.4600 884.4600 1347.0600 884.9400 ;
        RECT 1300.4600 917.1000 1302.0600 917.5800 ;
        RECT 1300.4600 922.5400 1302.0600 923.0200 ;
        RECT 1293.3000 917.1000 1294.9000 917.5800 ;
        RECT 1293.3000 922.5400 1294.9000 923.0200 ;
        RECT 1300.4600 900.7800 1302.0600 901.2600 ;
        RECT 1300.4600 906.2200 1302.0600 906.7000 ;
        RECT 1300.4600 911.6600 1302.0600 912.1400 ;
        RECT 1293.3000 900.7800 1294.9000 901.2600 ;
        RECT 1293.3000 906.2200 1294.9000 906.7000 ;
        RECT 1293.3000 911.6600 1294.9000 912.1400 ;
        RECT 1300.4600 889.9000 1302.0600 890.3800 ;
        RECT 1300.4600 895.3400 1302.0600 895.8200 ;
        RECT 1293.3000 889.9000 1294.9000 890.3800 ;
        RECT 1293.3000 895.3400 1294.9000 895.8200 ;
        RECT 1293.3000 884.4600 1294.9000 884.9400 ;
        RECT 1300.4600 884.4600 1302.0600 884.9400 ;
        RECT 1290.3400 1086.6500 1500.5600 1088.2500 ;
        RECT 1290.3400 874.9500 1500.5600 876.5500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 872.1200 1294.9000 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 1090.1600 1294.9000 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 872.1200 1497.6000 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 1090.1600 1497.6000 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 874.9500 1291.9400 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 874.9500 1500.5600 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1086.6500 1291.9400 1088.2500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1086.6500 1500.5600 1088.2500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 645.3100 1482.0600 858.6100 ;
        RECT 1435.4600 645.3100 1437.0600 858.6100 ;
        RECT 1390.4600 645.3100 1392.0600 858.6100 ;
        RECT 1345.4600 645.3100 1347.0600 858.6100 ;
        RECT 1300.4600 645.3100 1302.0600 858.6100 ;
        RECT 1496.0000 642.4800 1497.6000 862.1200 ;
        RECT 1293.3000 642.4800 1294.9000 862.1200 ;
      LAYER met3 ;
        RECT 1480.4600 850.6600 1482.0600 851.1400 ;
        RECT 1496.0000 850.6600 1497.6000 851.1400 ;
        RECT 1496.0000 839.7800 1497.6000 840.2600 ;
        RECT 1496.0000 845.2200 1497.6000 845.7000 ;
        RECT 1480.4600 839.7800 1482.0600 840.2600 ;
        RECT 1480.4600 845.2200 1482.0600 845.7000 ;
        RECT 1496.0000 823.4600 1497.6000 823.9400 ;
        RECT 1496.0000 828.9000 1497.6000 829.3800 ;
        RECT 1480.4600 823.4600 1482.0600 823.9400 ;
        RECT 1480.4600 828.9000 1482.0600 829.3800 ;
        RECT 1496.0000 812.5800 1497.6000 813.0600 ;
        RECT 1496.0000 818.0200 1497.6000 818.5000 ;
        RECT 1480.4600 812.5800 1482.0600 813.0600 ;
        RECT 1480.4600 818.0200 1482.0600 818.5000 ;
        RECT 1480.4600 834.3400 1482.0600 834.8200 ;
        RECT 1496.0000 834.3400 1497.6000 834.8200 ;
        RECT 1435.4600 839.7800 1437.0600 840.2600 ;
        RECT 1435.4600 845.2200 1437.0600 845.7000 ;
        RECT 1435.4600 850.6600 1437.0600 851.1400 ;
        RECT 1435.4600 823.4600 1437.0600 823.9400 ;
        RECT 1435.4600 828.9000 1437.0600 829.3800 ;
        RECT 1435.4600 818.0200 1437.0600 818.5000 ;
        RECT 1435.4600 812.5800 1437.0600 813.0600 ;
        RECT 1435.4600 834.3400 1437.0600 834.8200 ;
        RECT 1496.0000 796.2600 1497.6000 796.7400 ;
        RECT 1496.0000 801.7000 1497.6000 802.1800 ;
        RECT 1480.4600 796.2600 1482.0600 796.7400 ;
        RECT 1480.4600 801.7000 1482.0600 802.1800 ;
        RECT 1496.0000 779.9400 1497.6000 780.4200 ;
        RECT 1496.0000 785.3800 1497.6000 785.8600 ;
        RECT 1496.0000 790.8200 1497.6000 791.3000 ;
        RECT 1480.4600 779.9400 1482.0600 780.4200 ;
        RECT 1480.4600 785.3800 1482.0600 785.8600 ;
        RECT 1480.4600 790.8200 1482.0600 791.3000 ;
        RECT 1496.0000 769.0600 1497.6000 769.5400 ;
        RECT 1496.0000 774.5000 1497.6000 774.9800 ;
        RECT 1480.4600 769.0600 1482.0600 769.5400 ;
        RECT 1480.4600 774.5000 1482.0600 774.9800 ;
        RECT 1496.0000 752.7400 1497.6000 753.2200 ;
        RECT 1496.0000 758.1800 1497.6000 758.6600 ;
        RECT 1496.0000 763.6200 1497.6000 764.1000 ;
        RECT 1480.4600 752.7400 1482.0600 753.2200 ;
        RECT 1480.4600 758.1800 1482.0600 758.6600 ;
        RECT 1480.4600 763.6200 1482.0600 764.1000 ;
        RECT 1435.4600 796.2600 1437.0600 796.7400 ;
        RECT 1435.4600 801.7000 1437.0600 802.1800 ;
        RECT 1435.4600 779.9400 1437.0600 780.4200 ;
        RECT 1435.4600 785.3800 1437.0600 785.8600 ;
        RECT 1435.4600 790.8200 1437.0600 791.3000 ;
        RECT 1435.4600 769.0600 1437.0600 769.5400 ;
        RECT 1435.4600 774.5000 1437.0600 774.9800 ;
        RECT 1435.4600 752.7400 1437.0600 753.2200 ;
        RECT 1435.4600 758.1800 1437.0600 758.6600 ;
        RECT 1435.4600 763.6200 1437.0600 764.1000 ;
        RECT 1435.4600 807.1400 1437.0600 807.6200 ;
        RECT 1480.4600 807.1400 1482.0600 807.6200 ;
        RECT 1496.0000 807.1400 1497.6000 807.6200 ;
        RECT 1390.4600 839.7800 1392.0600 840.2600 ;
        RECT 1390.4600 845.2200 1392.0600 845.7000 ;
        RECT 1390.4600 850.6600 1392.0600 851.1400 ;
        RECT 1345.4600 839.7800 1347.0600 840.2600 ;
        RECT 1345.4600 845.2200 1347.0600 845.7000 ;
        RECT 1345.4600 850.6600 1347.0600 851.1400 ;
        RECT 1390.4600 823.4600 1392.0600 823.9400 ;
        RECT 1390.4600 828.9000 1392.0600 829.3800 ;
        RECT 1390.4600 812.5800 1392.0600 813.0600 ;
        RECT 1390.4600 818.0200 1392.0600 818.5000 ;
        RECT 1345.4600 823.4600 1347.0600 823.9400 ;
        RECT 1345.4600 828.9000 1347.0600 829.3800 ;
        RECT 1345.4600 812.5800 1347.0600 813.0600 ;
        RECT 1345.4600 818.0200 1347.0600 818.5000 ;
        RECT 1345.4600 834.3400 1347.0600 834.8200 ;
        RECT 1390.4600 834.3400 1392.0600 834.8200 ;
        RECT 1293.3000 850.6600 1294.9000 851.1400 ;
        RECT 1300.4600 850.6600 1302.0600 851.1400 ;
        RECT 1300.4600 839.7800 1302.0600 840.2600 ;
        RECT 1300.4600 845.2200 1302.0600 845.7000 ;
        RECT 1293.3000 839.7800 1294.9000 840.2600 ;
        RECT 1293.3000 845.2200 1294.9000 845.7000 ;
        RECT 1300.4600 823.4600 1302.0600 823.9400 ;
        RECT 1300.4600 828.9000 1302.0600 829.3800 ;
        RECT 1293.3000 823.4600 1294.9000 823.9400 ;
        RECT 1293.3000 828.9000 1294.9000 829.3800 ;
        RECT 1300.4600 812.5800 1302.0600 813.0600 ;
        RECT 1300.4600 818.0200 1302.0600 818.5000 ;
        RECT 1293.3000 812.5800 1294.9000 813.0600 ;
        RECT 1293.3000 818.0200 1294.9000 818.5000 ;
        RECT 1293.3000 834.3400 1294.9000 834.8200 ;
        RECT 1300.4600 834.3400 1302.0600 834.8200 ;
        RECT 1390.4600 796.2600 1392.0600 796.7400 ;
        RECT 1390.4600 801.7000 1392.0600 802.1800 ;
        RECT 1390.4600 779.9400 1392.0600 780.4200 ;
        RECT 1390.4600 785.3800 1392.0600 785.8600 ;
        RECT 1390.4600 790.8200 1392.0600 791.3000 ;
        RECT 1345.4600 796.2600 1347.0600 796.7400 ;
        RECT 1345.4600 801.7000 1347.0600 802.1800 ;
        RECT 1345.4600 779.9400 1347.0600 780.4200 ;
        RECT 1345.4600 785.3800 1347.0600 785.8600 ;
        RECT 1345.4600 790.8200 1347.0600 791.3000 ;
        RECT 1390.4600 769.0600 1392.0600 769.5400 ;
        RECT 1390.4600 774.5000 1392.0600 774.9800 ;
        RECT 1390.4600 752.7400 1392.0600 753.2200 ;
        RECT 1390.4600 758.1800 1392.0600 758.6600 ;
        RECT 1390.4600 763.6200 1392.0600 764.1000 ;
        RECT 1345.4600 769.0600 1347.0600 769.5400 ;
        RECT 1345.4600 774.5000 1347.0600 774.9800 ;
        RECT 1345.4600 752.7400 1347.0600 753.2200 ;
        RECT 1345.4600 758.1800 1347.0600 758.6600 ;
        RECT 1345.4600 763.6200 1347.0600 764.1000 ;
        RECT 1300.4600 796.2600 1302.0600 796.7400 ;
        RECT 1300.4600 801.7000 1302.0600 802.1800 ;
        RECT 1293.3000 796.2600 1294.9000 796.7400 ;
        RECT 1293.3000 801.7000 1294.9000 802.1800 ;
        RECT 1300.4600 779.9400 1302.0600 780.4200 ;
        RECT 1300.4600 785.3800 1302.0600 785.8600 ;
        RECT 1300.4600 790.8200 1302.0600 791.3000 ;
        RECT 1293.3000 779.9400 1294.9000 780.4200 ;
        RECT 1293.3000 785.3800 1294.9000 785.8600 ;
        RECT 1293.3000 790.8200 1294.9000 791.3000 ;
        RECT 1300.4600 769.0600 1302.0600 769.5400 ;
        RECT 1300.4600 774.5000 1302.0600 774.9800 ;
        RECT 1293.3000 769.0600 1294.9000 769.5400 ;
        RECT 1293.3000 774.5000 1294.9000 774.9800 ;
        RECT 1300.4600 752.7400 1302.0600 753.2200 ;
        RECT 1300.4600 758.1800 1302.0600 758.6600 ;
        RECT 1300.4600 763.6200 1302.0600 764.1000 ;
        RECT 1293.3000 752.7400 1294.9000 753.2200 ;
        RECT 1293.3000 758.1800 1294.9000 758.6600 ;
        RECT 1293.3000 763.6200 1294.9000 764.1000 ;
        RECT 1293.3000 807.1400 1294.9000 807.6200 ;
        RECT 1300.4600 807.1400 1302.0600 807.6200 ;
        RECT 1345.4600 807.1400 1347.0600 807.6200 ;
        RECT 1390.4600 807.1400 1392.0600 807.6200 ;
        RECT 1496.0000 741.8600 1497.6000 742.3400 ;
        RECT 1496.0000 747.3000 1497.6000 747.7800 ;
        RECT 1480.4600 741.8600 1482.0600 742.3400 ;
        RECT 1480.4600 747.3000 1482.0600 747.7800 ;
        RECT 1496.0000 725.5400 1497.6000 726.0200 ;
        RECT 1496.0000 730.9800 1497.6000 731.4600 ;
        RECT 1496.0000 736.4200 1497.6000 736.9000 ;
        RECT 1480.4600 725.5400 1482.0600 726.0200 ;
        RECT 1480.4600 730.9800 1482.0600 731.4600 ;
        RECT 1480.4600 736.4200 1482.0600 736.9000 ;
        RECT 1496.0000 714.6600 1497.6000 715.1400 ;
        RECT 1496.0000 720.1000 1497.6000 720.5800 ;
        RECT 1480.4600 714.6600 1482.0600 715.1400 ;
        RECT 1480.4600 720.1000 1482.0600 720.5800 ;
        RECT 1496.0000 698.3400 1497.6000 698.8200 ;
        RECT 1496.0000 703.7800 1497.6000 704.2600 ;
        RECT 1496.0000 709.2200 1497.6000 709.7000 ;
        RECT 1480.4600 698.3400 1482.0600 698.8200 ;
        RECT 1480.4600 703.7800 1482.0600 704.2600 ;
        RECT 1480.4600 709.2200 1482.0600 709.7000 ;
        RECT 1435.4600 741.8600 1437.0600 742.3400 ;
        RECT 1435.4600 747.3000 1437.0600 747.7800 ;
        RECT 1435.4600 725.5400 1437.0600 726.0200 ;
        RECT 1435.4600 730.9800 1437.0600 731.4600 ;
        RECT 1435.4600 736.4200 1437.0600 736.9000 ;
        RECT 1435.4600 714.6600 1437.0600 715.1400 ;
        RECT 1435.4600 720.1000 1437.0600 720.5800 ;
        RECT 1435.4600 698.3400 1437.0600 698.8200 ;
        RECT 1435.4600 703.7800 1437.0600 704.2600 ;
        RECT 1435.4600 709.2200 1437.0600 709.7000 ;
        RECT 1496.0000 687.4600 1497.6000 687.9400 ;
        RECT 1496.0000 692.9000 1497.6000 693.3800 ;
        RECT 1480.4600 687.4600 1482.0600 687.9400 ;
        RECT 1480.4600 692.9000 1482.0600 693.3800 ;
        RECT 1496.0000 671.1400 1497.6000 671.6200 ;
        RECT 1496.0000 676.5800 1497.6000 677.0600 ;
        RECT 1496.0000 682.0200 1497.6000 682.5000 ;
        RECT 1480.4600 671.1400 1482.0600 671.6200 ;
        RECT 1480.4600 676.5800 1482.0600 677.0600 ;
        RECT 1480.4600 682.0200 1482.0600 682.5000 ;
        RECT 1496.0000 660.2600 1497.6000 660.7400 ;
        RECT 1496.0000 665.7000 1497.6000 666.1800 ;
        RECT 1480.4600 660.2600 1482.0600 660.7400 ;
        RECT 1480.4600 665.7000 1482.0600 666.1800 ;
        RECT 1480.4600 654.8200 1482.0600 655.3000 ;
        RECT 1496.0000 654.8200 1497.6000 655.3000 ;
        RECT 1435.4600 687.4600 1437.0600 687.9400 ;
        RECT 1435.4600 692.9000 1437.0600 693.3800 ;
        RECT 1435.4600 671.1400 1437.0600 671.6200 ;
        RECT 1435.4600 676.5800 1437.0600 677.0600 ;
        RECT 1435.4600 682.0200 1437.0600 682.5000 ;
        RECT 1435.4600 660.2600 1437.0600 660.7400 ;
        RECT 1435.4600 665.7000 1437.0600 666.1800 ;
        RECT 1435.4600 654.8200 1437.0600 655.3000 ;
        RECT 1390.4600 741.8600 1392.0600 742.3400 ;
        RECT 1390.4600 747.3000 1392.0600 747.7800 ;
        RECT 1390.4600 725.5400 1392.0600 726.0200 ;
        RECT 1390.4600 730.9800 1392.0600 731.4600 ;
        RECT 1390.4600 736.4200 1392.0600 736.9000 ;
        RECT 1345.4600 741.8600 1347.0600 742.3400 ;
        RECT 1345.4600 747.3000 1347.0600 747.7800 ;
        RECT 1345.4600 725.5400 1347.0600 726.0200 ;
        RECT 1345.4600 730.9800 1347.0600 731.4600 ;
        RECT 1345.4600 736.4200 1347.0600 736.9000 ;
        RECT 1390.4600 714.6600 1392.0600 715.1400 ;
        RECT 1390.4600 720.1000 1392.0600 720.5800 ;
        RECT 1390.4600 698.3400 1392.0600 698.8200 ;
        RECT 1390.4600 703.7800 1392.0600 704.2600 ;
        RECT 1390.4600 709.2200 1392.0600 709.7000 ;
        RECT 1345.4600 714.6600 1347.0600 715.1400 ;
        RECT 1345.4600 720.1000 1347.0600 720.5800 ;
        RECT 1345.4600 698.3400 1347.0600 698.8200 ;
        RECT 1345.4600 703.7800 1347.0600 704.2600 ;
        RECT 1345.4600 709.2200 1347.0600 709.7000 ;
        RECT 1300.4600 741.8600 1302.0600 742.3400 ;
        RECT 1300.4600 747.3000 1302.0600 747.7800 ;
        RECT 1293.3000 741.8600 1294.9000 742.3400 ;
        RECT 1293.3000 747.3000 1294.9000 747.7800 ;
        RECT 1300.4600 725.5400 1302.0600 726.0200 ;
        RECT 1300.4600 730.9800 1302.0600 731.4600 ;
        RECT 1300.4600 736.4200 1302.0600 736.9000 ;
        RECT 1293.3000 725.5400 1294.9000 726.0200 ;
        RECT 1293.3000 730.9800 1294.9000 731.4600 ;
        RECT 1293.3000 736.4200 1294.9000 736.9000 ;
        RECT 1300.4600 714.6600 1302.0600 715.1400 ;
        RECT 1300.4600 720.1000 1302.0600 720.5800 ;
        RECT 1293.3000 714.6600 1294.9000 715.1400 ;
        RECT 1293.3000 720.1000 1294.9000 720.5800 ;
        RECT 1300.4600 698.3400 1302.0600 698.8200 ;
        RECT 1300.4600 703.7800 1302.0600 704.2600 ;
        RECT 1300.4600 709.2200 1302.0600 709.7000 ;
        RECT 1293.3000 698.3400 1294.9000 698.8200 ;
        RECT 1293.3000 703.7800 1294.9000 704.2600 ;
        RECT 1293.3000 709.2200 1294.9000 709.7000 ;
        RECT 1390.4600 687.4600 1392.0600 687.9400 ;
        RECT 1390.4600 692.9000 1392.0600 693.3800 ;
        RECT 1390.4600 671.1400 1392.0600 671.6200 ;
        RECT 1390.4600 676.5800 1392.0600 677.0600 ;
        RECT 1390.4600 682.0200 1392.0600 682.5000 ;
        RECT 1345.4600 687.4600 1347.0600 687.9400 ;
        RECT 1345.4600 692.9000 1347.0600 693.3800 ;
        RECT 1345.4600 671.1400 1347.0600 671.6200 ;
        RECT 1345.4600 676.5800 1347.0600 677.0600 ;
        RECT 1345.4600 682.0200 1347.0600 682.5000 ;
        RECT 1390.4600 665.7000 1392.0600 666.1800 ;
        RECT 1390.4600 660.2600 1392.0600 660.7400 ;
        RECT 1390.4600 654.8200 1392.0600 655.3000 ;
        RECT 1345.4600 665.7000 1347.0600 666.1800 ;
        RECT 1345.4600 660.2600 1347.0600 660.7400 ;
        RECT 1345.4600 654.8200 1347.0600 655.3000 ;
        RECT 1300.4600 687.4600 1302.0600 687.9400 ;
        RECT 1300.4600 692.9000 1302.0600 693.3800 ;
        RECT 1293.3000 687.4600 1294.9000 687.9400 ;
        RECT 1293.3000 692.9000 1294.9000 693.3800 ;
        RECT 1300.4600 671.1400 1302.0600 671.6200 ;
        RECT 1300.4600 676.5800 1302.0600 677.0600 ;
        RECT 1300.4600 682.0200 1302.0600 682.5000 ;
        RECT 1293.3000 671.1400 1294.9000 671.6200 ;
        RECT 1293.3000 676.5800 1294.9000 677.0600 ;
        RECT 1293.3000 682.0200 1294.9000 682.5000 ;
        RECT 1300.4600 660.2600 1302.0600 660.7400 ;
        RECT 1300.4600 665.7000 1302.0600 666.1800 ;
        RECT 1293.3000 660.2600 1294.9000 660.7400 ;
        RECT 1293.3000 665.7000 1294.9000 666.1800 ;
        RECT 1293.3000 654.8200 1294.9000 655.3000 ;
        RECT 1300.4600 654.8200 1302.0600 655.3000 ;
        RECT 1290.3400 857.0100 1500.5600 858.6100 ;
        RECT 1290.3400 645.3100 1500.5600 646.9100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 642.4800 1294.9000 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 860.5200 1294.9000 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 642.4800 1497.6000 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 860.5200 1497.6000 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 645.3100 1291.9400 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 645.3100 1500.5600 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 857.0100 1291.9400 858.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 857.0100 1500.5600 858.6100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1480.4600 415.6700 1482.0600 628.9700 ;
        RECT 1435.4600 415.6700 1437.0600 628.9700 ;
        RECT 1390.4600 415.6700 1392.0600 628.9700 ;
        RECT 1345.4600 415.6700 1347.0600 628.9700 ;
        RECT 1300.4600 415.6700 1302.0600 628.9700 ;
        RECT 1496.0000 412.8400 1497.6000 632.4800 ;
        RECT 1293.3000 412.8400 1294.9000 632.4800 ;
      LAYER met3 ;
        RECT 1480.4600 621.0200 1482.0600 621.5000 ;
        RECT 1496.0000 621.0200 1497.6000 621.5000 ;
        RECT 1496.0000 610.1400 1497.6000 610.6200 ;
        RECT 1496.0000 615.5800 1497.6000 616.0600 ;
        RECT 1480.4600 610.1400 1482.0600 610.6200 ;
        RECT 1480.4600 615.5800 1482.0600 616.0600 ;
        RECT 1496.0000 593.8200 1497.6000 594.3000 ;
        RECT 1496.0000 599.2600 1497.6000 599.7400 ;
        RECT 1480.4600 593.8200 1482.0600 594.3000 ;
        RECT 1480.4600 599.2600 1482.0600 599.7400 ;
        RECT 1496.0000 582.9400 1497.6000 583.4200 ;
        RECT 1496.0000 588.3800 1497.6000 588.8600 ;
        RECT 1480.4600 582.9400 1482.0600 583.4200 ;
        RECT 1480.4600 588.3800 1482.0600 588.8600 ;
        RECT 1480.4600 604.7000 1482.0600 605.1800 ;
        RECT 1496.0000 604.7000 1497.6000 605.1800 ;
        RECT 1435.4600 610.1400 1437.0600 610.6200 ;
        RECT 1435.4600 615.5800 1437.0600 616.0600 ;
        RECT 1435.4600 621.0200 1437.0600 621.5000 ;
        RECT 1435.4600 593.8200 1437.0600 594.3000 ;
        RECT 1435.4600 599.2600 1437.0600 599.7400 ;
        RECT 1435.4600 588.3800 1437.0600 588.8600 ;
        RECT 1435.4600 582.9400 1437.0600 583.4200 ;
        RECT 1435.4600 604.7000 1437.0600 605.1800 ;
        RECT 1496.0000 566.6200 1497.6000 567.1000 ;
        RECT 1496.0000 572.0600 1497.6000 572.5400 ;
        RECT 1480.4600 566.6200 1482.0600 567.1000 ;
        RECT 1480.4600 572.0600 1482.0600 572.5400 ;
        RECT 1496.0000 550.3000 1497.6000 550.7800 ;
        RECT 1496.0000 555.7400 1497.6000 556.2200 ;
        RECT 1496.0000 561.1800 1497.6000 561.6600 ;
        RECT 1480.4600 550.3000 1482.0600 550.7800 ;
        RECT 1480.4600 555.7400 1482.0600 556.2200 ;
        RECT 1480.4600 561.1800 1482.0600 561.6600 ;
        RECT 1496.0000 539.4200 1497.6000 539.9000 ;
        RECT 1496.0000 544.8600 1497.6000 545.3400 ;
        RECT 1480.4600 539.4200 1482.0600 539.9000 ;
        RECT 1480.4600 544.8600 1482.0600 545.3400 ;
        RECT 1496.0000 523.1000 1497.6000 523.5800 ;
        RECT 1496.0000 528.5400 1497.6000 529.0200 ;
        RECT 1496.0000 533.9800 1497.6000 534.4600 ;
        RECT 1480.4600 523.1000 1482.0600 523.5800 ;
        RECT 1480.4600 528.5400 1482.0600 529.0200 ;
        RECT 1480.4600 533.9800 1482.0600 534.4600 ;
        RECT 1435.4600 566.6200 1437.0600 567.1000 ;
        RECT 1435.4600 572.0600 1437.0600 572.5400 ;
        RECT 1435.4600 550.3000 1437.0600 550.7800 ;
        RECT 1435.4600 555.7400 1437.0600 556.2200 ;
        RECT 1435.4600 561.1800 1437.0600 561.6600 ;
        RECT 1435.4600 539.4200 1437.0600 539.9000 ;
        RECT 1435.4600 544.8600 1437.0600 545.3400 ;
        RECT 1435.4600 523.1000 1437.0600 523.5800 ;
        RECT 1435.4600 528.5400 1437.0600 529.0200 ;
        RECT 1435.4600 533.9800 1437.0600 534.4600 ;
        RECT 1435.4600 577.5000 1437.0600 577.9800 ;
        RECT 1480.4600 577.5000 1482.0600 577.9800 ;
        RECT 1496.0000 577.5000 1497.6000 577.9800 ;
        RECT 1390.4600 610.1400 1392.0600 610.6200 ;
        RECT 1390.4600 615.5800 1392.0600 616.0600 ;
        RECT 1390.4600 621.0200 1392.0600 621.5000 ;
        RECT 1345.4600 610.1400 1347.0600 610.6200 ;
        RECT 1345.4600 615.5800 1347.0600 616.0600 ;
        RECT 1345.4600 621.0200 1347.0600 621.5000 ;
        RECT 1390.4600 593.8200 1392.0600 594.3000 ;
        RECT 1390.4600 599.2600 1392.0600 599.7400 ;
        RECT 1390.4600 582.9400 1392.0600 583.4200 ;
        RECT 1390.4600 588.3800 1392.0600 588.8600 ;
        RECT 1345.4600 593.8200 1347.0600 594.3000 ;
        RECT 1345.4600 599.2600 1347.0600 599.7400 ;
        RECT 1345.4600 582.9400 1347.0600 583.4200 ;
        RECT 1345.4600 588.3800 1347.0600 588.8600 ;
        RECT 1345.4600 604.7000 1347.0600 605.1800 ;
        RECT 1390.4600 604.7000 1392.0600 605.1800 ;
        RECT 1293.3000 621.0200 1294.9000 621.5000 ;
        RECT 1300.4600 621.0200 1302.0600 621.5000 ;
        RECT 1300.4600 610.1400 1302.0600 610.6200 ;
        RECT 1300.4600 615.5800 1302.0600 616.0600 ;
        RECT 1293.3000 610.1400 1294.9000 610.6200 ;
        RECT 1293.3000 615.5800 1294.9000 616.0600 ;
        RECT 1300.4600 593.8200 1302.0600 594.3000 ;
        RECT 1300.4600 599.2600 1302.0600 599.7400 ;
        RECT 1293.3000 593.8200 1294.9000 594.3000 ;
        RECT 1293.3000 599.2600 1294.9000 599.7400 ;
        RECT 1300.4600 582.9400 1302.0600 583.4200 ;
        RECT 1300.4600 588.3800 1302.0600 588.8600 ;
        RECT 1293.3000 582.9400 1294.9000 583.4200 ;
        RECT 1293.3000 588.3800 1294.9000 588.8600 ;
        RECT 1293.3000 604.7000 1294.9000 605.1800 ;
        RECT 1300.4600 604.7000 1302.0600 605.1800 ;
        RECT 1390.4600 566.6200 1392.0600 567.1000 ;
        RECT 1390.4600 572.0600 1392.0600 572.5400 ;
        RECT 1390.4600 550.3000 1392.0600 550.7800 ;
        RECT 1390.4600 555.7400 1392.0600 556.2200 ;
        RECT 1390.4600 561.1800 1392.0600 561.6600 ;
        RECT 1345.4600 566.6200 1347.0600 567.1000 ;
        RECT 1345.4600 572.0600 1347.0600 572.5400 ;
        RECT 1345.4600 550.3000 1347.0600 550.7800 ;
        RECT 1345.4600 555.7400 1347.0600 556.2200 ;
        RECT 1345.4600 561.1800 1347.0600 561.6600 ;
        RECT 1390.4600 539.4200 1392.0600 539.9000 ;
        RECT 1390.4600 544.8600 1392.0600 545.3400 ;
        RECT 1390.4600 523.1000 1392.0600 523.5800 ;
        RECT 1390.4600 528.5400 1392.0600 529.0200 ;
        RECT 1390.4600 533.9800 1392.0600 534.4600 ;
        RECT 1345.4600 539.4200 1347.0600 539.9000 ;
        RECT 1345.4600 544.8600 1347.0600 545.3400 ;
        RECT 1345.4600 523.1000 1347.0600 523.5800 ;
        RECT 1345.4600 528.5400 1347.0600 529.0200 ;
        RECT 1345.4600 533.9800 1347.0600 534.4600 ;
        RECT 1300.4600 566.6200 1302.0600 567.1000 ;
        RECT 1300.4600 572.0600 1302.0600 572.5400 ;
        RECT 1293.3000 566.6200 1294.9000 567.1000 ;
        RECT 1293.3000 572.0600 1294.9000 572.5400 ;
        RECT 1300.4600 550.3000 1302.0600 550.7800 ;
        RECT 1300.4600 555.7400 1302.0600 556.2200 ;
        RECT 1300.4600 561.1800 1302.0600 561.6600 ;
        RECT 1293.3000 550.3000 1294.9000 550.7800 ;
        RECT 1293.3000 555.7400 1294.9000 556.2200 ;
        RECT 1293.3000 561.1800 1294.9000 561.6600 ;
        RECT 1300.4600 539.4200 1302.0600 539.9000 ;
        RECT 1300.4600 544.8600 1302.0600 545.3400 ;
        RECT 1293.3000 539.4200 1294.9000 539.9000 ;
        RECT 1293.3000 544.8600 1294.9000 545.3400 ;
        RECT 1300.4600 523.1000 1302.0600 523.5800 ;
        RECT 1300.4600 528.5400 1302.0600 529.0200 ;
        RECT 1300.4600 533.9800 1302.0600 534.4600 ;
        RECT 1293.3000 523.1000 1294.9000 523.5800 ;
        RECT 1293.3000 528.5400 1294.9000 529.0200 ;
        RECT 1293.3000 533.9800 1294.9000 534.4600 ;
        RECT 1293.3000 577.5000 1294.9000 577.9800 ;
        RECT 1300.4600 577.5000 1302.0600 577.9800 ;
        RECT 1345.4600 577.5000 1347.0600 577.9800 ;
        RECT 1390.4600 577.5000 1392.0600 577.9800 ;
        RECT 1496.0000 512.2200 1497.6000 512.7000 ;
        RECT 1496.0000 517.6600 1497.6000 518.1400 ;
        RECT 1480.4600 512.2200 1482.0600 512.7000 ;
        RECT 1480.4600 517.6600 1482.0600 518.1400 ;
        RECT 1496.0000 495.9000 1497.6000 496.3800 ;
        RECT 1496.0000 501.3400 1497.6000 501.8200 ;
        RECT 1496.0000 506.7800 1497.6000 507.2600 ;
        RECT 1480.4600 495.9000 1482.0600 496.3800 ;
        RECT 1480.4600 501.3400 1482.0600 501.8200 ;
        RECT 1480.4600 506.7800 1482.0600 507.2600 ;
        RECT 1496.0000 485.0200 1497.6000 485.5000 ;
        RECT 1496.0000 490.4600 1497.6000 490.9400 ;
        RECT 1480.4600 485.0200 1482.0600 485.5000 ;
        RECT 1480.4600 490.4600 1482.0600 490.9400 ;
        RECT 1496.0000 468.7000 1497.6000 469.1800 ;
        RECT 1496.0000 474.1400 1497.6000 474.6200 ;
        RECT 1496.0000 479.5800 1497.6000 480.0600 ;
        RECT 1480.4600 468.7000 1482.0600 469.1800 ;
        RECT 1480.4600 474.1400 1482.0600 474.6200 ;
        RECT 1480.4600 479.5800 1482.0600 480.0600 ;
        RECT 1435.4600 512.2200 1437.0600 512.7000 ;
        RECT 1435.4600 517.6600 1437.0600 518.1400 ;
        RECT 1435.4600 495.9000 1437.0600 496.3800 ;
        RECT 1435.4600 501.3400 1437.0600 501.8200 ;
        RECT 1435.4600 506.7800 1437.0600 507.2600 ;
        RECT 1435.4600 485.0200 1437.0600 485.5000 ;
        RECT 1435.4600 490.4600 1437.0600 490.9400 ;
        RECT 1435.4600 468.7000 1437.0600 469.1800 ;
        RECT 1435.4600 474.1400 1437.0600 474.6200 ;
        RECT 1435.4600 479.5800 1437.0600 480.0600 ;
        RECT 1496.0000 457.8200 1497.6000 458.3000 ;
        RECT 1496.0000 463.2600 1497.6000 463.7400 ;
        RECT 1480.4600 457.8200 1482.0600 458.3000 ;
        RECT 1480.4600 463.2600 1482.0600 463.7400 ;
        RECT 1496.0000 441.5000 1497.6000 441.9800 ;
        RECT 1496.0000 446.9400 1497.6000 447.4200 ;
        RECT 1496.0000 452.3800 1497.6000 452.8600 ;
        RECT 1480.4600 441.5000 1482.0600 441.9800 ;
        RECT 1480.4600 446.9400 1482.0600 447.4200 ;
        RECT 1480.4600 452.3800 1482.0600 452.8600 ;
        RECT 1496.0000 430.6200 1497.6000 431.1000 ;
        RECT 1496.0000 436.0600 1497.6000 436.5400 ;
        RECT 1480.4600 430.6200 1482.0600 431.1000 ;
        RECT 1480.4600 436.0600 1482.0600 436.5400 ;
        RECT 1480.4600 425.1800 1482.0600 425.6600 ;
        RECT 1496.0000 425.1800 1497.6000 425.6600 ;
        RECT 1435.4600 457.8200 1437.0600 458.3000 ;
        RECT 1435.4600 463.2600 1437.0600 463.7400 ;
        RECT 1435.4600 441.5000 1437.0600 441.9800 ;
        RECT 1435.4600 446.9400 1437.0600 447.4200 ;
        RECT 1435.4600 452.3800 1437.0600 452.8600 ;
        RECT 1435.4600 430.6200 1437.0600 431.1000 ;
        RECT 1435.4600 436.0600 1437.0600 436.5400 ;
        RECT 1435.4600 425.1800 1437.0600 425.6600 ;
        RECT 1390.4600 512.2200 1392.0600 512.7000 ;
        RECT 1390.4600 517.6600 1392.0600 518.1400 ;
        RECT 1390.4600 495.9000 1392.0600 496.3800 ;
        RECT 1390.4600 501.3400 1392.0600 501.8200 ;
        RECT 1390.4600 506.7800 1392.0600 507.2600 ;
        RECT 1345.4600 512.2200 1347.0600 512.7000 ;
        RECT 1345.4600 517.6600 1347.0600 518.1400 ;
        RECT 1345.4600 495.9000 1347.0600 496.3800 ;
        RECT 1345.4600 501.3400 1347.0600 501.8200 ;
        RECT 1345.4600 506.7800 1347.0600 507.2600 ;
        RECT 1390.4600 485.0200 1392.0600 485.5000 ;
        RECT 1390.4600 490.4600 1392.0600 490.9400 ;
        RECT 1390.4600 468.7000 1392.0600 469.1800 ;
        RECT 1390.4600 474.1400 1392.0600 474.6200 ;
        RECT 1390.4600 479.5800 1392.0600 480.0600 ;
        RECT 1345.4600 485.0200 1347.0600 485.5000 ;
        RECT 1345.4600 490.4600 1347.0600 490.9400 ;
        RECT 1345.4600 468.7000 1347.0600 469.1800 ;
        RECT 1345.4600 474.1400 1347.0600 474.6200 ;
        RECT 1345.4600 479.5800 1347.0600 480.0600 ;
        RECT 1300.4600 512.2200 1302.0600 512.7000 ;
        RECT 1300.4600 517.6600 1302.0600 518.1400 ;
        RECT 1293.3000 512.2200 1294.9000 512.7000 ;
        RECT 1293.3000 517.6600 1294.9000 518.1400 ;
        RECT 1300.4600 495.9000 1302.0600 496.3800 ;
        RECT 1300.4600 501.3400 1302.0600 501.8200 ;
        RECT 1300.4600 506.7800 1302.0600 507.2600 ;
        RECT 1293.3000 495.9000 1294.9000 496.3800 ;
        RECT 1293.3000 501.3400 1294.9000 501.8200 ;
        RECT 1293.3000 506.7800 1294.9000 507.2600 ;
        RECT 1300.4600 485.0200 1302.0600 485.5000 ;
        RECT 1300.4600 490.4600 1302.0600 490.9400 ;
        RECT 1293.3000 485.0200 1294.9000 485.5000 ;
        RECT 1293.3000 490.4600 1294.9000 490.9400 ;
        RECT 1300.4600 468.7000 1302.0600 469.1800 ;
        RECT 1300.4600 474.1400 1302.0600 474.6200 ;
        RECT 1300.4600 479.5800 1302.0600 480.0600 ;
        RECT 1293.3000 468.7000 1294.9000 469.1800 ;
        RECT 1293.3000 474.1400 1294.9000 474.6200 ;
        RECT 1293.3000 479.5800 1294.9000 480.0600 ;
        RECT 1390.4600 457.8200 1392.0600 458.3000 ;
        RECT 1390.4600 463.2600 1392.0600 463.7400 ;
        RECT 1390.4600 441.5000 1392.0600 441.9800 ;
        RECT 1390.4600 446.9400 1392.0600 447.4200 ;
        RECT 1390.4600 452.3800 1392.0600 452.8600 ;
        RECT 1345.4600 457.8200 1347.0600 458.3000 ;
        RECT 1345.4600 463.2600 1347.0600 463.7400 ;
        RECT 1345.4600 441.5000 1347.0600 441.9800 ;
        RECT 1345.4600 446.9400 1347.0600 447.4200 ;
        RECT 1345.4600 452.3800 1347.0600 452.8600 ;
        RECT 1390.4600 436.0600 1392.0600 436.5400 ;
        RECT 1390.4600 430.6200 1392.0600 431.1000 ;
        RECT 1390.4600 425.1800 1392.0600 425.6600 ;
        RECT 1345.4600 436.0600 1347.0600 436.5400 ;
        RECT 1345.4600 430.6200 1347.0600 431.1000 ;
        RECT 1345.4600 425.1800 1347.0600 425.6600 ;
        RECT 1300.4600 457.8200 1302.0600 458.3000 ;
        RECT 1300.4600 463.2600 1302.0600 463.7400 ;
        RECT 1293.3000 457.8200 1294.9000 458.3000 ;
        RECT 1293.3000 463.2600 1294.9000 463.7400 ;
        RECT 1300.4600 441.5000 1302.0600 441.9800 ;
        RECT 1300.4600 446.9400 1302.0600 447.4200 ;
        RECT 1300.4600 452.3800 1302.0600 452.8600 ;
        RECT 1293.3000 441.5000 1294.9000 441.9800 ;
        RECT 1293.3000 446.9400 1294.9000 447.4200 ;
        RECT 1293.3000 452.3800 1294.9000 452.8600 ;
        RECT 1300.4600 430.6200 1302.0600 431.1000 ;
        RECT 1300.4600 436.0600 1302.0600 436.5400 ;
        RECT 1293.3000 430.6200 1294.9000 431.1000 ;
        RECT 1293.3000 436.0600 1294.9000 436.5400 ;
        RECT 1293.3000 425.1800 1294.9000 425.6600 ;
        RECT 1300.4600 425.1800 1302.0600 425.6600 ;
        RECT 1290.3400 627.3700 1500.5600 628.9700 ;
        RECT 1290.3400 415.6700 1500.5600 417.2700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 412.8400 1294.9000 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1293.3000 630.8800 1294.9000 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 412.8400 1497.6000 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1496.0000 630.8800 1497.6000 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 415.6700 1291.9400 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 415.6700 1500.5600 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 627.3700 1291.9400 628.9700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 627.3700 1500.5600 628.9700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1513.6200 2479.6000 1515.2200 2509.8600 ;
        RECT 1716.1200 2479.6000 1717.7200 2509.8600 ;
      LAYER met3 ;
        RECT 1716.1200 2500.1000 1717.7200 2500.5800 ;
        RECT 1513.6200 2500.1000 1515.2200 2500.5800 ;
        RECT 1716.1200 2489.2200 1717.7200 2489.7000 ;
        RECT 1513.6200 2489.2200 1515.2200 2489.7000 ;
        RECT 1716.1200 2494.6600 1717.7200 2495.1400 ;
        RECT 1513.6200 2494.6600 1515.2200 2495.1400 ;
        RECT 1510.5600 2505.5000 1720.7800 2507.1000 ;
        RECT 1510.5600 2481.1700 1720.7800 2482.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.6200 2479.6000 1515.2200 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.6200 2508.2600 1515.2200 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.1200 2479.6000 1717.7200 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.1200 2508.2600 1717.7200 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2481.1700 1512.1600 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2481.1700 1720.7800 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2505.5000 1512.1600 2507.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2505.5000 1720.7800 2507.1000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 186.0300 1702.2800 399.3300 ;
        RECT 1655.6800 186.0300 1657.2800 399.3300 ;
        RECT 1610.6800 186.0300 1612.2800 399.3300 ;
        RECT 1565.6800 186.0300 1567.2800 399.3300 ;
        RECT 1520.6800 186.0300 1522.2800 399.3300 ;
        RECT 1716.2200 183.2000 1717.8200 402.8400 ;
        RECT 1513.5200 183.2000 1515.1200 402.8400 ;
      LAYER met3 ;
        RECT 1700.6800 391.3800 1702.2800 391.8600 ;
        RECT 1716.2200 391.3800 1717.8200 391.8600 ;
        RECT 1716.2200 380.5000 1717.8200 380.9800 ;
        RECT 1716.2200 385.9400 1717.8200 386.4200 ;
        RECT 1700.6800 380.5000 1702.2800 380.9800 ;
        RECT 1700.6800 385.9400 1702.2800 386.4200 ;
        RECT 1716.2200 364.1800 1717.8200 364.6600 ;
        RECT 1716.2200 369.6200 1717.8200 370.1000 ;
        RECT 1700.6800 364.1800 1702.2800 364.6600 ;
        RECT 1700.6800 369.6200 1702.2800 370.1000 ;
        RECT 1716.2200 353.3000 1717.8200 353.7800 ;
        RECT 1716.2200 358.7400 1717.8200 359.2200 ;
        RECT 1700.6800 353.3000 1702.2800 353.7800 ;
        RECT 1700.6800 358.7400 1702.2800 359.2200 ;
        RECT 1700.6800 375.0600 1702.2800 375.5400 ;
        RECT 1716.2200 375.0600 1717.8200 375.5400 ;
        RECT 1655.6800 380.5000 1657.2800 380.9800 ;
        RECT 1655.6800 385.9400 1657.2800 386.4200 ;
        RECT 1655.6800 391.3800 1657.2800 391.8600 ;
        RECT 1655.6800 364.1800 1657.2800 364.6600 ;
        RECT 1655.6800 369.6200 1657.2800 370.1000 ;
        RECT 1655.6800 358.7400 1657.2800 359.2200 ;
        RECT 1655.6800 353.3000 1657.2800 353.7800 ;
        RECT 1655.6800 375.0600 1657.2800 375.5400 ;
        RECT 1716.2200 336.9800 1717.8200 337.4600 ;
        RECT 1716.2200 342.4200 1717.8200 342.9000 ;
        RECT 1700.6800 336.9800 1702.2800 337.4600 ;
        RECT 1700.6800 342.4200 1702.2800 342.9000 ;
        RECT 1716.2200 320.6600 1717.8200 321.1400 ;
        RECT 1716.2200 326.1000 1717.8200 326.5800 ;
        RECT 1716.2200 331.5400 1717.8200 332.0200 ;
        RECT 1700.6800 320.6600 1702.2800 321.1400 ;
        RECT 1700.6800 326.1000 1702.2800 326.5800 ;
        RECT 1700.6800 331.5400 1702.2800 332.0200 ;
        RECT 1716.2200 309.7800 1717.8200 310.2600 ;
        RECT 1716.2200 315.2200 1717.8200 315.7000 ;
        RECT 1700.6800 309.7800 1702.2800 310.2600 ;
        RECT 1700.6800 315.2200 1702.2800 315.7000 ;
        RECT 1716.2200 293.4600 1717.8200 293.9400 ;
        RECT 1716.2200 298.9000 1717.8200 299.3800 ;
        RECT 1716.2200 304.3400 1717.8200 304.8200 ;
        RECT 1700.6800 293.4600 1702.2800 293.9400 ;
        RECT 1700.6800 298.9000 1702.2800 299.3800 ;
        RECT 1700.6800 304.3400 1702.2800 304.8200 ;
        RECT 1655.6800 336.9800 1657.2800 337.4600 ;
        RECT 1655.6800 342.4200 1657.2800 342.9000 ;
        RECT 1655.6800 320.6600 1657.2800 321.1400 ;
        RECT 1655.6800 326.1000 1657.2800 326.5800 ;
        RECT 1655.6800 331.5400 1657.2800 332.0200 ;
        RECT 1655.6800 309.7800 1657.2800 310.2600 ;
        RECT 1655.6800 315.2200 1657.2800 315.7000 ;
        RECT 1655.6800 293.4600 1657.2800 293.9400 ;
        RECT 1655.6800 298.9000 1657.2800 299.3800 ;
        RECT 1655.6800 304.3400 1657.2800 304.8200 ;
        RECT 1655.6800 347.8600 1657.2800 348.3400 ;
        RECT 1700.6800 347.8600 1702.2800 348.3400 ;
        RECT 1716.2200 347.8600 1717.8200 348.3400 ;
        RECT 1610.6800 380.5000 1612.2800 380.9800 ;
        RECT 1610.6800 385.9400 1612.2800 386.4200 ;
        RECT 1610.6800 391.3800 1612.2800 391.8600 ;
        RECT 1565.6800 380.5000 1567.2800 380.9800 ;
        RECT 1565.6800 385.9400 1567.2800 386.4200 ;
        RECT 1565.6800 391.3800 1567.2800 391.8600 ;
        RECT 1610.6800 364.1800 1612.2800 364.6600 ;
        RECT 1610.6800 369.6200 1612.2800 370.1000 ;
        RECT 1610.6800 353.3000 1612.2800 353.7800 ;
        RECT 1610.6800 358.7400 1612.2800 359.2200 ;
        RECT 1565.6800 364.1800 1567.2800 364.6600 ;
        RECT 1565.6800 369.6200 1567.2800 370.1000 ;
        RECT 1565.6800 353.3000 1567.2800 353.7800 ;
        RECT 1565.6800 358.7400 1567.2800 359.2200 ;
        RECT 1565.6800 375.0600 1567.2800 375.5400 ;
        RECT 1610.6800 375.0600 1612.2800 375.5400 ;
        RECT 1513.5200 391.3800 1515.1200 391.8600 ;
        RECT 1520.6800 391.3800 1522.2800 391.8600 ;
        RECT 1520.6800 380.5000 1522.2800 380.9800 ;
        RECT 1520.6800 385.9400 1522.2800 386.4200 ;
        RECT 1513.5200 380.5000 1515.1200 380.9800 ;
        RECT 1513.5200 385.9400 1515.1200 386.4200 ;
        RECT 1520.6800 364.1800 1522.2800 364.6600 ;
        RECT 1520.6800 369.6200 1522.2800 370.1000 ;
        RECT 1513.5200 364.1800 1515.1200 364.6600 ;
        RECT 1513.5200 369.6200 1515.1200 370.1000 ;
        RECT 1520.6800 353.3000 1522.2800 353.7800 ;
        RECT 1520.6800 358.7400 1522.2800 359.2200 ;
        RECT 1513.5200 353.3000 1515.1200 353.7800 ;
        RECT 1513.5200 358.7400 1515.1200 359.2200 ;
        RECT 1513.5200 375.0600 1515.1200 375.5400 ;
        RECT 1520.6800 375.0600 1522.2800 375.5400 ;
        RECT 1610.6800 336.9800 1612.2800 337.4600 ;
        RECT 1610.6800 342.4200 1612.2800 342.9000 ;
        RECT 1610.6800 320.6600 1612.2800 321.1400 ;
        RECT 1610.6800 326.1000 1612.2800 326.5800 ;
        RECT 1610.6800 331.5400 1612.2800 332.0200 ;
        RECT 1565.6800 336.9800 1567.2800 337.4600 ;
        RECT 1565.6800 342.4200 1567.2800 342.9000 ;
        RECT 1565.6800 320.6600 1567.2800 321.1400 ;
        RECT 1565.6800 326.1000 1567.2800 326.5800 ;
        RECT 1565.6800 331.5400 1567.2800 332.0200 ;
        RECT 1610.6800 309.7800 1612.2800 310.2600 ;
        RECT 1610.6800 315.2200 1612.2800 315.7000 ;
        RECT 1610.6800 293.4600 1612.2800 293.9400 ;
        RECT 1610.6800 298.9000 1612.2800 299.3800 ;
        RECT 1610.6800 304.3400 1612.2800 304.8200 ;
        RECT 1565.6800 309.7800 1567.2800 310.2600 ;
        RECT 1565.6800 315.2200 1567.2800 315.7000 ;
        RECT 1565.6800 293.4600 1567.2800 293.9400 ;
        RECT 1565.6800 298.9000 1567.2800 299.3800 ;
        RECT 1565.6800 304.3400 1567.2800 304.8200 ;
        RECT 1520.6800 336.9800 1522.2800 337.4600 ;
        RECT 1520.6800 342.4200 1522.2800 342.9000 ;
        RECT 1513.5200 336.9800 1515.1200 337.4600 ;
        RECT 1513.5200 342.4200 1515.1200 342.9000 ;
        RECT 1520.6800 320.6600 1522.2800 321.1400 ;
        RECT 1520.6800 326.1000 1522.2800 326.5800 ;
        RECT 1520.6800 331.5400 1522.2800 332.0200 ;
        RECT 1513.5200 320.6600 1515.1200 321.1400 ;
        RECT 1513.5200 326.1000 1515.1200 326.5800 ;
        RECT 1513.5200 331.5400 1515.1200 332.0200 ;
        RECT 1520.6800 309.7800 1522.2800 310.2600 ;
        RECT 1520.6800 315.2200 1522.2800 315.7000 ;
        RECT 1513.5200 309.7800 1515.1200 310.2600 ;
        RECT 1513.5200 315.2200 1515.1200 315.7000 ;
        RECT 1520.6800 293.4600 1522.2800 293.9400 ;
        RECT 1520.6800 298.9000 1522.2800 299.3800 ;
        RECT 1520.6800 304.3400 1522.2800 304.8200 ;
        RECT 1513.5200 293.4600 1515.1200 293.9400 ;
        RECT 1513.5200 298.9000 1515.1200 299.3800 ;
        RECT 1513.5200 304.3400 1515.1200 304.8200 ;
        RECT 1513.5200 347.8600 1515.1200 348.3400 ;
        RECT 1520.6800 347.8600 1522.2800 348.3400 ;
        RECT 1565.6800 347.8600 1567.2800 348.3400 ;
        RECT 1610.6800 347.8600 1612.2800 348.3400 ;
        RECT 1716.2200 282.5800 1717.8200 283.0600 ;
        RECT 1716.2200 288.0200 1717.8200 288.5000 ;
        RECT 1700.6800 282.5800 1702.2800 283.0600 ;
        RECT 1700.6800 288.0200 1702.2800 288.5000 ;
        RECT 1716.2200 266.2600 1717.8200 266.7400 ;
        RECT 1716.2200 271.7000 1717.8200 272.1800 ;
        RECT 1716.2200 277.1400 1717.8200 277.6200 ;
        RECT 1700.6800 266.2600 1702.2800 266.7400 ;
        RECT 1700.6800 271.7000 1702.2800 272.1800 ;
        RECT 1700.6800 277.1400 1702.2800 277.6200 ;
        RECT 1716.2200 255.3800 1717.8200 255.8600 ;
        RECT 1716.2200 260.8200 1717.8200 261.3000 ;
        RECT 1700.6800 255.3800 1702.2800 255.8600 ;
        RECT 1700.6800 260.8200 1702.2800 261.3000 ;
        RECT 1716.2200 239.0600 1717.8200 239.5400 ;
        RECT 1716.2200 244.5000 1717.8200 244.9800 ;
        RECT 1716.2200 249.9400 1717.8200 250.4200 ;
        RECT 1700.6800 239.0600 1702.2800 239.5400 ;
        RECT 1700.6800 244.5000 1702.2800 244.9800 ;
        RECT 1700.6800 249.9400 1702.2800 250.4200 ;
        RECT 1655.6800 282.5800 1657.2800 283.0600 ;
        RECT 1655.6800 288.0200 1657.2800 288.5000 ;
        RECT 1655.6800 266.2600 1657.2800 266.7400 ;
        RECT 1655.6800 271.7000 1657.2800 272.1800 ;
        RECT 1655.6800 277.1400 1657.2800 277.6200 ;
        RECT 1655.6800 255.3800 1657.2800 255.8600 ;
        RECT 1655.6800 260.8200 1657.2800 261.3000 ;
        RECT 1655.6800 239.0600 1657.2800 239.5400 ;
        RECT 1655.6800 244.5000 1657.2800 244.9800 ;
        RECT 1655.6800 249.9400 1657.2800 250.4200 ;
        RECT 1716.2200 228.1800 1717.8200 228.6600 ;
        RECT 1716.2200 233.6200 1717.8200 234.1000 ;
        RECT 1700.6800 228.1800 1702.2800 228.6600 ;
        RECT 1700.6800 233.6200 1702.2800 234.1000 ;
        RECT 1716.2200 211.8600 1717.8200 212.3400 ;
        RECT 1716.2200 217.3000 1717.8200 217.7800 ;
        RECT 1716.2200 222.7400 1717.8200 223.2200 ;
        RECT 1700.6800 211.8600 1702.2800 212.3400 ;
        RECT 1700.6800 217.3000 1702.2800 217.7800 ;
        RECT 1700.6800 222.7400 1702.2800 223.2200 ;
        RECT 1716.2200 200.9800 1717.8200 201.4600 ;
        RECT 1716.2200 206.4200 1717.8200 206.9000 ;
        RECT 1700.6800 200.9800 1702.2800 201.4600 ;
        RECT 1700.6800 206.4200 1702.2800 206.9000 ;
        RECT 1700.6800 195.5400 1702.2800 196.0200 ;
        RECT 1716.2200 195.5400 1717.8200 196.0200 ;
        RECT 1655.6800 228.1800 1657.2800 228.6600 ;
        RECT 1655.6800 233.6200 1657.2800 234.1000 ;
        RECT 1655.6800 211.8600 1657.2800 212.3400 ;
        RECT 1655.6800 217.3000 1657.2800 217.7800 ;
        RECT 1655.6800 222.7400 1657.2800 223.2200 ;
        RECT 1655.6800 200.9800 1657.2800 201.4600 ;
        RECT 1655.6800 206.4200 1657.2800 206.9000 ;
        RECT 1655.6800 195.5400 1657.2800 196.0200 ;
        RECT 1610.6800 282.5800 1612.2800 283.0600 ;
        RECT 1610.6800 288.0200 1612.2800 288.5000 ;
        RECT 1610.6800 266.2600 1612.2800 266.7400 ;
        RECT 1610.6800 271.7000 1612.2800 272.1800 ;
        RECT 1610.6800 277.1400 1612.2800 277.6200 ;
        RECT 1565.6800 282.5800 1567.2800 283.0600 ;
        RECT 1565.6800 288.0200 1567.2800 288.5000 ;
        RECT 1565.6800 266.2600 1567.2800 266.7400 ;
        RECT 1565.6800 271.7000 1567.2800 272.1800 ;
        RECT 1565.6800 277.1400 1567.2800 277.6200 ;
        RECT 1610.6800 255.3800 1612.2800 255.8600 ;
        RECT 1610.6800 260.8200 1612.2800 261.3000 ;
        RECT 1610.6800 239.0600 1612.2800 239.5400 ;
        RECT 1610.6800 244.5000 1612.2800 244.9800 ;
        RECT 1610.6800 249.9400 1612.2800 250.4200 ;
        RECT 1565.6800 255.3800 1567.2800 255.8600 ;
        RECT 1565.6800 260.8200 1567.2800 261.3000 ;
        RECT 1565.6800 239.0600 1567.2800 239.5400 ;
        RECT 1565.6800 244.5000 1567.2800 244.9800 ;
        RECT 1565.6800 249.9400 1567.2800 250.4200 ;
        RECT 1520.6800 282.5800 1522.2800 283.0600 ;
        RECT 1520.6800 288.0200 1522.2800 288.5000 ;
        RECT 1513.5200 282.5800 1515.1200 283.0600 ;
        RECT 1513.5200 288.0200 1515.1200 288.5000 ;
        RECT 1520.6800 266.2600 1522.2800 266.7400 ;
        RECT 1520.6800 271.7000 1522.2800 272.1800 ;
        RECT 1520.6800 277.1400 1522.2800 277.6200 ;
        RECT 1513.5200 266.2600 1515.1200 266.7400 ;
        RECT 1513.5200 271.7000 1515.1200 272.1800 ;
        RECT 1513.5200 277.1400 1515.1200 277.6200 ;
        RECT 1520.6800 255.3800 1522.2800 255.8600 ;
        RECT 1520.6800 260.8200 1522.2800 261.3000 ;
        RECT 1513.5200 255.3800 1515.1200 255.8600 ;
        RECT 1513.5200 260.8200 1515.1200 261.3000 ;
        RECT 1520.6800 239.0600 1522.2800 239.5400 ;
        RECT 1520.6800 244.5000 1522.2800 244.9800 ;
        RECT 1520.6800 249.9400 1522.2800 250.4200 ;
        RECT 1513.5200 239.0600 1515.1200 239.5400 ;
        RECT 1513.5200 244.5000 1515.1200 244.9800 ;
        RECT 1513.5200 249.9400 1515.1200 250.4200 ;
        RECT 1610.6800 228.1800 1612.2800 228.6600 ;
        RECT 1610.6800 233.6200 1612.2800 234.1000 ;
        RECT 1610.6800 211.8600 1612.2800 212.3400 ;
        RECT 1610.6800 217.3000 1612.2800 217.7800 ;
        RECT 1610.6800 222.7400 1612.2800 223.2200 ;
        RECT 1565.6800 228.1800 1567.2800 228.6600 ;
        RECT 1565.6800 233.6200 1567.2800 234.1000 ;
        RECT 1565.6800 211.8600 1567.2800 212.3400 ;
        RECT 1565.6800 217.3000 1567.2800 217.7800 ;
        RECT 1565.6800 222.7400 1567.2800 223.2200 ;
        RECT 1610.6800 206.4200 1612.2800 206.9000 ;
        RECT 1610.6800 200.9800 1612.2800 201.4600 ;
        RECT 1610.6800 195.5400 1612.2800 196.0200 ;
        RECT 1565.6800 206.4200 1567.2800 206.9000 ;
        RECT 1565.6800 200.9800 1567.2800 201.4600 ;
        RECT 1565.6800 195.5400 1567.2800 196.0200 ;
        RECT 1520.6800 228.1800 1522.2800 228.6600 ;
        RECT 1520.6800 233.6200 1522.2800 234.1000 ;
        RECT 1513.5200 228.1800 1515.1200 228.6600 ;
        RECT 1513.5200 233.6200 1515.1200 234.1000 ;
        RECT 1520.6800 211.8600 1522.2800 212.3400 ;
        RECT 1520.6800 217.3000 1522.2800 217.7800 ;
        RECT 1520.6800 222.7400 1522.2800 223.2200 ;
        RECT 1513.5200 211.8600 1515.1200 212.3400 ;
        RECT 1513.5200 217.3000 1515.1200 217.7800 ;
        RECT 1513.5200 222.7400 1515.1200 223.2200 ;
        RECT 1520.6800 200.9800 1522.2800 201.4600 ;
        RECT 1520.6800 206.4200 1522.2800 206.9000 ;
        RECT 1513.5200 200.9800 1515.1200 201.4600 ;
        RECT 1513.5200 206.4200 1515.1200 206.9000 ;
        RECT 1513.5200 195.5400 1515.1200 196.0200 ;
        RECT 1520.6800 195.5400 1522.2800 196.0200 ;
        RECT 1510.5600 397.7300 1720.7800 399.3300 ;
        RECT 1510.5600 186.0300 1720.7800 187.6300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 183.2000 1515.1200 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 401.2400 1515.1200 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 183.2000 1717.8200 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 401.2400 1717.8200 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 186.0300 1512.1600 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 186.0300 1720.7800 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 397.7300 1512.1600 399.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 397.7300 1720.7800 399.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1513.6200 142.9400 1515.2200 173.2000 ;
        RECT 1716.1200 142.9400 1717.7200 173.2000 ;
      LAYER met3 ;
        RECT 1716.1200 163.4400 1717.7200 163.9200 ;
        RECT 1513.6200 163.4400 1515.2200 163.9200 ;
        RECT 1716.1200 152.5600 1717.7200 153.0400 ;
        RECT 1513.6200 152.5600 1515.2200 153.0400 ;
        RECT 1716.1200 158.0000 1717.7200 158.4800 ;
        RECT 1513.6200 158.0000 1515.2200 158.4800 ;
        RECT 1510.5600 168.8400 1720.7800 170.4400 ;
        RECT 1510.5600 144.5100 1720.7800 146.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.6200 142.9400 1515.2200 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.6200 171.6000 1515.2200 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.1200 142.9400 1717.7200 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.1200 171.6000 1717.7200 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 144.5100 1512.1600 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 144.5100 1720.7800 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 168.8400 1512.1600 170.4400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 168.8400 1720.7800 170.4400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 2252.7900 1702.2800 2466.0900 ;
        RECT 1655.6800 2252.7900 1657.2800 2466.0900 ;
        RECT 1610.6800 2252.7900 1612.2800 2466.0900 ;
        RECT 1565.6800 2252.7900 1567.2800 2466.0900 ;
        RECT 1520.6800 2252.7900 1522.2800 2466.0900 ;
        RECT 1716.2200 2249.9600 1717.8200 2469.6000 ;
        RECT 1513.5200 2249.9600 1515.1200 2469.6000 ;
      LAYER met3 ;
        RECT 1700.6800 2458.1400 1702.2800 2458.6200 ;
        RECT 1716.2200 2458.1400 1717.8200 2458.6200 ;
        RECT 1716.2200 2447.2600 1717.8200 2447.7400 ;
        RECT 1716.2200 2452.7000 1717.8200 2453.1800 ;
        RECT 1700.6800 2447.2600 1702.2800 2447.7400 ;
        RECT 1700.6800 2452.7000 1702.2800 2453.1800 ;
        RECT 1716.2200 2430.9400 1717.8200 2431.4200 ;
        RECT 1716.2200 2436.3800 1717.8200 2436.8600 ;
        RECT 1700.6800 2430.9400 1702.2800 2431.4200 ;
        RECT 1700.6800 2436.3800 1702.2800 2436.8600 ;
        RECT 1716.2200 2420.0600 1717.8200 2420.5400 ;
        RECT 1716.2200 2425.5000 1717.8200 2425.9800 ;
        RECT 1700.6800 2420.0600 1702.2800 2420.5400 ;
        RECT 1700.6800 2425.5000 1702.2800 2425.9800 ;
        RECT 1700.6800 2441.8200 1702.2800 2442.3000 ;
        RECT 1716.2200 2441.8200 1717.8200 2442.3000 ;
        RECT 1655.6800 2447.2600 1657.2800 2447.7400 ;
        RECT 1655.6800 2452.7000 1657.2800 2453.1800 ;
        RECT 1655.6800 2458.1400 1657.2800 2458.6200 ;
        RECT 1655.6800 2430.9400 1657.2800 2431.4200 ;
        RECT 1655.6800 2436.3800 1657.2800 2436.8600 ;
        RECT 1655.6800 2425.5000 1657.2800 2425.9800 ;
        RECT 1655.6800 2420.0600 1657.2800 2420.5400 ;
        RECT 1655.6800 2441.8200 1657.2800 2442.3000 ;
        RECT 1716.2200 2403.7400 1717.8200 2404.2200 ;
        RECT 1716.2200 2409.1800 1717.8200 2409.6600 ;
        RECT 1700.6800 2403.7400 1702.2800 2404.2200 ;
        RECT 1700.6800 2409.1800 1702.2800 2409.6600 ;
        RECT 1716.2200 2387.4200 1717.8200 2387.9000 ;
        RECT 1716.2200 2392.8600 1717.8200 2393.3400 ;
        RECT 1716.2200 2398.3000 1717.8200 2398.7800 ;
        RECT 1700.6800 2387.4200 1702.2800 2387.9000 ;
        RECT 1700.6800 2392.8600 1702.2800 2393.3400 ;
        RECT 1700.6800 2398.3000 1702.2800 2398.7800 ;
        RECT 1716.2200 2376.5400 1717.8200 2377.0200 ;
        RECT 1716.2200 2381.9800 1717.8200 2382.4600 ;
        RECT 1700.6800 2376.5400 1702.2800 2377.0200 ;
        RECT 1700.6800 2381.9800 1702.2800 2382.4600 ;
        RECT 1716.2200 2360.2200 1717.8200 2360.7000 ;
        RECT 1716.2200 2365.6600 1717.8200 2366.1400 ;
        RECT 1716.2200 2371.1000 1717.8200 2371.5800 ;
        RECT 1700.6800 2360.2200 1702.2800 2360.7000 ;
        RECT 1700.6800 2365.6600 1702.2800 2366.1400 ;
        RECT 1700.6800 2371.1000 1702.2800 2371.5800 ;
        RECT 1655.6800 2403.7400 1657.2800 2404.2200 ;
        RECT 1655.6800 2409.1800 1657.2800 2409.6600 ;
        RECT 1655.6800 2387.4200 1657.2800 2387.9000 ;
        RECT 1655.6800 2392.8600 1657.2800 2393.3400 ;
        RECT 1655.6800 2398.3000 1657.2800 2398.7800 ;
        RECT 1655.6800 2376.5400 1657.2800 2377.0200 ;
        RECT 1655.6800 2381.9800 1657.2800 2382.4600 ;
        RECT 1655.6800 2360.2200 1657.2800 2360.7000 ;
        RECT 1655.6800 2365.6600 1657.2800 2366.1400 ;
        RECT 1655.6800 2371.1000 1657.2800 2371.5800 ;
        RECT 1655.6800 2414.6200 1657.2800 2415.1000 ;
        RECT 1700.6800 2414.6200 1702.2800 2415.1000 ;
        RECT 1716.2200 2414.6200 1717.8200 2415.1000 ;
        RECT 1610.6800 2447.2600 1612.2800 2447.7400 ;
        RECT 1610.6800 2452.7000 1612.2800 2453.1800 ;
        RECT 1610.6800 2458.1400 1612.2800 2458.6200 ;
        RECT 1565.6800 2447.2600 1567.2800 2447.7400 ;
        RECT 1565.6800 2452.7000 1567.2800 2453.1800 ;
        RECT 1565.6800 2458.1400 1567.2800 2458.6200 ;
        RECT 1610.6800 2430.9400 1612.2800 2431.4200 ;
        RECT 1610.6800 2436.3800 1612.2800 2436.8600 ;
        RECT 1610.6800 2420.0600 1612.2800 2420.5400 ;
        RECT 1610.6800 2425.5000 1612.2800 2425.9800 ;
        RECT 1565.6800 2430.9400 1567.2800 2431.4200 ;
        RECT 1565.6800 2436.3800 1567.2800 2436.8600 ;
        RECT 1565.6800 2420.0600 1567.2800 2420.5400 ;
        RECT 1565.6800 2425.5000 1567.2800 2425.9800 ;
        RECT 1565.6800 2441.8200 1567.2800 2442.3000 ;
        RECT 1610.6800 2441.8200 1612.2800 2442.3000 ;
        RECT 1513.5200 2458.1400 1515.1200 2458.6200 ;
        RECT 1520.6800 2458.1400 1522.2800 2458.6200 ;
        RECT 1520.6800 2447.2600 1522.2800 2447.7400 ;
        RECT 1520.6800 2452.7000 1522.2800 2453.1800 ;
        RECT 1513.5200 2447.2600 1515.1200 2447.7400 ;
        RECT 1513.5200 2452.7000 1515.1200 2453.1800 ;
        RECT 1520.6800 2430.9400 1522.2800 2431.4200 ;
        RECT 1520.6800 2436.3800 1522.2800 2436.8600 ;
        RECT 1513.5200 2430.9400 1515.1200 2431.4200 ;
        RECT 1513.5200 2436.3800 1515.1200 2436.8600 ;
        RECT 1520.6800 2420.0600 1522.2800 2420.5400 ;
        RECT 1520.6800 2425.5000 1522.2800 2425.9800 ;
        RECT 1513.5200 2420.0600 1515.1200 2420.5400 ;
        RECT 1513.5200 2425.5000 1515.1200 2425.9800 ;
        RECT 1513.5200 2441.8200 1515.1200 2442.3000 ;
        RECT 1520.6800 2441.8200 1522.2800 2442.3000 ;
        RECT 1610.6800 2403.7400 1612.2800 2404.2200 ;
        RECT 1610.6800 2409.1800 1612.2800 2409.6600 ;
        RECT 1610.6800 2387.4200 1612.2800 2387.9000 ;
        RECT 1610.6800 2392.8600 1612.2800 2393.3400 ;
        RECT 1610.6800 2398.3000 1612.2800 2398.7800 ;
        RECT 1565.6800 2403.7400 1567.2800 2404.2200 ;
        RECT 1565.6800 2409.1800 1567.2800 2409.6600 ;
        RECT 1565.6800 2387.4200 1567.2800 2387.9000 ;
        RECT 1565.6800 2392.8600 1567.2800 2393.3400 ;
        RECT 1565.6800 2398.3000 1567.2800 2398.7800 ;
        RECT 1610.6800 2376.5400 1612.2800 2377.0200 ;
        RECT 1610.6800 2381.9800 1612.2800 2382.4600 ;
        RECT 1610.6800 2360.2200 1612.2800 2360.7000 ;
        RECT 1610.6800 2365.6600 1612.2800 2366.1400 ;
        RECT 1610.6800 2371.1000 1612.2800 2371.5800 ;
        RECT 1565.6800 2376.5400 1567.2800 2377.0200 ;
        RECT 1565.6800 2381.9800 1567.2800 2382.4600 ;
        RECT 1565.6800 2360.2200 1567.2800 2360.7000 ;
        RECT 1565.6800 2365.6600 1567.2800 2366.1400 ;
        RECT 1565.6800 2371.1000 1567.2800 2371.5800 ;
        RECT 1520.6800 2403.7400 1522.2800 2404.2200 ;
        RECT 1520.6800 2409.1800 1522.2800 2409.6600 ;
        RECT 1513.5200 2403.7400 1515.1200 2404.2200 ;
        RECT 1513.5200 2409.1800 1515.1200 2409.6600 ;
        RECT 1520.6800 2387.4200 1522.2800 2387.9000 ;
        RECT 1520.6800 2392.8600 1522.2800 2393.3400 ;
        RECT 1520.6800 2398.3000 1522.2800 2398.7800 ;
        RECT 1513.5200 2387.4200 1515.1200 2387.9000 ;
        RECT 1513.5200 2392.8600 1515.1200 2393.3400 ;
        RECT 1513.5200 2398.3000 1515.1200 2398.7800 ;
        RECT 1520.6800 2376.5400 1522.2800 2377.0200 ;
        RECT 1520.6800 2381.9800 1522.2800 2382.4600 ;
        RECT 1513.5200 2376.5400 1515.1200 2377.0200 ;
        RECT 1513.5200 2381.9800 1515.1200 2382.4600 ;
        RECT 1520.6800 2360.2200 1522.2800 2360.7000 ;
        RECT 1520.6800 2365.6600 1522.2800 2366.1400 ;
        RECT 1520.6800 2371.1000 1522.2800 2371.5800 ;
        RECT 1513.5200 2360.2200 1515.1200 2360.7000 ;
        RECT 1513.5200 2365.6600 1515.1200 2366.1400 ;
        RECT 1513.5200 2371.1000 1515.1200 2371.5800 ;
        RECT 1513.5200 2414.6200 1515.1200 2415.1000 ;
        RECT 1520.6800 2414.6200 1522.2800 2415.1000 ;
        RECT 1565.6800 2414.6200 1567.2800 2415.1000 ;
        RECT 1610.6800 2414.6200 1612.2800 2415.1000 ;
        RECT 1716.2200 2349.3400 1717.8200 2349.8200 ;
        RECT 1716.2200 2354.7800 1717.8200 2355.2600 ;
        RECT 1700.6800 2349.3400 1702.2800 2349.8200 ;
        RECT 1700.6800 2354.7800 1702.2800 2355.2600 ;
        RECT 1716.2200 2333.0200 1717.8200 2333.5000 ;
        RECT 1716.2200 2338.4600 1717.8200 2338.9400 ;
        RECT 1716.2200 2343.9000 1717.8200 2344.3800 ;
        RECT 1700.6800 2333.0200 1702.2800 2333.5000 ;
        RECT 1700.6800 2338.4600 1702.2800 2338.9400 ;
        RECT 1700.6800 2343.9000 1702.2800 2344.3800 ;
        RECT 1716.2200 2322.1400 1717.8200 2322.6200 ;
        RECT 1716.2200 2327.5800 1717.8200 2328.0600 ;
        RECT 1700.6800 2322.1400 1702.2800 2322.6200 ;
        RECT 1700.6800 2327.5800 1702.2800 2328.0600 ;
        RECT 1716.2200 2305.8200 1717.8200 2306.3000 ;
        RECT 1716.2200 2311.2600 1717.8200 2311.7400 ;
        RECT 1716.2200 2316.7000 1717.8200 2317.1800 ;
        RECT 1700.6800 2305.8200 1702.2800 2306.3000 ;
        RECT 1700.6800 2311.2600 1702.2800 2311.7400 ;
        RECT 1700.6800 2316.7000 1702.2800 2317.1800 ;
        RECT 1655.6800 2349.3400 1657.2800 2349.8200 ;
        RECT 1655.6800 2354.7800 1657.2800 2355.2600 ;
        RECT 1655.6800 2333.0200 1657.2800 2333.5000 ;
        RECT 1655.6800 2338.4600 1657.2800 2338.9400 ;
        RECT 1655.6800 2343.9000 1657.2800 2344.3800 ;
        RECT 1655.6800 2322.1400 1657.2800 2322.6200 ;
        RECT 1655.6800 2327.5800 1657.2800 2328.0600 ;
        RECT 1655.6800 2305.8200 1657.2800 2306.3000 ;
        RECT 1655.6800 2311.2600 1657.2800 2311.7400 ;
        RECT 1655.6800 2316.7000 1657.2800 2317.1800 ;
        RECT 1716.2200 2294.9400 1717.8200 2295.4200 ;
        RECT 1716.2200 2300.3800 1717.8200 2300.8600 ;
        RECT 1700.6800 2294.9400 1702.2800 2295.4200 ;
        RECT 1700.6800 2300.3800 1702.2800 2300.8600 ;
        RECT 1716.2200 2278.6200 1717.8200 2279.1000 ;
        RECT 1716.2200 2284.0600 1717.8200 2284.5400 ;
        RECT 1716.2200 2289.5000 1717.8200 2289.9800 ;
        RECT 1700.6800 2278.6200 1702.2800 2279.1000 ;
        RECT 1700.6800 2284.0600 1702.2800 2284.5400 ;
        RECT 1700.6800 2289.5000 1702.2800 2289.9800 ;
        RECT 1716.2200 2267.7400 1717.8200 2268.2200 ;
        RECT 1716.2200 2273.1800 1717.8200 2273.6600 ;
        RECT 1700.6800 2267.7400 1702.2800 2268.2200 ;
        RECT 1700.6800 2273.1800 1702.2800 2273.6600 ;
        RECT 1700.6800 2262.3000 1702.2800 2262.7800 ;
        RECT 1716.2200 2262.3000 1717.8200 2262.7800 ;
        RECT 1655.6800 2294.9400 1657.2800 2295.4200 ;
        RECT 1655.6800 2300.3800 1657.2800 2300.8600 ;
        RECT 1655.6800 2278.6200 1657.2800 2279.1000 ;
        RECT 1655.6800 2284.0600 1657.2800 2284.5400 ;
        RECT 1655.6800 2289.5000 1657.2800 2289.9800 ;
        RECT 1655.6800 2267.7400 1657.2800 2268.2200 ;
        RECT 1655.6800 2273.1800 1657.2800 2273.6600 ;
        RECT 1655.6800 2262.3000 1657.2800 2262.7800 ;
        RECT 1610.6800 2349.3400 1612.2800 2349.8200 ;
        RECT 1610.6800 2354.7800 1612.2800 2355.2600 ;
        RECT 1610.6800 2333.0200 1612.2800 2333.5000 ;
        RECT 1610.6800 2338.4600 1612.2800 2338.9400 ;
        RECT 1610.6800 2343.9000 1612.2800 2344.3800 ;
        RECT 1565.6800 2349.3400 1567.2800 2349.8200 ;
        RECT 1565.6800 2354.7800 1567.2800 2355.2600 ;
        RECT 1565.6800 2333.0200 1567.2800 2333.5000 ;
        RECT 1565.6800 2338.4600 1567.2800 2338.9400 ;
        RECT 1565.6800 2343.9000 1567.2800 2344.3800 ;
        RECT 1610.6800 2322.1400 1612.2800 2322.6200 ;
        RECT 1610.6800 2327.5800 1612.2800 2328.0600 ;
        RECT 1610.6800 2305.8200 1612.2800 2306.3000 ;
        RECT 1610.6800 2311.2600 1612.2800 2311.7400 ;
        RECT 1610.6800 2316.7000 1612.2800 2317.1800 ;
        RECT 1565.6800 2322.1400 1567.2800 2322.6200 ;
        RECT 1565.6800 2327.5800 1567.2800 2328.0600 ;
        RECT 1565.6800 2305.8200 1567.2800 2306.3000 ;
        RECT 1565.6800 2311.2600 1567.2800 2311.7400 ;
        RECT 1565.6800 2316.7000 1567.2800 2317.1800 ;
        RECT 1520.6800 2349.3400 1522.2800 2349.8200 ;
        RECT 1520.6800 2354.7800 1522.2800 2355.2600 ;
        RECT 1513.5200 2349.3400 1515.1200 2349.8200 ;
        RECT 1513.5200 2354.7800 1515.1200 2355.2600 ;
        RECT 1520.6800 2333.0200 1522.2800 2333.5000 ;
        RECT 1520.6800 2338.4600 1522.2800 2338.9400 ;
        RECT 1520.6800 2343.9000 1522.2800 2344.3800 ;
        RECT 1513.5200 2333.0200 1515.1200 2333.5000 ;
        RECT 1513.5200 2338.4600 1515.1200 2338.9400 ;
        RECT 1513.5200 2343.9000 1515.1200 2344.3800 ;
        RECT 1520.6800 2322.1400 1522.2800 2322.6200 ;
        RECT 1520.6800 2327.5800 1522.2800 2328.0600 ;
        RECT 1513.5200 2322.1400 1515.1200 2322.6200 ;
        RECT 1513.5200 2327.5800 1515.1200 2328.0600 ;
        RECT 1520.6800 2305.8200 1522.2800 2306.3000 ;
        RECT 1520.6800 2311.2600 1522.2800 2311.7400 ;
        RECT 1520.6800 2316.7000 1522.2800 2317.1800 ;
        RECT 1513.5200 2305.8200 1515.1200 2306.3000 ;
        RECT 1513.5200 2311.2600 1515.1200 2311.7400 ;
        RECT 1513.5200 2316.7000 1515.1200 2317.1800 ;
        RECT 1610.6800 2294.9400 1612.2800 2295.4200 ;
        RECT 1610.6800 2300.3800 1612.2800 2300.8600 ;
        RECT 1610.6800 2278.6200 1612.2800 2279.1000 ;
        RECT 1610.6800 2284.0600 1612.2800 2284.5400 ;
        RECT 1610.6800 2289.5000 1612.2800 2289.9800 ;
        RECT 1565.6800 2294.9400 1567.2800 2295.4200 ;
        RECT 1565.6800 2300.3800 1567.2800 2300.8600 ;
        RECT 1565.6800 2278.6200 1567.2800 2279.1000 ;
        RECT 1565.6800 2284.0600 1567.2800 2284.5400 ;
        RECT 1565.6800 2289.5000 1567.2800 2289.9800 ;
        RECT 1610.6800 2273.1800 1612.2800 2273.6600 ;
        RECT 1610.6800 2267.7400 1612.2800 2268.2200 ;
        RECT 1610.6800 2262.3000 1612.2800 2262.7800 ;
        RECT 1565.6800 2273.1800 1567.2800 2273.6600 ;
        RECT 1565.6800 2267.7400 1567.2800 2268.2200 ;
        RECT 1565.6800 2262.3000 1567.2800 2262.7800 ;
        RECT 1520.6800 2294.9400 1522.2800 2295.4200 ;
        RECT 1520.6800 2300.3800 1522.2800 2300.8600 ;
        RECT 1513.5200 2294.9400 1515.1200 2295.4200 ;
        RECT 1513.5200 2300.3800 1515.1200 2300.8600 ;
        RECT 1520.6800 2278.6200 1522.2800 2279.1000 ;
        RECT 1520.6800 2284.0600 1522.2800 2284.5400 ;
        RECT 1520.6800 2289.5000 1522.2800 2289.9800 ;
        RECT 1513.5200 2278.6200 1515.1200 2279.1000 ;
        RECT 1513.5200 2284.0600 1515.1200 2284.5400 ;
        RECT 1513.5200 2289.5000 1515.1200 2289.9800 ;
        RECT 1520.6800 2267.7400 1522.2800 2268.2200 ;
        RECT 1520.6800 2273.1800 1522.2800 2273.6600 ;
        RECT 1513.5200 2267.7400 1515.1200 2268.2200 ;
        RECT 1513.5200 2273.1800 1515.1200 2273.6600 ;
        RECT 1513.5200 2262.3000 1515.1200 2262.7800 ;
        RECT 1520.6800 2262.3000 1522.2800 2262.7800 ;
        RECT 1510.5600 2464.4900 1720.7800 2466.0900 ;
        RECT 1510.5600 2252.7900 1720.7800 2254.3900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 2249.9600 1515.1200 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 2468.0000 1515.1200 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 2249.9600 1717.8200 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 2468.0000 1717.8200 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2252.7900 1512.1600 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2252.7900 1720.7800 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2464.4900 1512.1600 2466.0900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2464.4900 1720.7800 2466.0900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 2023.1500 1702.2800 2236.4500 ;
        RECT 1655.6800 2023.1500 1657.2800 2236.4500 ;
        RECT 1610.6800 2023.1500 1612.2800 2236.4500 ;
        RECT 1565.6800 2023.1500 1567.2800 2236.4500 ;
        RECT 1520.6800 2023.1500 1522.2800 2236.4500 ;
        RECT 1716.2200 2020.3200 1717.8200 2239.9600 ;
        RECT 1513.5200 2020.3200 1515.1200 2239.9600 ;
      LAYER met3 ;
        RECT 1700.6800 2228.5000 1702.2800 2228.9800 ;
        RECT 1716.2200 2228.5000 1717.8200 2228.9800 ;
        RECT 1716.2200 2217.6200 1717.8200 2218.1000 ;
        RECT 1716.2200 2223.0600 1717.8200 2223.5400 ;
        RECT 1700.6800 2217.6200 1702.2800 2218.1000 ;
        RECT 1700.6800 2223.0600 1702.2800 2223.5400 ;
        RECT 1716.2200 2201.3000 1717.8200 2201.7800 ;
        RECT 1716.2200 2206.7400 1717.8200 2207.2200 ;
        RECT 1700.6800 2201.3000 1702.2800 2201.7800 ;
        RECT 1700.6800 2206.7400 1702.2800 2207.2200 ;
        RECT 1716.2200 2190.4200 1717.8200 2190.9000 ;
        RECT 1716.2200 2195.8600 1717.8200 2196.3400 ;
        RECT 1700.6800 2190.4200 1702.2800 2190.9000 ;
        RECT 1700.6800 2195.8600 1702.2800 2196.3400 ;
        RECT 1700.6800 2212.1800 1702.2800 2212.6600 ;
        RECT 1716.2200 2212.1800 1717.8200 2212.6600 ;
        RECT 1655.6800 2217.6200 1657.2800 2218.1000 ;
        RECT 1655.6800 2223.0600 1657.2800 2223.5400 ;
        RECT 1655.6800 2228.5000 1657.2800 2228.9800 ;
        RECT 1655.6800 2201.3000 1657.2800 2201.7800 ;
        RECT 1655.6800 2206.7400 1657.2800 2207.2200 ;
        RECT 1655.6800 2195.8600 1657.2800 2196.3400 ;
        RECT 1655.6800 2190.4200 1657.2800 2190.9000 ;
        RECT 1655.6800 2212.1800 1657.2800 2212.6600 ;
        RECT 1716.2200 2174.1000 1717.8200 2174.5800 ;
        RECT 1716.2200 2179.5400 1717.8200 2180.0200 ;
        RECT 1700.6800 2174.1000 1702.2800 2174.5800 ;
        RECT 1700.6800 2179.5400 1702.2800 2180.0200 ;
        RECT 1716.2200 2157.7800 1717.8200 2158.2600 ;
        RECT 1716.2200 2163.2200 1717.8200 2163.7000 ;
        RECT 1716.2200 2168.6600 1717.8200 2169.1400 ;
        RECT 1700.6800 2157.7800 1702.2800 2158.2600 ;
        RECT 1700.6800 2163.2200 1702.2800 2163.7000 ;
        RECT 1700.6800 2168.6600 1702.2800 2169.1400 ;
        RECT 1716.2200 2146.9000 1717.8200 2147.3800 ;
        RECT 1716.2200 2152.3400 1717.8200 2152.8200 ;
        RECT 1700.6800 2146.9000 1702.2800 2147.3800 ;
        RECT 1700.6800 2152.3400 1702.2800 2152.8200 ;
        RECT 1716.2200 2130.5800 1717.8200 2131.0600 ;
        RECT 1716.2200 2136.0200 1717.8200 2136.5000 ;
        RECT 1716.2200 2141.4600 1717.8200 2141.9400 ;
        RECT 1700.6800 2130.5800 1702.2800 2131.0600 ;
        RECT 1700.6800 2136.0200 1702.2800 2136.5000 ;
        RECT 1700.6800 2141.4600 1702.2800 2141.9400 ;
        RECT 1655.6800 2174.1000 1657.2800 2174.5800 ;
        RECT 1655.6800 2179.5400 1657.2800 2180.0200 ;
        RECT 1655.6800 2157.7800 1657.2800 2158.2600 ;
        RECT 1655.6800 2163.2200 1657.2800 2163.7000 ;
        RECT 1655.6800 2168.6600 1657.2800 2169.1400 ;
        RECT 1655.6800 2146.9000 1657.2800 2147.3800 ;
        RECT 1655.6800 2152.3400 1657.2800 2152.8200 ;
        RECT 1655.6800 2130.5800 1657.2800 2131.0600 ;
        RECT 1655.6800 2136.0200 1657.2800 2136.5000 ;
        RECT 1655.6800 2141.4600 1657.2800 2141.9400 ;
        RECT 1655.6800 2184.9800 1657.2800 2185.4600 ;
        RECT 1700.6800 2184.9800 1702.2800 2185.4600 ;
        RECT 1716.2200 2184.9800 1717.8200 2185.4600 ;
        RECT 1610.6800 2217.6200 1612.2800 2218.1000 ;
        RECT 1610.6800 2223.0600 1612.2800 2223.5400 ;
        RECT 1610.6800 2228.5000 1612.2800 2228.9800 ;
        RECT 1565.6800 2217.6200 1567.2800 2218.1000 ;
        RECT 1565.6800 2223.0600 1567.2800 2223.5400 ;
        RECT 1565.6800 2228.5000 1567.2800 2228.9800 ;
        RECT 1610.6800 2201.3000 1612.2800 2201.7800 ;
        RECT 1610.6800 2206.7400 1612.2800 2207.2200 ;
        RECT 1610.6800 2190.4200 1612.2800 2190.9000 ;
        RECT 1610.6800 2195.8600 1612.2800 2196.3400 ;
        RECT 1565.6800 2201.3000 1567.2800 2201.7800 ;
        RECT 1565.6800 2206.7400 1567.2800 2207.2200 ;
        RECT 1565.6800 2190.4200 1567.2800 2190.9000 ;
        RECT 1565.6800 2195.8600 1567.2800 2196.3400 ;
        RECT 1565.6800 2212.1800 1567.2800 2212.6600 ;
        RECT 1610.6800 2212.1800 1612.2800 2212.6600 ;
        RECT 1513.5200 2228.5000 1515.1200 2228.9800 ;
        RECT 1520.6800 2228.5000 1522.2800 2228.9800 ;
        RECT 1520.6800 2217.6200 1522.2800 2218.1000 ;
        RECT 1520.6800 2223.0600 1522.2800 2223.5400 ;
        RECT 1513.5200 2217.6200 1515.1200 2218.1000 ;
        RECT 1513.5200 2223.0600 1515.1200 2223.5400 ;
        RECT 1520.6800 2201.3000 1522.2800 2201.7800 ;
        RECT 1520.6800 2206.7400 1522.2800 2207.2200 ;
        RECT 1513.5200 2201.3000 1515.1200 2201.7800 ;
        RECT 1513.5200 2206.7400 1515.1200 2207.2200 ;
        RECT 1520.6800 2190.4200 1522.2800 2190.9000 ;
        RECT 1520.6800 2195.8600 1522.2800 2196.3400 ;
        RECT 1513.5200 2190.4200 1515.1200 2190.9000 ;
        RECT 1513.5200 2195.8600 1515.1200 2196.3400 ;
        RECT 1513.5200 2212.1800 1515.1200 2212.6600 ;
        RECT 1520.6800 2212.1800 1522.2800 2212.6600 ;
        RECT 1610.6800 2174.1000 1612.2800 2174.5800 ;
        RECT 1610.6800 2179.5400 1612.2800 2180.0200 ;
        RECT 1610.6800 2157.7800 1612.2800 2158.2600 ;
        RECT 1610.6800 2163.2200 1612.2800 2163.7000 ;
        RECT 1610.6800 2168.6600 1612.2800 2169.1400 ;
        RECT 1565.6800 2174.1000 1567.2800 2174.5800 ;
        RECT 1565.6800 2179.5400 1567.2800 2180.0200 ;
        RECT 1565.6800 2157.7800 1567.2800 2158.2600 ;
        RECT 1565.6800 2163.2200 1567.2800 2163.7000 ;
        RECT 1565.6800 2168.6600 1567.2800 2169.1400 ;
        RECT 1610.6800 2146.9000 1612.2800 2147.3800 ;
        RECT 1610.6800 2152.3400 1612.2800 2152.8200 ;
        RECT 1610.6800 2130.5800 1612.2800 2131.0600 ;
        RECT 1610.6800 2136.0200 1612.2800 2136.5000 ;
        RECT 1610.6800 2141.4600 1612.2800 2141.9400 ;
        RECT 1565.6800 2146.9000 1567.2800 2147.3800 ;
        RECT 1565.6800 2152.3400 1567.2800 2152.8200 ;
        RECT 1565.6800 2130.5800 1567.2800 2131.0600 ;
        RECT 1565.6800 2136.0200 1567.2800 2136.5000 ;
        RECT 1565.6800 2141.4600 1567.2800 2141.9400 ;
        RECT 1520.6800 2174.1000 1522.2800 2174.5800 ;
        RECT 1520.6800 2179.5400 1522.2800 2180.0200 ;
        RECT 1513.5200 2174.1000 1515.1200 2174.5800 ;
        RECT 1513.5200 2179.5400 1515.1200 2180.0200 ;
        RECT 1520.6800 2157.7800 1522.2800 2158.2600 ;
        RECT 1520.6800 2163.2200 1522.2800 2163.7000 ;
        RECT 1520.6800 2168.6600 1522.2800 2169.1400 ;
        RECT 1513.5200 2157.7800 1515.1200 2158.2600 ;
        RECT 1513.5200 2163.2200 1515.1200 2163.7000 ;
        RECT 1513.5200 2168.6600 1515.1200 2169.1400 ;
        RECT 1520.6800 2146.9000 1522.2800 2147.3800 ;
        RECT 1520.6800 2152.3400 1522.2800 2152.8200 ;
        RECT 1513.5200 2146.9000 1515.1200 2147.3800 ;
        RECT 1513.5200 2152.3400 1515.1200 2152.8200 ;
        RECT 1520.6800 2130.5800 1522.2800 2131.0600 ;
        RECT 1520.6800 2136.0200 1522.2800 2136.5000 ;
        RECT 1520.6800 2141.4600 1522.2800 2141.9400 ;
        RECT 1513.5200 2130.5800 1515.1200 2131.0600 ;
        RECT 1513.5200 2136.0200 1515.1200 2136.5000 ;
        RECT 1513.5200 2141.4600 1515.1200 2141.9400 ;
        RECT 1513.5200 2184.9800 1515.1200 2185.4600 ;
        RECT 1520.6800 2184.9800 1522.2800 2185.4600 ;
        RECT 1565.6800 2184.9800 1567.2800 2185.4600 ;
        RECT 1610.6800 2184.9800 1612.2800 2185.4600 ;
        RECT 1716.2200 2119.7000 1717.8200 2120.1800 ;
        RECT 1716.2200 2125.1400 1717.8200 2125.6200 ;
        RECT 1700.6800 2119.7000 1702.2800 2120.1800 ;
        RECT 1700.6800 2125.1400 1702.2800 2125.6200 ;
        RECT 1716.2200 2103.3800 1717.8200 2103.8600 ;
        RECT 1716.2200 2108.8200 1717.8200 2109.3000 ;
        RECT 1716.2200 2114.2600 1717.8200 2114.7400 ;
        RECT 1700.6800 2103.3800 1702.2800 2103.8600 ;
        RECT 1700.6800 2108.8200 1702.2800 2109.3000 ;
        RECT 1700.6800 2114.2600 1702.2800 2114.7400 ;
        RECT 1716.2200 2092.5000 1717.8200 2092.9800 ;
        RECT 1716.2200 2097.9400 1717.8200 2098.4200 ;
        RECT 1700.6800 2092.5000 1702.2800 2092.9800 ;
        RECT 1700.6800 2097.9400 1702.2800 2098.4200 ;
        RECT 1716.2200 2076.1800 1717.8200 2076.6600 ;
        RECT 1716.2200 2081.6200 1717.8200 2082.1000 ;
        RECT 1716.2200 2087.0600 1717.8200 2087.5400 ;
        RECT 1700.6800 2076.1800 1702.2800 2076.6600 ;
        RECT 1700.6800 2081.6200 1702.2800 2082.1000 ;
        RECT 1700.6800 2087.0600 1702.2800 2087.5400 ;
        RECT 1655.6800 2119.7000 1657.2800 2120.1800 ;
        RECT 1655.6800 2125.1400 1657.2800 2125.6200 ;
        RECT 1655.6800 2103.3800 1657.2800 2103.8600 ;
        RECT 1655.6800 2108.8200 1657.2800 2109.3000 ;
        RECT 1655.6800 2114.2600 1657.2800 2114.7400 ;
        RECT 1655.6800 2092.5000 1657.2800 2092.9800 ;
        RECT 1655.6800 2097.9400 1657.2800 2098.4200 ;
        RECT 1655.6800 2076.1800 1657.2800 2076.6600 ;
        RECT 1655.6800 2081.6200 1657.2800 2082.1000 ;
        RECT 1655.6800 2087.0600 1657.2800 2087.5400 ;
        RECT 1716.2200 2065.3000 1717.8200 2065.7800 ;
        RECT 1716.2200 2070.7400 1717.8200 2071.2200 ;
        RECT 1700.6800 2065.3000 1702.2800 2065.7800 ;
        RECT 1700.6800 2070.7400 1702.2800 2071.2200 ;
        RECT 1716.2200 2048.9800 1717.8200 2049.4600 ;
        RECT 1716.2200 2054.4200 1717.8200 2054.9000 ;
        RECT 1716.2200 2059.8600 1717.8200 2060.3400 ;
        RECT 1700.6800 2048.9800 1702.2800 2049.4600 ;
        RECT 1700.6800 2054.4200 1702.2800 2054.9000 ;
        RECT 1700.6800 2059.8600 1702.2800 2060.3400 ;
        RECT 1716.2200 2038.1000 1717.8200 2038.5800 ;
        RECT 1716.2200 2043.5400 1717.8200 2044.0200 ;
        RECT 1700.6800 2038.1000 1702.2800 2038.5800 ;
        RECT 1700.6800 2043.5400 1702.2800 2044.0200 ;
        RECT 1700.6800 2032.6600 1702.2800 2033.1400 ;
        RECT 1716.2200 2032.6600 1717.8200 2033.1400 ;
        RECT 1655.6800 2065.3000 1657.2800 2065.7800 ;
        RECT 1655.6800 2070.7400 1657.2800 2071.2200 ;
        RECT 1655.6800 2048.9800 1657.2800 2049.4600 ;
        RECT 1655.6800 2054.4200 1657.2800 2054.9000 ;
        RECT 1655.6800 2059.8600 1657.2800 2060.3400 ;
        RECT 1655.6800 2038.1000 1657.2800 2038.5800 ;
        RECT 1655.6800 2043.5400 1657.2800 2044.0200 ;
        RECT 1655.6800 2032.6600 1657.2800 2033.1400 ;
        RECT 1610.6800 2119.7000 1612.2800 2120.1800 ;
        RECT 1610.6800 2125.1400 1612.2800 2125.6200 ;
        RECT 1610.6800 2103.3800 1612.2800 2103.8600 ;
        RECT 1610.6800 2108.8200 1612.2800 2109.3000 ;
        RECT 1610.6800 2114.2600 1612.2800 2114.7400 ;
        RECT 1565.6800 2119.7000 1567.2800 2120.1800 ;
        RECT 1565.6800 2125.1400 1567.2800 2125.6200 ;
        RECT 1565.6800 2103.3800 1567.2800 2103.8600 ;
        RECT 1565.6800 2108.8200 1567.2800 2109.3000 ;
        RECT 1565.6800 2114.2600 1567.2800 2114.7400 ;
        RECT 1610.6800 2092.5000 1612.2800 2092.9800 ;
        RECT 1610.6800 2097.9400 1612.2800 2098.4200 ;
        RECT 1610.6800 2076.1800 1612.2800 2076.6600 ;
        RECT 1610.6800 2081.6200 1612.2800 2082.1000 ;
        RECT 1610.6800 2087.0600 1612.2800 2087.5400 ;
        RECT 1565.6800 2092.5000 1567.2800 2092.9800 ;
        RECT 1565.6800 2097.9400 1567.2800 2098.4200 ;
        RECT 1565.6800 2076.1800 1567.2800 2076.6600 ;
        RECT 1565.6800 2081.6200 1567.2800 2082.1000 ;
        RECT 1565.6800 2087.0600 1567.2800 2087.5400 ;
        RECT 1520.6800 2119.7000 1522.2800 2120.1800 ;
        RECT 1520.6800 2125.1400 1522.2800 2125.6200 ;
        RECT 1513.5200 2119.7000 1515.1200 2120.1800 ;
        RECT 1513.5200 2125.1400 1515.1200 2125.6200 ;
        RECT 1520.6800 2103.3800 1522.2800 2103.8600 ;
        RECT 1520.6800 2108.8200 1522.2800 2109.3000 ;
        RECT 1520.6800 2114.2600 1522.2800 2114.7400 ;
        RECT 1513.5200 2103.3800 1515.1200 2103.8600 ;
        RECT 1513.5200 2108.8200 1515.1200 2109.3000 ;
        RECT 1513.5200 2114.2600 1515.1200 2114.7400 ;
        RECT 1520.6800 2092.5000 1522.2800 2092.9800 ;
        RECT 1520.6800 2097.9400 1522.2800 2098.4200 ;
        RECT 1513.5200 2092.5000 1515.1200 2092.9800 ;
        RECT 1513.5200 2097.9400 1515.1200 2098.4200 ;
        RECT 1520.6800 2076.1800 1522.2800 2076.6600 ;
        RECT 1520.6800 2081.6200 1522.2800 2082.1000 ;
        RECT 1520.6800 2087.0600 1522.2800 2087.5400 ;
        RECT 1513.5200 2076.1800 1515.1200 2076.6600 ;
        RECT 1513.5200 2081.6200 1515.1200 2082.1000 ;
        RECT 1513.5200 2087.0600 1515.1200 2087.5400 ;
        RECT 1610.6800 2065.3000 1612.2800 2065.7800 ;
        RECT 1610.6800 2070.7400 1612.2800 2071.2200 ;
        RECT 1610.6800 2048.9800 1612.2800 2049.4600 ;
        RECT 1610.6800 2054.4200 1612.2800 2054.9000 ;
        RECT 1610.6800 2059.8600 1612.2800 2060.3400 ;
        RECT 1565.6800 2065.3000 1567.2800 2065.7800 ;
        RECT 1565.6800 2070.7400 1567.2800 2071.2200 ;
        RECT 1565.6800 2048.9800 1567.2800 2049.4600 ;
        RECT 1565.6800 2054.4200 1567.2800 2054.9000 ;
        RECT 1565.6800 2059.8600 1567.2800 2060.3400 ;
        RECT 1610.6800 2043.5400 1612.2800 2044.0200 ;
        RECT 1610.6800 2038.1000 1612.2800 2038.5800 ;
        RECT 1610.6800 2032.6600 1612.2800 2033.1400 ;
        RECT 1565.6800 2043.5400 1567.2800 2044.0200 ;
        RECT 1565.6800 2038.1000 1567.2800 2038.5800 ;
        RECT 1565.6800 2032.6600 1567.2800 2033.1400 ;
        RECT 1520.6800 2065.3000 1522.2800 2065.7800 ;
        RECT 1520.6800 2070.7400 1522.2800 2071.2200 ;
        RECT 1513.5200 2065.3000 1515.1200 2065.7800 ;
        RECT 1513.5200 2070.7400 1515.1200 2071.2200 ;
        RECT 1520.6800 2048.9800 1522.2800 2049.4600 ;
        RECT 1520.6800 2054.4200 1522.2800 2054.9000 ;
        RECT 1520.6800 2059.8600 1522.2800 2060.3400 ;
        RECT 1513.5200 2048.9800 1515.1200 2049.4600 ;
        RECT 1513.5200 2054.4200 1515.1200 2054.9000 ;
        RECT 1513.5200 2059.8600 1515.1200 2060.3400 ;
        RECT 1520.6800 2038.1000 1522.2800 2038.5800 ;
        RECT 1520.6800 2043.5400 1522.2800 2044.0200 ;
        RECT 1513.5200 2038.1000 1515.1200 2038.5800 ;
        RECT 1513.5200 2043.5400 1515.1200 2044.0200 ;
        RECT 1513.5200 2032.6600 1515.1200 2033.1400 ;
        RECT 1520.6800 2032.6600 1522.2800 2033.1400 ;
        RECT 1510.5600 2234.8500 1720.7800 2236.4500 ;
        RECT 1510.5600 2023.1500 1720.7800 2024.7500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 2020.3200 1515.1200 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 2238.3600 1515.1200 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 2020.3200 1717.8200 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 2238.3600 1717.8200 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2023.1500 1512.1600 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2023.1500 1720.7800 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2234.8500 1512.1600 2236.4500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2234.8500 1720.7800 2236.4500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 1793.5100 1702.2800 2006.8100 ;
        RECT 1655.6800 1793.5100 1657.2800 2006.8100 ;
        RECT 1610.6800 1793.5100 1612.2800 2006.8100 ;
        RECT 1565.6800 1793.5100 1567.2800 2006.8100 ;
        RECT 1520.6800 1793.5100 1522.2800 2006.8100 ;
        RECT 1716.2200 1790.6800 1717.8200 2010.3200 ;
        RECT 1513.5200 1790.6800 1515.1200 2010.3200 ;
      LAYER met3 ;
        RECT 1700.6800 1998.8600 1702.2800 1999.3400 ;
        RECT 1716.2200 1998.8600 1717.8200 1999.3400 ;
        RECT 1716.2200 1987.9800 1717.8200 1988.4600 ;
        RECT 1716.2200 1993.4200 1717.8200 1993.9000 ;
        RECT 1700.6800 1987.9800 1702.2800 1988.4600 ;
        RECT 1700.6800 1993.4200 1702.2800 1993.9000 ;
        RECT 1716.2200 1971.6600 1717.8200 1972.1400 ;
        RECT 1716.2200 1977.1000 1717.8200 1977.5800 ;
        RECT 1700.6800 1971.6600 1702.2800 1972.1400 ;
        RECT 1700.6800 1977.1000 1702.2800 1977.5800 ;
        RECT 1716.2200 1960.7800 1717.8200 1961.2600 ;
        RECT 1716.2200 1966.2200 1717.8200 1966.7000 ;
        RECT 1700.6800 1960.7800 1702.2800 1961.2600 ;
        RECT 1700.6800 1966.2200 1702.2800 1966.7000 ;
        RECT 1700.6800 1982.5400 1702.2800 1983.0200 ;
        RECT 1716.2200 1982.5400 1717.8200 1983.0200 ;
        RECT 1655.6800 1987.9800 1657.2800 1988.4600 ;
        RECT 1655.6800 1993.4200 1657.2800 1993.9000 ;
        RECT 1655.6800 1998.8600 1657.2800 1999.3400 ;
        RECT 1655.6800 1971.6600 1657.2800 1972.1400 ;
        RECT 1655.6800 1977.1000 1657.2800 1977.5800 ;
        RECT 1655.6800 1966.2200 1657.2800 1966.7000 ;
        RECT 1655.6800 1960.7800 1657.2800 1961.2600 ;
        RECT 1655.6800 1982.5400 1657.2800 1983.0200 ;
        RECT 1716.2200 1944.4600 1717.8200 1944.9400 ;
        RECT 1716.2200 1949.9000 1717.8200 1950.3800 ;
        RECT 1700.6800 1944.4600 1702.2800 1944.9400 ;
        RECT 1700.6800 1949.9000 1702.2800 1950.3800 ;
        RECT 1716.2200 1928.1400 1717.8200 1928.6200 ;
        RECT 1716.2200 1933.5800 1717.8200 1934.0600 ;
        RECT 1716.2200 1939.0200 1717.8200 1939.5000 ;
        RECT 1700.6800 1928.1400 1702.2800 1928.6200 ;
        RECT 1700.6800 1933.5800 1702.2800 1934.0600 ;
        RECT 1700.6800 1939.0200 1702.2800 1939.5000 ;
        RECT 1716.2200 1917.2600 1717.8200 1917.7400 ;
        RECT 1716.2200 1922.7000 1717.8200 1923.1800 ;
        RECT 1700.6800 1917.2600 1702.2800 1917.7400 ;
        RECT 1700.6800 1922.7000 1702.2800 1923.1800 ;
        RECT 1716.2200 1900.9400 1717.8200 1901.4200 ;
        RECT 1716.2200 1906.3800 1717.8200 1906.8600 ;
        RECT 1716.2200 1911.8200 1717.8200 1912.3000 ;
        RECT 1700.6800 1900.9400 1702.2800 1901.4200 ;
        RECT 1700.6800 1906.3800 1702.2800 1906.8600 ;
        RECT 1700.6800 1911.8200 1702.2800 1912.3000 ;
        RECT 1655.6800 1944.4600 1657.2800 1944.9400 ;
        RECT 1655.6800 1949.9000 1657.2800 1950.3800 ;
        RECT 1655.6800 1928.1400 1657.2800 1928.6200 ;
        RECT 1655.6800 1933.5800 1657.2800 1934.0600 ;
        RECT 1655.6800 1939.0200 1657.2800 1939.5000 ;
        RECT 1655.6800 1917.2600 1657.2800 1917.7400 ;
        RECT 1655.6800 1922.7000 1657.2800 1923.1800 ;
        RECT 1655.6800 1900.9400 1657.2800 1901.4200 ;
        RECT 1655.6800 1906.3800 1657.2800 1906.8600 ;
        RECT 1655.6800 1911.8200 1657.2800 1912.3000 ;
        RECT 1655.6800 1955.3400 1657.2800 1955.8200 ;
        RECT 1700.6800 1955.3400 1702.2800 1955.8200 ;
        RECT 1716.2200 1955.3400 1717.8200 1955.8200 ;
        RECT 1610.6800 1987.9800 1612.2800 1988.4600 ;
        RECT 1610.6800 1993.4200 1612.2800 1993.9000 ;
        RECT 1610.6800 1998.8600 1612.2800 1999.3400 ;
        RECT 1565.6800 1987.9800 1567.2800 1988.4600 ;
        RECT 1565.6800 1993.4200 1567.2800 1993.9000 ;
        RECT 1565.6800 1998.8600 1567.2800 1999.3400 ;
        RECT 1610.6800 1971.6600 1612.2800 1972.1400 ;
        RECT 1610.6800 1977.1000 1612.2800 1977.5800 ;
        RECT 1610.6800 1960.7800 1612.2800 1961.2600 ;
        RECT 1610.6800 1966.2200 1612.2800 1966.7000 ;
        RECT 1565.6800 1971.6600 1567.2800 1972.1400 ;
        RECT 1565.6800 1977.1000 1567.2800 1977.5800 ;
        RECT 1565.6800 1960.7800 1567.2800 1961.2600 ;
        RECT 1565.6800 1966.2200 1567.2800 1966.7000 ;
        RECT 1565.6800 1982.5400 1567.2800 1983.0200 ;
        RECT 1610.6800 1982.5400 1612.2800 1983.0200 ;
        RECT 1513.5200 1998.8600 1515.1200 1999.3400 ;
        RECT 1520.6800 1998.8600 1522.2800 1999.3400 ;
        RECT 1520.6800 1987.9800 1522.2800 1988.4600 ;
        RECT 1520.6800 1993.4200 1522.2800 1993.9000 ;
        RECT 1513.5200 1987.9800 1515.1200 1988.4600 ;
        RECT 1513.5200 1993.4200 1515.1200 1993.9000 ;
        RECT 1520.6800 1971.6600 1522.2800 1972.1400 ;
        RECT 1520.6800 1977.1000 1522.2800 1977.5800 ;
        RECT 1513.5200 1971.6600 1515.1200 1972.1400 ;
        RECT 1513.5200 1977.1000 1515.1200 1977.5800 ;
        RECT 1520.6800 1960.7800 1522.2800 1961.2600 ;
        RECT 1520.6800 1966.2200 1522.2800 1966.7000 ;
        RECT 1513.5200 1960.7800 1515.1200 1961.2600 ;
        RECT 1513.5200 1966.2200 1515.1200 1966.7000 ;
        RECT 1513.5200 1982.5400 1515.1200 1983.0200 ;
        RECT 1520.6800 1982.5400 1522.2800 1983.0200 ;
        RECT 1610.6800 1944.4600 1612.2800 1944.9400 ;
        RECT 1610.6800 1949.9000 1612.2800 1950.3800 ;
        RECT 1610.6800 1928.1400 1612.2800 1928.6200 ;
        RECT 1610.6800 1933.5800 1612.2800 1934.0600 ;
        RECT 1610.6800 1939.0200 1612.2800 1939.5000 ;
        RECT 1565.6800 1944.4600 1567.2800 1944.9400 ;
        RECT 1565.6800 1949.9000 1567.2800 1950.3800 ;
        RECT 1565.6800 1928.1400 1567.2800 1928.6200 ;
        RECT 1565.6800 1933.5800 1567.2800 1934.0600 ;
        RECT 1565.6800 1939.0200 1567.2800 1939.5000 ;
        RECT 1610.6800 1917.2600 1612.2800 1917.7400 ;
        RECT 1610.6800 1922.7000 1612.2800 1923.1800 ;
        RECT 1610.6800 1900.9400 1612.2800 1901.4200 ;
        RECT 1610.6800 1906.3800 1612.2800 1906.8600 ;
        RECT 1610.6800 1911.8200 1612.2800 1912.3000 ;
        RECT 1565.6800 1917.2600 1567.2800 1917.7400 ;
        RECT 1565.6800 1922.7000 1567.2800 1923.1800 ;
        RECT 1565.6800 1900.9400 1567.2800 1901.4200 ;
        RECT 1565.6800 1906.3800 1567.2800 1906.8600 ;
        RECT 1565.6800 1911.8200 1567.2800 1912.3000 ;
        RECT 1520.6800 1944.4600 1522.2800 1944.9400 ;
        RECT 1520.6800 1949.9000 1522.2800 1950.3800 ;
        RECT 1513.5200 1944.4600 1515.1200 1944.9400 ;
        RECT 1513.5200 1949.9000 1515.1200 1950.3800 ;
        RECT 1520.6800 1928.1400 1522.2800 1928.6200 ;
        RECT 1520.6800 1933.5800 1522.2800 1934.0600 ;
        RECT 1520.6800 1939.0200 1522.2800 1939.5000 ;
        RECT 1513.5200 1928.1400 1515.1200 1928.6200 ;
        RECT 1513.5200 1933.5800 1515.1200 1934.0600 ;
        RECT 1513.5200 1939.0200 1515.1200 1939.5000 ;
        RECT 1520.6800 1917.2600 1522.2800 1917.7400 ;
        RECT 1520.6800 1922.7000 1522.2800 1923.1800 ;
        RECT 1513.5200 1917.2600 1515.1200 1917.7400 ;
        RECT 1513.5200 1922.7000 1515.1200 1923.1800 ;
        RECT 1520.6800 1900.9400 1522.2800 1901.4200 ;
        RECT 1520.6800 1906.3800 1522.2800 1906.8600 ;
        RECT 1520.6800 1911.8200 1522.2800 1912.3000 ;
        RECT 1513.5200 1900.9400 1515.1200 1901.4200 ;
        RECT 1513.5200 1906.3800 1515.1200 1906.8600 ;
        RECT 1513.5200 1911.8200 1515.1200 1912.3000 ;
        RECT 1513.5200 1955.3400 1515.1200 1955.8200 ;
        RECT 1520.6800 1955.3400 1522.2800 1955.8200 ;
        RECT 1565.6800 1955.3400 1567.2800 1955.8200 ;
        RECT 1610.6800 1955.3400 1612.2800 1955.8200 ;
        RECT 1716.2200 1890.0600 1717.8200 1890.5400 ;
        RECT 1716.2200 1895.5000 1717.8200 1895.9800 ;
        RECT 1700.6800 1890.0600 1702.2800 1890.5400 ;
        RECT 1700.6800 1895.5000 1702.2800 1895.9800 ;
        RECT 1716.2200 1873.7400 1717.8200 1874.2200 ;
        RECT 1716.2200 1879.1800 1717.8200 1879.6600 ;
        RECT 1716.2200 1884.6200 1717.8200 1885.1000 ;
        RECT 1700.6800 1873.7400 1702.2800 1874.2200 ;
        RECT 1700.6800 1879.1800 1702.2800 1879.6600 ;
        RECT 1700.6800 1884.6200 1702.2800 1885.1000 ;
        RECT 1716.2200 1862.8600 1717.8200 1863.3400 ;
        RECT 1716.2200 1868.3000 1717.8200 1868.7800 ;
        RECT 1700.6800 1862.8600 1702.2800 1863.3400 ;
        RECT 1700.6800 1868.3000 1702.2800 1868.7800 ;
        RECT 1716.2200 1846.5400 1717.8200 1847.0200 ;
        RECT 1716.2200 1851.9800 1717.8200 1852.4600 ;
        RECT 1716.2200 1857.4200 1717.8200 1857.9000 ;
        RECT 1700.6800 1846.5400 1702.2800 1847.0200 ;
        RECT 1700.6800 1851.9800 1702.2800 1852.4600 ;
        RECT 1700.6800 1857.4200 1702.2800 1857.9000 ;
        RECT 1655.6800 1890.0600 1657.2800 1890.5400 ;
        RECT 1655.6800 1895.5000 1657.2800 1895.9800 ;
        RECT 1655.6800 1873.7400 1657.2800 1874.2200 ;
        RECT 1655.6800 1879.1800 1657.2800 1879.6600 ;
        RECT 1655.6800 1884.6200 1657.2800 1885.1000 ;
        RECT 1655.6800 1862.8600 1657.2800 1863.3400 ;
        RECT 1655.6800 1868.3000 1657.2800 1868.7800 ;
        RECT 1655.6800 1846.5400 1657.2800 1847.0200 ;
        RECT 1655.6800 1851.9800 1657.2800 1852.4600 ;
        RECT 1655.6800 1857.4200 1657.2800 1857.9000 ;
        RECT 1716.2200 1835.6600 1717.8200 1836.1400 ;
        RECT 1716.2200 1841.1000 1717.8200 1841.5800 ;
        RECT 1700.6800 1835.6600 1702.2800 1836.1400 ;
        RECT 1700.6800 1841.1000 1702.2800 1841.5800 ;
        RECT 1716.2200 1819.3400 1717.8200 1819.8200 ;
        RECT 1716.2200 1824.7800 1717.8200 1825.2600 ;
        RECT 1716.2200 1830.2200 1717.8200 1830.7000 ;
        RECT 1700.6800 1819.3400 1702.2800 1819.8200 ;
        RECT 1700.6800 1824.7800 1702.2800 1825.2600 ;
        RECT 1700.6800 1830.2200 1702.2800 1830.7000 ;
        RECT 1716.2200 1808.4600 1717.8200 1808.9400 ;
        RECT 1716.2200 1813.9000 1717.8200 1814.3800 ;
        RECT 1700.6800 1808.4600 1702.2800 1808.9400 ;
        RECT 1700.6800 1813.9000 1702.2800 1814.3800 ;
        RECT 1700.6800 1803.0200 1702.2800 1803.5000 ;
        RECT 1716.2200 1803.0200 1717.8200 1803.5000 ;
        RECT 1655.6800 1835.6600 1657.2800 1836.1400 ;
        RECT 1655.6800 1841.1000 1657.2800 1841.5800 ;
        RECT 1655.6800 1819.3400 1657.2800 1819.8200 ;
        RECT 1655.6800 1824.7800 1657.2800 1825.2600 ;
        RECT 1655.6800 1830.2200 1657.2800 1830.7000 ;
        RECT 1655.6800 1808.4600 1657.2800 1808.9400 ;
        RECT 1655.6800 1813.9000 1657.2800 1814.3800 ;
        RECT 1655.6800 1803.0200 1657.2800 1803.5000 ;
        RECT 1610.6800 1890.0600 1612.2800 1890.5400 ;
        RECT 1610.6800 1895.5000 1612.2800 1895.9800 ;
        RECT 1610.6800 1873.7400 1612.2800 1874.2200 ;
        RECT 1610.6800 1879.1800 1612.2800 1879.6600 ;
        RECT 1610.6800 1884.6200 1612.2800 1885.1000 ;
        RECT 1565.6800 1890.0600 1567.2800 1890.5400 ;
        RECT 1565.6800 1895.5000 1567.2800 1895.9800 ;
        RECT 1565.6800 1873.7400 1567.2800 1874.2200 ;
        RECT 1565.6800 1879.1800 1567.2800 1879.6600 ;
        RECT 1565.6800 1884.6200 1567.2800 1885.1000 ;
        RECT 1610.6800 1862.8600 1612.2800 1863.3400 ;
        RECT 1610.6800 1868.3000 1612.2800 1868.7800 ;
        RECT 1610.6800 1846.5400 1612.2800 1847.0200 ;
        RECT 1610.6800 1851.9800 1612.2800 1852.4600 ;
        RECT 1610.6800 1857.4200 1612.2800 1857.9000 ;
        RECT 1565.6800 1862.8600 1567.2800 1863.3400 ;
        RECT 1565.6800 1868.3000 1567.2800 1868.7800 ;
        RECT 1565.6800 1846.5400 1567.2800 1847.0200 ;
        RECT 1565.6800 1851.9800 1567.2800 1852.4600 ;
        RECT 1565.6800 1857.4200 1567.2800 1857.9000 ;
        RECT 1520.6800 1890.0600 1522.2800 1890.5400 ;
        RECT 1520.6800 1895.5000 1522.2800 1895.9800 ;
        RECT 1513.5200 1890.0600 1515.1200 1890.5400 ;
        RECT 1513.5200 1895.5000 1515.1200 1895.9800 ;
        RECT 1520.6800 1873.7400 1522.2800 1874.2200 ;
        RECT 1520.6800 1879.1800 1522.2800 1879.6600 ;
        RECT 1520.6800 1884.6200 1522.2800 1885.1000 ;
        RECT 1513.5200 1873.7400 1515.1200 1874.2200 ;
        RECT 1513.5200 1879.1800 1515.1200 1879.6600 ;
        RECT 1513.5200 1884.6200 1515.1200 1885.1000 ;
        RECT 1520.6800 1862.8600 1522.2800 1863.3400 ;
        RECT 1520.6800 1868.3000 1522.2800 1868.7800 ;
        RECT 1513.5200 1862.8600 1515.1200 1863.3400 ;
        RECT 1513.5200 1868.3000 1515.1200 1868.7800 ;
        RECT 1520.6800 1846.5400 1522.2800 1847.0200 ;
        RECT 1520.6800 1851.9800 1522.2800 1852.4600 ;
        RECT 1520.6800 1857.4200 1522.2800 1857.9000 ;
        RECT 1513.5200 1846.5400 1515.1200 1847.0200 ;
        RECT 1513.5200 1851.9800 1515.1200 1852.4600 ;
        RECT 1513.5200 1857.4200 1515.1200 1857.9000 ;
        RECT 1610.6800 1835.6600 1612.2800 1836.1400 ;
        RECT 1610.6800 1841.1000 1612.2800 1841.5800 ;
        RECT 1610.6800 1819.3400 1612.2800 1819.8200 ;
        RECT 1610.6800 1824.7800 1612.2800 1825.2600 ;
        RECT 1610.6800 1830.2200 1612.2800 1830.7000 ;
        RECT 1565.6800 1835.6600 1567.2800 1836.1400 ;
        RECT 1565.6800 1841.1000 1567.2800 1841.5800 ;
        RECT 1565.6800 1819.3400 1567.2800 1819.8200 ;
        RECT 1565.6800 1824.7800 1567.2800 1825.2600 ;
        RECT 1565.6800 1830.2200 1567.2800 1830.7000 ;
        RECT 1610.6800 1813.9000 1612.2800 1814.3800 ;
        RECT 1610.6800 1808.4600 1612.2800 1808.9400 ;
        RECT 1610.6800 1803.0200 1612.2800 1803.5000 ;
        RECT 1565.6800 1813.9000 1567.2800 1814.3800 ;
        RECT 1565.6800 1808.4600 1567.2800 1808.9400 ;
        RECT 1565.6800 1803.0200 1567.2800 1803.5000 ;
        RECT 1520.6800 1835.6600 1522.2800 1836.1400 ;
        RECT 1520.6800 1841.1000 1522.2800 1841.5800 ;
        RECT 1513.5200 1835.6600 1515.1200 1836.1400 ;
        RECT 1513.5200 1841.1000 1515.1200 1841.5800 ;
        RECT 1520.6800 1819.3400 1522.2800 1819.8200 ;
        RECT 1520.6800 1824.7800 1522.2800 1825.2600 ;
        RECT 1520.6800 1830.2200 1522.2800 1830.7000 ;
        RECT 1513.5200 1819.3400 1515.1200 1819.8200 ;
        RECT 1513.5200 1824.7800 1515.1200 1825.2600 ;
        RECT 1513.5200 1830.2200 1515.1200 1830.7000 ;
        RECT 1520.6800 1808.4600 1522.2800 1808.9400 ;
        RECT 1520.6800 1813.9000 1522.2800 1814.3800 ;
        RECT 1513.5200 1808.4600 1515.1200 1808.9400 ;
        RECT 1513.5200 1813.9000 1515.1200 1814.3800 ;
        RECT 1513.5200 1803.0200 1515.1200 1803.5000 ;
        RECT 1520.6800 1803.0200 1522.2800 1803.5000 ;
        RECT 1510.5600 2005.2100 1720.7800 2006.8100 ;
        RECT 1510.5600 1793.5100 1720.7800 1795.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1790.6800 1515.1200 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 2008.7200 1515.1200 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1790.6800 1717.8200 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 2008.7200 1717.8200 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1793.5100 1512.1600 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1793.5100 1720.7800 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2005.2100 1512.1600 2006.8100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2005.2100 1720.7800 2006.8100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 1563.8700 1702.2800 1777.1700 ;
        RECT 1655.6800 1563.8700 1657.2800 1777.1700 ;
        RECT 1610.6800 1563.8700 1612.2800 1777.1700 ;
        RECT 1565.6800 1563.8700 1567.2800 1777.1700 ;
        RECT 1520.6800 1563.8700 1522.2800 1777.1700 ;
        RECT 1716.2200 1561.0400 1717.8200 1780.6800 ;
        RECT 1513.5200 1561.0400 1515.1200 1780.6800 ;
      LAYER met3 ;
        RECT 1700.6800 1769.2200 1702.2800 1769.7000 ;
        RECT 1716.2200 1769.2200 1717.8200 1769.7000 ;
        RECT 1716.2200 1758.3400 1717.8200 1758.8200 ;
        RECT 1716.2200 1763.7800 1717.8200 1764.2600 ;
        RECT 1700.6800 1758.3400 1702.2800 1758.8200 ;
        RECT 1700.6800 1763.7800 1702.2800 1764.2600 ;
        RECT 1716.2200 1742.0200 1717.8200 1742.5000 ;
        RECT 1716.2200 1747.4600 1717.8200 1747.9400 ;
        RECT 1700.6800 1742.0200 1702.2800 1742.5000 ;
        RECT 1700.6800 1747.4600 1702.2800 1747.9400 ;
        RECT 1716.2200 1731.1400 1717.8200 1731.6200 ;
        RECT 1716.2200 1736.5800 1717.8200 1737.0600 ;
        RECT 1700.6800 1731.1400 1702.2800 1731.6200 ;
        RECT 1700.6800 1736.5800 1702.2800 1737.0600 ;
        RECT 1700.6800 1752.9000 1702.2800 1753.3800 ;
        RECT 1716.2200 1752.9000 1717.8200 1753.3800 ;
        RECT 1655.6800 1758.3400 1657.2800 1758.8200 ;
        RECT 1655.6800 1763.7800 1657.2800 1764.2600 ;
        RECT 1655.6800 1769.2200 1657.2800 1769.7000 ;
        RECT 1655.6800 1742.0200 1657.2800 1742.5000 ;
        RECT 1655.6800 1747.4600 1657.2800 1747.9400 ;
        RECT 1655.6800 1736.5800 1657.2800 1737.0600 ;
        RECT 1655.6800 1731.1400 1657.2800 1731.6200 ;
        RECT 1655.6800 1752.9000 1657.2800 1753.3800 ;
        RECT 1716.2200 1714.8200 1717.8200 1715.3000 ;
        RECT 1716.2200 1720.2600 1717.8200 1720.7400 ;
        RECT 1700.6800 1714.8200 1702.2800 1715.3000 ;
        RECT 1700.6800 1720.2600 1702.2800 1720.7400 ;
        RECT 1716.2200 1698.5000 1717.8200 1698.9800 ;
        RECT 1716.2200 1703.9400 1717.8200 1704.4200 ;
        RECT 1716.2200 1709.3800 1717.8200 1709.8600 ;
        RECT 1700.6800 1698.5000 1702.2800 1698.9800 ;
        RECT 1700.6800 1703.9400 1702.2800 1704.4200 ;
        RECT 1700.6800 1709.3800 1702.2800 1709.8600 ;
        RECT 1716.2200 1687.6200 1717.8200 1688.1000 ;
        RECT 1716.2200 1693.0600 1717.8200 1693.5400 ;
        RECT 1700.6800 1687.6200 1702.2800 1688.1000 ;
        RECT 1700.6800 1693.0600 1702.2800 1693.5400 ;
        RECT 1716.2200 1671.3000 1717.8200 1671.7800 ;
        RECT 1716.2200 1676.7400 1717.8200 1677.2200 ;
        RECT 1716.2200 1682.1800 1717.8200 1682.6600 ;
        RECT 1700.6800 1671.3000 1702.2800 1671.7800 ;
        RECT 1700.6800 1676.7400 1702.2800 1677.2200 ;
        RECT 1700.6800 1682.1800 1702.2800 1682.6600 ;
        RECT 1655.6800 1714.8200 1657.2800 1715.3000 ;
        RECT 1655.6800 1720.2600 1657.2800 1720.7400 ;
        RECT 1655.6800 1698.5000 1657.2800 1698.9800 ;
        RECT 1655.6800 1703.9400 1657.2800 1704.4200 ;
        RECT 1655.6800 1709.3800 1657.2800 1709.8600 ;
        RECT 1655.6800 1687.6200 1657.2800 1688.1000 ;
        RECT 1655.6800 1693.0600 1657.2800 1693.5400 ;
        RECT 1655.6800 1671.3000 1657.2800 1671.7800 ;
        RECT 1655.6800 1676.7400 1657.2800 1677.2200 ;
        RECT 1655.6800 1682.1800 1657.2800 1682.6600 ;
        RECT 1655.6800 1725.7000 1657.2800 1726.1800 ;
        RECT 1700.6800 1725.7000 1702.2800 1726.1800 ;
        RECT 1716.2200 1725.7000 1717.8200 1726.1800 ;
        RECT 1610.6800 1758.3400 1612.2800 1758.8200 ;
        RECT 1610.6800 1763.7800 1612.2800 1764.2600 ;
        RECT 1610.6800 1769.2200 1612.2800 1769.7000 ;
        RECT 1565.6800 1758.3400 1567.2800 1758.8200 ;
        RECT 1565.6800 1763.7800 1567.2800 1764.2600 ;
        RECT 1565.6800 1769.2200 1567.2800 1769.7000 ;
        RECT 1610.6800 1742.0200 1612.2800 1742.5000 ;
        RECT 1610.6800 1747.4600 1612.2800 1747.9400 ;
        RECT 1610.6800 1731.1400 1612.2800 1731.6200 ;
        RECT 1610.6800 1736.5800 1612.2800 1737.0600 ;
        RECT 1565.6800 1742.0200 1567.2800 1742.5000 ;
        RECT 1565.6800 1747.4600 1567.2800 1747.9400 ;
        RECT 1565.6800 1731.1400 1567.2800 1731.6200 ;
        RECT 1565.6800 1736.5800 1567.2800 1737.0600 ;
        RECT 1565.6800 1752.9000 1567.2800 1753.3800 ;
        RECT 1610.6800 1752.9000 1612.2800 1753.3800 ;
        RECT 1513.5200 1769.2200 1515.1200 1769.7000 ;
        RECT 1520.6800 1769.2200 1522.2800 1769.7000 ;
        RECT 1520.6800 1758.3400 1522.2800 1758.8200 ;
        RECT 1520.6800 1763.7800 1522.2800 1764.2600 ;
        RECT 1513.5200 1758.3400 1515.1200 1758.8200 ;
        RECT 1513.5200 1763.7800 1515.1200 1764.2600 ;
        RECT 1520.6800 1742.0200 1522.2800 1742.5000 ;
        RECT 1520.6800 1747.4600 1522.2800 1747.9400 ;
        RECT 1513.5200 1742.0200 1515.1200 1742.5000 ;
        RECT 1513.5200 1747.4600 1515.1200 1747.9400 ;
        RECT 1520.6800 1731.1400 1522.2800 1731.6200 ;
        RECT 1520.6800 1736.5800 1522.2800 1737.0600 ;
        RECT 1513.5200 1731.1400 1515.1200 1731.6200 ;
        RECT 1513.5200 1736.5800 1515.1200 1737.0600 ;
        RECT 1513.5200 1752.9000 1515.1200 1753.3800 ;
        RECT 1520.6800 1752.9000 1522.2800 1753.3800 ;
        RECT 1610.6800 1714.8200 1612.2800 1715.3000 ;
        RECT 1610.6800 1720.2600 1612.2800 1720.7400 ;
        RECT 1610.6800 1698.5000 1612.2800 1698.9800 ;
        RECT 1610.6800 1703.9400 1612.2800 1704.4200 ;
        RECT 1610.6800 1709.3800 1612.2800 1709.8600 ;
        RECT 1565.6800 1714.8200 1567.2800 1715.3000 ;
        RECT 1565.6800 1720.2600 1567.2800 1720.7400 ;
        RECT 1565.6800 1698.5000 1567.2800 1698.9800 ;
        RECT 1565.6800 1703.9400 1567.2800 1704.4200 ;
        RECT 1565.6800 1709.3800 1567.2800 1709.8600 ;
        RECT 1610.6800 1687.6200 1612.2800 1688.1000 ;
        RECT 1610.6800 1693.0600 1612.2800 1693.5400 ;
        RECT 1610.6800 1671.3000 1612.2800 1671.7800 ;
        RECT 1610.6800 1676.7400 1612.2800 1677.2200 ;
        RECT 1610.6800 1682.1800 1612.2800 1682.6600 ;
        RECT 1565.6800 1687.6200 1567.2800 1688.1000 ;
        RECT 1565.6800 1693.0600 1567.2800 1693.5400 ;
        RECT 1565.6800 1671.3000 1567.2800 1671.7800 ;
        RECT 1565.6800 1676.7400 1567.2800 1677.2200 ;
        RECT 1565.6800 1682.1800 1567.2800 1682.6600 ;
        RECT 1520.6800 1714.8200 1522.2800 1715.3000 ;
        RECT 1520.6800 1720.2600 1522.2800 1720.7400 ;
        RECT 1513.5200 1714.8200 1515.1200 1715.3000 ;
        RECT 1513.5200 1720.2600 1515.1200 1720.7400 ;
        RECT 1520.6800 1698.5000 1522.2800 1698.9800 ;
        RECT 1520.6800 1703.9400 1522.2800 1704.4200 ;
        RECT 1520.6800 1709.3800 1522.2800 1709.8600 ;
        RECT 1513.5200 1698.5000 1515.1200 1698.9800 ;
        RECT 1513.5200 1703.9400 1515.1200 1704.4200 ;
        RECT 1513.5200 1709.3800 1515.1200 1709.8600 ;
        RECT 1520.6800 1687.6200 1522.2800 1688.1000 ;
        RECT 1520.6800 1693.0600 1522.2800 1693.5400 ;
        RECT 1513.5200 1687.6200 1515.1200 1688.1000 ;
        RECT 1513.5200 1693.0600 1515.1200 1693.5400 ;
        RECT 1520.6800 1671.3000 1522.2800 1671.7800 ;
        RECT 1520.6800 1676.7400 1522.2800 1677.2200 ;
        RECT 1520.6800 1682.1800 1522.2800 1682.6600 ;
        RECT 1513.5200 1671.3000 1515.1200 1671.7800 ;
        RECT 1513.5200 1676.7400 1515.1200 1677.2200 ;
        RECT 1513.5200 1682.1800 1515.1200 1682.6600 ;
        RECT 1513.5200 1725.7000 1515.1200 1726.1800 ;
        RECT 1520.6800 1725.7000 1522.2800 1726.1800 ;
        RECT 1565.6800 1725.7000 1567.2800 1726.1800 ;
        RECT 1610.6800 1725.7000 1612.2800 1726.1800 ;
        RECT 1716.2200 1660.4200 1717.8200 1660.9000 ;
        RECT 1716.2200 1665.8600 1717.8200 1666.3400 ;
        RECT 1700.6800 1660.4200 1702.2800 1660.9000 ;
        RECT 1700.6800 1665.8600 1702.2800 1666.3400 ;
        RECT 1716.2200 1644.1000 1717.8200 1644.5800 ;
        RECT 1716.2200 1649.5400 1717.8200 1650.0200 ;
        RECT 1716.2200 1654.9800 1717.8200 1655.4600 ;
        RECT 1700.6800 1644.1000 1702.2800 1644.5800 ;
        RECT 1700.6800 1649.5400 1702.2800 1650.0200 ;
        RECT 1700.6800 1654.9800 1702.2800 1655.4600 ;
        RECT 1716.2200 1633.2200 1717.8200 1633.7000 ;
        RECT 1716.2200 1638.6600 1717.8200 1639.1400 ;
        RECT 1700.6800 1633.2200 1702.2800 1633.7000 ;
        RECT 1700.6800 1638.6600 1702.2800 1639.1400 ;
        RECT 1716.2200 1616.9000 1717.8200 1617.3800 ;
        RECT 1716.2200 1622.3400 1717.8200 1622.8200 ;
        RECT 1716.2200 1627.7800 1717.8200 1628.2600 ;
        RECT 1700.6800 1616.9000 1702.2800 1617.3800 ;
        RECT 1700.6800 1622.3400 1702.2800 1622.8200 ;
        RECT 1700.6800 1627.7800 1702.2800 1628.2600 ;
        RECT 1655.6800 1660.4200 1657.2800 1660.9000 ;
        RECT 1655.6800 1665.8600 1657.2800 1666.3400 ;
        RECT 1655.6800 1644.1000 1657.2800 1644.5800 ;
        RECT 1655.6800 1649.5400 1657.2800 1650.0200 ;
        RECT 1655.6800 1654.9800 1657.2800 1655.4600 ;
        RECT 1655.6800 1633.2200 1657.2800 1633.7000 ;
        RECT 1655.6800 1638.6600 1657.2800 1639.1400 ;
        RECT 1655.6800 1616.9000 1657.2800 1617.3800 ;
        RECT 1655.6800 1622.3400 1657.2800 1622.8200 ;
        RECT 1655.6800 1627.7800 1657.2800 1628.2600 ;
        RECT 1716.2200 1606.0200 1717.8200 1606.5000 ;
        RECT 1716.2200 1611.4600 1717.8200 1611.9400 ;
        RECT 1700.6800 1606.0200 1702.2800 1606.5000 ;
        RECT 1700.6800 1611.4600 1702.2800 1611.9400 ;
        RECT 1716.2200 1589.7000 1717.8200 1590.1800 ;
        RECT 1716.2200 1595.1400 1717.8200 1595.6200 ;
        RECT 1716.2200 1600.5800 1717.8200 1601.0600 ;
        RECT 1700.6800 1589.7000 1702.2800 1590.1800 ;
        RECT 1700.6800 1595.1400 1702.2800 1595.6200 ;
        RECT 1700.6800 1600.5800 1702.2800 1601.0600 ;
        RECT 1716.2200 1578.8200 1717.8200 1579.3000 ;
        RECT 1716.2200 1584.2600 1717.8200 1584.7400 ;
        RECT 1700.6800 1578.8200 1702.2800 1579.3000 ;
        RECT 1700.6800 1584.2600 1702.2800 1584.7400 ;
        RECT 1700.6800 1573.3800 1702.2800 1573.8600 ;
        RECT 1716.2200 1573.3800 1717.8200 1573.8600 ;
        RECT 1655.6800 1606.0200 1657.2800 1606.5000 ;
        RECT 1655.6800 1611.4600 1657.2800 1611.9400 ;
        RECT 1655.6800 1589.7000 1657.2800 1590.1800 ;
        RECT 1655.6800 1595.1400 1657.2800 1595.6200 ;
        RECT 1655.6800 1600.5800 1657.2800 1601.0600 ;
        RECT 1655.6800 1578.8200 1657.2800 1579.3000 ;
        RECT 1655.6800 1584.2600 1657.2800 1584.7400 ;
        RECT 1655.6800 1573.3800 1657.2800 1573.8600 ;
        RECT 1610.6800 1660.4200 1612.2800 1660.9000 ;
        RECT 1610.6800 1665.8600 1612.2800 1666.3400 ;
        RECT 1610.6800 1644.1000 1612.2800 1644.5800 ;
        RECT 1610.6800 1649.5400 1612.2800 1650.0200 ;
        RECT 1610.6800 1654.9800 1612.2800 1655.4600 ;
        RECT 1565.6800 1660.4200 1567.2800 1660.9000 ;
        RECT 1565.6800 1665.8600 1567.2800 1666.3400 ;
        RECT 1565.6800 1644.1000 1567.2800 1644.5800 ;
        RECT 1565.6800 1649.5400 1567.2800 1650.0200 ;
        RECT 1565.6800 1654.9800 1567.2800 1655.4600 ;
        RECT 1610.6800 1633.2200 1612.2800 1633.7000 ;
        RECT 1610.6800 1638.6600 1612.2800 1639.1400 ;
        RECT 1610.6800 1616.9000 1612.2800 1617.3800 ;
        RECT 1610.6800 1622.3400 1612.2800 1622.8200 ;
        RECT 1610.6800 1627.7800 1612.2800 1628.2600 ;
        RECT 1565.6800 1633.2200 1567.2800 1633.7000 ;
        RECT 1565.6800 1638.6600 1567.2800 1639.1400 ;
        RECT 1565.6800 1616.9000 1567.2800 1617.3800 ;
        RECT 1565.6800 1622.3400 1567.2800 1622.8200 ;
        RECT 1565.6800 1627.7800 1567.2800 1628.2600 ;
        RECT 1520.6800 1660.4200 1522.2800 1660.9000 ;
        RECT 1520.6800 1665.8600 1522.2800 1666.3400 ;
        RECT 1513.5200 1660.4200 1515.1200 1660.9000 ;
        RECT 1513.5200 1665.8600 1515.1200 1666.3400 ;
        RECT 1520.6800 1644.1000 1522.2800 1644.5800 ;
        RECT 1520.6800 1649.5400 1522.2800 1650.0200 ;
        RECT 1520.6800 1654.9800 1522.2800 1655.4600 ;
        RECT 1513.5200 1644.1000 1515.1200 1644.5800 ;
        RECT 1513.5200 1649.5400 1515.1200 1650.0200 ;
        RECT 1513.5200 1654.9800 1515.1200 1655.4600 ;
        RECT 1520.6800 1633.2200 1522.2800 1633.7000 ;
        RECT 1520.6800 1638.6600 1522.2800 1639.1400 ;
        RECT 1513.5200 1633.2200 1515.1200 1633.7000 ;
        RECT 1513.5200 1638.6600 1515.1200 1639.1400 ;
        RECT 1520.6800 1616.9000 1522.2800 1617.3800 ;
        RECT 1520.6800 1622.3400 1522.2800 1622.8200 ;
        RECT 1520.6800 1627.7800 1522.2800 1628.2600 ;
        RECT 1513.5200 1616.9000 1515.1200 1617.3800 ;
        RECT 1513.5200 1622.3400 1515.1200 1622.8200 ;
        RECT 1513.5200 1627.7800 1515.1200 1628.2600 ;
        RECT 1610.6800 1606.0200 1612.2800 1606.5000 ;
        RECT 1610.6800 1611.4600 1612.2800 1611.9400 ;
        RECT 1610.6800 1589.7000 1612.2800 1590.1800 ;
        RECT 1610.6800 1595.1400 1612.2800 1595.6200 ;
        RECT 1610.6800 1600.5800 1612.2800 1601.0600 ;
        RECT 1565.6800 1606.0200 1567.2800 1606.5000 ;
        RECT 1565.6800 1611.4600 1567.2800 1611.9400 ;
        RECT 1565.6800 1589.7000 1567.2800 1590.1800 ;
        RECT 1565.6800 1595.1400 1567.2800 1595.6200 ;
        RECT 1565.6800 1600.5800 1567.2800 1601.0600 ;
        RECT 1610.6800 1584.2600 1612.2800 1584.7400 ;
        RECT 1610.6800 1578.8200 1612.2800 1579.3000 ;
        RECT 1610.6800 1573.3800 1612.2800 1573.8600 ;
        RECT 1565.6800 1584.2600 1567.2800 1584.7400 ;
        RECT 1565.6800 1578.8200 1567.2800 1579.3000 ;
        RECT 1565.6800 1573.3800 1567.2800 1573.8600 ;
        RECT 1520.6800 1606.0200 1522.2800 1606.5000 ;
        RECT 1520.6800 1611.4600 1522.2800 1611.9400 ;
        RECT 1513.5200 1606.0200 1515.1200 1606.5000 ;
        RECT 1513.5200 1611.4600 1515.1200 1611.9400 ;
        RECT 1520.6800 1589.7000 1522.2800 1590.1800 ;
        RECT 1520.6800 1595.1400 1522.2800 1595.6200 ;
        RECT 1520.6800 1600.5800 1522.2800 1601.0600 ;
        RECT 1513.5200 1589.7000 1515.1200 1590.1800 ;
        RECT 1513.5200 1595.1400 1515.1200 1595.6200 ;
        RECT 1513.5200 1600.5800 1515.1200 1601.0600 ;
        RECT 1520.6800 1578.8200 1522.2800 1579.3000 ;
        RECT 1520.6800 1584.2600 1522.2800 1584.7400 ;
        RECT 1513.5200 1578.8200 1515.1200 1579.3000 ;
        RECT 1513.5200 1584.2600 1515.1200 1584.7400 ;
        RECT 1513.5200 1573.3800 1515.1200 1573.8600 ;
        RECT 1520.6800 1573.3800 1522.2800 1573.8600 ;
        RECT 1510.5600 1775.5700 1720.7800 1777.1700 ;
        RECT 1510.5600 1563.8700 1720.7800 1565.4700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1561.0400 1515.1200 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1779.0800 1515.1200 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1561.0400 1717.8200 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1779.0800 1717.8200 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1563.8700 1512.1600 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1563.8700 1720.7800 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1775.5700 1512.1600 1777.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1775.5700 1720.7800 1777.1700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 1334.2300 1702.2800 1547.5300 ;
        RECT 1655.6800 1334.2300 1657.2800 1547.5300 ;
        RECT 1610.6800 1334.2300 1612.2800 1547.5300 ;
        RECT 1565.6800 1334.2300 1567.2800 1547.5300 ;
        RECT 1520.6800 1334.2300 1522.2800 1547.5300 ;
        RECT 1716.2200 1331.4000 1717.8200 1551.0400 ;
        RECT 1513.5200 1331.4000 1515.1200 1551.0400 ;
      LAYER met3 ;
        RECT 1700.6800 1539.5800 1702.2800 1540.0600 ;
        RECT 1716.2200 1539.5800 1717.8200 1540.0600 ;
        RECT 1716.2200 1528.7000 1717.8200 1529.1800 ;
        RECT 1716.2200 1534.1400 1717.8200 1534.6200 ;
        RECT 1700.6800 1528.7000 1702.2800 1529.1800 ;
        RECT 1700.6800 1534.1400 1702.2800 1534.6200 ;
        RECT 1716.2200 1512.3800 1717.8200 1512.8600 ;
        RECT 1716.2200 1517.8200 1717.8200 1518.3000 ;
        RECT 1700.6800 1512.3800 1702.2800 1512.8600 ;
        RECT 1700.6800 1517.8200 1702.2800 1518.3000 ;
        RECT 1716.2200 1501.5000 1717.8200 1501.9800 ;
        RECT 1716.2200 1506.9400 1717.8200 1507.4200 ;
        RECT 1700.6800 1501.5000 1702.2800 1501.9800 ;
        RECT 1700.6800 1506.9400 1702.2800 1507.4200 ;
        RECT 1700.6800 1523.2600 1702.2800 1523.7400 ;
        RECT 1716.2200 1523.2600 1717.8200 1523.7400 ;
        RECT 1655.6800 1528.7000 1657.2800 1529.1800 ;
        RECT 1655.6800 1534.1400 1657.2800 1534.6200 ;
        RECT 1655.6800 1539.5800 1657.2800 1540.0600 ;
        RECT 1655.6800 1512.3800 1657.2800 1512.8600 ;
        RECT 1655.6800 1517.8200 1657.2800 1518.3000 ;
        RECT 1655.6800 1506.9400 1657.2800 1507.4200 ;
        RECT 1655.6800 1501.5000 1657.2800 1501.9800 ;
        RECT 1655.6800 1523.2600 1657.2800 1523.7400 ;
        RECT 1716.2200 1485.1800 1717.8200 1485.6600 ;
        RECT 1716.2200 1490.6200 1717.8200 1491.1000 ;
        RECT 1700.6800 1485.1800 1702.2800 1485.6600 ;
        RECT 1700.6800 1490.6200 1702.2800 1491.1000 ;
        RECT 1716.2200 1468.8600 1717.8200 1469.3400 ;
        RECT 1716.2200 1474.3000 1717.8200 1474.7800 ;
        RECT 1716.2200 1479.7400 1717.8200 1480.2200 ;
        RECT 1700.6800 1468.8600 1702.2800 1469.3400 ;
        RECT 1700.6800 1474.3000 1702.2800 1474.7800 ;
        RECT 1700.6800 1479.7400 1702.2800 1480.2200 ;
        RECT 1716.2200 1457.9800 1717.8200 1458.4600 ;
        RECT 1716.2200 1463.4200 1717.8200 1463.9000 ;
        RECT 1700.6800 1457.9800 1702.2800 1458.4600 ;
        RECT 1700.6800 1463.4200 1702.2800 1463.9000 ;
        RECT 1716.2200 1441.6600 1717.8200 1442.1400 ;
        RECT 1716.2200 1447.1000 1717.8200 1447.5800 ;
        RECT 1716.2200 1452.5400 1717.8200 1453.0200 ;
        RECT 1700.6800 1441.6600 1702.2800 1442.1400 ;
        RECT 1700.6800 1447.1000 1702.2800 1447.5800 ;
        RECT 1700.6800 1452.5400 1702.2800 1453.0200 ;
        RECT 1655.6800 1485.1800 1657.2800 1485.6600 ;
        RECT 1655.6800 1490.6200 1657.2800 1491.1000 ;
        RECT 1655.6800 1468.8600 1657.2800 1469.3400 ;
        RECT 1655.6800 1474.3000 1657.2800 1474.7800 ;
        RECT 1655.6800 1479.7400 1657.2800 1480.2200 ;
        RECT 1655.6800 1457.9800 1657.2800 1458.4600 ;
        RECT 1655.6800 1463.4200 1657.2800 1463.9000 ;
        RECT 1655.6800 1441.6600 1657.2800 1442.1400 ;
        RECT 1655.6800 1447.1000 1657.2800 1447.5800 ;
        RECT 1655.6800 1452.5400 1657.2800 1453.0200 ;
        RECT 1655.6800 1496.0600 1657.2800 1496.5400 ;
        RECT 1700.6800 1496.0600 1702.2800 1496.5400 ;
        RECT 1716.2200 1496.0600 1717.8200 1496.5400 ;
        RECT 1610.6800 1528.7000 1612.2800 1529.1800 ;
        RECT 1610.6800 1534.1400 1612.2800 1534.6200 ;
        RECT 1610.6800 1539.5800 1612.2800 1540.0600 ;
        RECT 1565.6800 1528.7000 1567.2800 1529.1800 ;
        RECT 1565.6800 1534.1400 1567.2800 1534.6200 ;
        RECT 1565.6800 1539.5800 1567.2800 1540.0600 ;
        RECT 1610.6800 1512.3800 1612.2800 1512.8600 ;
        RECT 1610.6800 1517.8200 1612.2800 1518.3000 ;
        RECT 1610.6800 1501.5000 1612.2800 1501.9800 ;
        RECT 1610.6800 1506.9400 1612.2800 1507.4200 ;
        RECT 1565.6800 1512.3800 1567.2800 1512.8600 ;
        RECT 1565.6800 1517.8200 1567.2800 1518.3000 ;
        RECT 1565.6800 1501.5000 1567.2800 1501.9800 ;
        RECT 1565.6800 1506.9400 1567.2800 1507.4200 ;
        RECT 1565.6800 1523.2600 1567.2800 1523.7400 ;
        RECT 1610.6800 1523.2600 1612.2800 1523.7400 ;
        RECT 1513.5200 1539.5800 1515.1200 1540.0600 ;
        RECT 1520.6800 1539.5800 1522.2800 1540.0600 ;
        RECT 1520.6800 1528.7000 1522.2800 1529.1800 ;
        RECT 1520.6800 1534.1400 1522.2800 1534.6200 ;
        RECT 1513.5200 1528.7000 1515.1200 1529.1800 ;
        RECT 1513.5200 1534.1400 1515.1200 1534.6200 ;
        RECT 1520.6800 1512.3800 1522.2800 1512.8600 ;
        RECT 1520.6800 1517.8200 1522.2800 1518.3000 ;
        RECT 1513.5200 1512.3800 1515.1200 1512.8600 ;
        RECT 1513.5200 1517.8200 1515.1200 1518.3000 ;
        RECT 1520.6800 1501.5000 1522.2800 1501.9800 ;
        RECT 1520.6800 1506.9400 1522.2800 1507.4200 ;
        RECT 1513.5200 1501.5000 1515.1200 1501.9800 ;
        RECT 1513.5200 1506.9400 1515.1200 1507.4200 ;
        RECT 1513.5200 1523.2600 1515.1200 1523.7400 ;
        RECT 1520.6800 1523.2600 1522.2800 1523.7400 ;
        RECT 1610.6800 1485.1800 1612.2800 1485.6600 ;
        RECT 1610.6800 1490.6200 1612.2800 1491.1000 ;
        RECT 1610.6800 1468.8600 1612.2800 1469.3400 ;
        RECT 1610.6800 1474.3000 1612.2800 1474.7800 ;
        RECT 1610.6800 1479.7400 1612.2800 1480.2200 ;
        RECT 1565.6800 1485.1800 1567.2800 1485.6600 ;
        RECT 1565.6800 1490.6200 1567.2800 1491.1000 ;
        RECT 1565.6800 1468.8600 1567.2800 1469.3400 ;
        RECT 1565.6800 1474.3000 1567.2800 1474.7800 ;
        RECT 1565.6800 1479.7400 1567.2800 1480.2200 ;
        RECT 1610.6800 1457.9800 1612.2800 1458.4600 ;
        RECT 1610.6800 1463.4200 1612.2800 1463.9000 ;
        RECT 1610.6800 1441.6600 1612.2800 1442.1400 ;
        RECT 1610.6800 1447.1000 1612.2800 1447.5800 ;
        RECT 1610.6800 1452.5400 1612.2800 1453.0200 ;
        RECT 1565.6800 1457.9800 1567.2800 1458.4600 ;
        RECT 1565.6800 1463.4200 1567.2800 1463.9000 ;
        RECT 1565.6800 1441.6600 1567.2800 1442.1400 ;
        RECT 1565.6800 1447.1000 1567.2800 1447.5800 ;
        RECT 1565.6800 1452.5400 1567.2800 1453.0200 ;
        RECT 1520.6800 1485.1800 1522.2800 1485.6600 ;
        RECT 1520.6800 1490.6200 1522.2800 1491.1000 ;
        RECT 1513.5200 1485.1800 1515.1200 1485.6600 ;
        RECT 1513.5200 1490.6200 1515.1200 1491.1000 ;
        RECT 1520.6800 1468.8600 1522.2800 1469.3400 ;
        RECT 1520.6800 1474.3000 1522.2800 1474.7800 ;
        RECT 1520.6800 1479.7400 1522.2800 1480.2200 ;
        RECT 1513.5200 1468.8600 1515.1200 1469.3400 ;
        RECT 1513.5200 1474.3000 1515.1200 1474.7800 ;
        RECT 1513.5200 1479.7400 1515.1200 1480.2200 ;
        RECT 1520.6800 1457.9800 1522.2800 1458.4600 ;
        RECT 1520.6800 1463.4200 1522.2800 1463.9000 ;
        RECT 1513.5200 1457.9800 1515.1200 1458.4600 ;
        RECT 1513.5200 1463.4200 1515.1200 1463.9000 ;
        RECT 1520.6800 1441.6600 1522.2800 1442.1400 ;
        RECT 1520.6800 1447.1000 1522.2800 1447.5800 ;
        RECT 1520.6800 1452.5400 1522.2800 1453.0200 ;
        RECT 1513.5200 1441.6600 1515.1200 1442.1400 ;
        RECT 1513.5200 1447.1000 1515.1200 1447.5800 ;
        RECT 1513.5200 1452.5400 1515.1200 1453.0200 ;
        RECT 1513.5200 1496.0600 1515.1200 1496.5400 ;
        RECT 1520.6800 1496.0600 1522.2800 1496.5400 ;
        RECT 1565.6800 1496.0600 1567.2800 1496.5400 ;
        RECT 1610.6800 1496.0600 1612.2800 1496.5400 ;
        RECT 1716.2200 1430.7800 1717.8200 1431.2600 ;
        RECT 1716.2200 1436.2200 1717.8200 1436.7000 ;
        RECT 1700.6800 1430.7800 1702.2800 1431.2600 ;
        RECT 1700.6800 1436.2200 1702.2800 1436.7000 ;
        RECT 1716.2200 1414.4600 1717.8200 1414.9400 ;
        RECT 1716.2200 1419.9000 1717.8200 1420.3800 ;
        RECT 1716.2200 1425.3400 1717.8200 1425.8200 ;
        RECT 1700.6800 1414.4600 1702.2800 1414.9400 ;
        RECT 1700.6800 1419.9000 1702.2800 1420.3800 ;
        RECT 1700.6800 1425.3400 1702.2800 1425.8200 ;
        RECT 1716.2200 1403.5800 1717.8200 1404.0600 ;
        RECT 1716.2200 1409.0200 1717.8200 1409.5000 ;
        RECT 1700.6800 1403.5800 1702.2800 1404.0600 ;
        RECT 1700.6800 1409.0200 1702.2800 1409.5000 ;
        RECT 1716.2200 1387.2600 1717.8200 1387.7400 ;
        RECT 1716.2200 1392.7000 1717.8200 1393.1800 ;
        RECT 1716.2200 1398.1400 1717.8200 1398.6200 ;
        RECT 1700.6800 1387.2600 1702.2800 1387.7400 ;
        RECT 1700.6800 1392.7000 1702.2800 1393.1800 ;
        RECT 1700.6800 1398.1400 1702.2800 1398.6200 ;
        RECT 1655.6800 1430.7800 1657.2800 1431.2600 ;
        RECT 1655.6800 1436.2200 1657.2800 1436.7000 ;
        RECT 1655.6800 1414.4600 1657.2800 1414.9400 ;
        RECT 1655.6800 1419.9000 1657.2800 1420.3800 ;
        RECT 1655.6800 1425.3400 1657.2800 1425.8200 ;
        RECT 1655.6800 1403.5800 1657.2800 1404.0600 ;
        RECT 1655.6800 1409.0200 1657.2800 1409.5000 ;
        RECT 1655.6800 1387.2600 1657.2800 1387.7400 ;
        RECT 1655.6800 1392.7000 1657.2800 1393.1800 ;
        RECT 1655.6800 1398.1400 1657.2800 1398.6200 ;
        RECT 1716.2200 1376.3800 1717.8200 1376.8600 ;
        RECT 1716.2200 1381.8200 1717.8200 1382.3000 ;
        RECT 1700.6800 1376.3800 1702.2800 1376.8600 ;
        RECT 1700.6800 1381.8200 1702.2800 1382.3000 ;
        RECT 1716.2200 1360.0600 1717.8200 1360.5400 ;
        RECT 1716.2200 1365.5000 1717.8200 1365.9800 ;
        RECT 1716.2200 1370.9400 1717.8200 1371.4200 ;
        RECT 1700.6800 1360.0600 1702.2800 1360.5400 ;
        RECT 1700.6800 1365.5000 1702.2800 1365.9800 ;
        RECT 1700.6800 1370.9400 1702.2800 1371.4200 ;
        RECT 1716.2200 1349.1800 1717.8200 1349.6600 ;
        RECT 1716.2200 1354.6200 1717.8200 1355.1000 ;
        RECT 1700.6800 1349.1800 1702.2800 1349.6600 ;
        RECT 1700.6800 1354.6200 1702.2800 1355.1000 ;
        RECT 1700.6800 1343.7400 1702.2800 1344.2200 ;
        RECT 1716.2200 1343.7400 1717.8200 1344.2200 ;
        RECT 1655.6800 1376.3800 1657.2800 1376.8600 ;
        RECT 1655.6800 1381.8200 1657.2800 1382.3000 ;
        RECT 1655.6800 1360.0600 1657.2800 1360.5400 ;
        RECT 1655.6800 1365.5000 1657.2800 1365.9800 ;
        RECT 1655.6800 1370.9400 1657.2800 1371.4200 ;
        RECT 1655.6800 1349.1800 1657.2800 1349.6600 ;
        RECT 1655.6800 1354.6200 1657.2800 1355.1000 ;
        RECT 1655.6800 1343.7400 1657.2800 1344.2200 ;
        RECT 1610.6800 1430.7800 1612.2800 1431.2600 ;
        RECT 1610.6800 1436.2200 1612.2800 1436.7000 ;
        RECT 1610.6800 1414.4600 1612.2800 1414.9400 ;
        RECT 1610.6800 1419.9000 1612.2800 1420.3800 ;
        RECT 1610.6800 1425.3400 1612.2800 1425.8200 ;
        RECT 1565.6800 1430.7800 1567.2800 1431.2600 ;
        RECT 1565.6800 1436.2200 1567.2800 1436.7000 ;
        RECT 1565.6800 1414.4600 1567.2800 1414.9400 ;
        RECT 1565.6800 1419.9000 1567.2800 1420.3800 ;
        RECT 1565.6800 1425.3400 1567.2800 1425.8200 ;
        RECT 1610.6800 1403.5800 1612.2800 1404.0600 ;
        RECT 1610.6800 1409.0200 1612.2800 1409.5000 ;
        RECT 1610.6800 1387.2600 1612.2800 1387.7400 ;
        RECT 1610.6800 1392.7000 1612.2800 1393.1800 ;
        RECT 1610.6800 1398.1400 1612.2800 1398.6200 ;
        RECT 1565.6800 1403.5800 1567.2800 1404.0600 ;
        RECT 1565.6800 1409.0200 1567.2800 1409.5000 ;
        RECT 1565.6800 1387.2600 1567.2800 1387.7400 ;
        RECT 1565.6800 1392.7000 1567.2800 1393.1800 ;
        RECT 1565.6800 1398.1400 1567.2800 1398.6200 ;
        RECT 1520.6800 1430.7800 1522.2800 1431.2600 ;
        RECT 1520.6800 1436.2200 1522.2800 1436.7000 ;
        RECT 1513.5200 1430.7800 1515.1200 1431.2600 ;
        RECT 1513.5200 1436.2200 1515.1200 1436.7000 ;
        RECT 1520.6800 1414.4600 1522.2800 1414.9400 ;
        RECT 1520.6800 1419.9000 1522.2800 1420.3800 ;
        RECT 1520.6800 1425.3400 1522.2800 1425.8200 ;
        RECT 1513.5200 1414.4600 1515.1200 1414.9400 ;
        RECT 1513.5200 1419.9000 1515.1200 1420.3800 ;
        RECT 1513.5200 1425.3400 1515.1200 1425.8200 ;
        RECT 1520.6800 1403.5800 1522.2800 1404.0600 ;
        RECT 1520.6800 1409.0200 1522.2800 1409.5000 ;
        RECT 1513.5200 1403.5800 1515.1200 1404.0600 ;
        RECT 1513.5200 1409.0200 1515.1200 1409.5000 ;
        RECT 1520.6800 1387.2600 1522.2800 1387.7400 ;
        RECT 1520.6800 1392.7000 1522.2800 1393.1800 ;
        RECT 1520.6800 1398.1400 1522.2800 1398.6200 ;
        RECT 1513.5200 1387.2600 1515.1200 1387.7400 ;
        RECT 1513.5200 1392.7000 1515.1200 1393.1800 ;
        RECT 1513.5200 1398.1400 1515.1200 1398.6200 ;
        RECT 1610.6800 1376.3800 1612.2800 1376.8600 ;
        RECT 1610.6800 1381.8200 1612.2800 1382.3000 ;
        RECT 1610.6800 1360.0600 1612.2800 1360.5400 ;
        RECT 1610.6800 1365.5000 1612.2800 1365.9800 ;
        RECT 1610.6800 1370.9400 1612.2800 1371.4200 ;
        RECT 1565.6800 1376.3800 1567.2800 1376.8600 ;
        RECT 1565.6800 1381.8200 1567.2800 1382.3000 ;
        RECT 1565.6800 1360.0600 1567.2800 1360.5400 ;
        RECT 1565.6800 1365.5000 1567.2800 1365.9800 ;
        RECT 1565.6800 1370.9400 1567.2800 1371.4200 ;
        RECT 1610.6800 1354.6200 1612.2800 1355.1000 ;
        RECT 1610.6800 1349.1800 1612.2800 1349.6600 ;
        RECT 1610.6800 1343.7400 1612.2800 1344.2200 ;
        RECT 1565.6800 1354.6200 1567.2800 1355.1000 ;
        RECT 1565.6800 1349.1800 1567.2800 1349.6600 ;
        RECT 1565.6800 1343.7400 1567.2800 1344.2200 ;
        RECT 1520.6800 1376.3800 1522.2800 1376.8600 ;
        RECT 1520.6800 1381.8200 1522.2800 1382.3000 ;
        RECT 1513.5200 1376.3800 1515.1200 1376.8600 ;
        RECT 1513.5200 1381.8200 1515.1200 1382.3000 ;
        RECT 1520.6800 1360.0600 1522.2800 1360.5400 ;
        RECT 1520.6800 1365.5000 1522.2800 1365.9800 ;
        RECT 1520.6800 1370.9400 1522.2800 1371.4200 ;
        RECT 1513.5200 1360.0600 1515.1200 1360.5400 ;
        RECT 1513.5200 1365.5000 1515.1200 1365.9800 ;
        RECT 1513.5200 1370.9400 1515.1200 1371.4200 ;
        RECT 1520.6800 1349.1800 1522.2800 1349.6600 ;
        RECT 1520.6800 1354.6200 1522.2800 1355.1000 ;
        RECT 1513.5200 1349.1800 1515.1200 1349.6600 ;
        RECT 1513.5200 1354.6200 1515.1200 1355.1000 ;
        RECT 1513.5200 1343.7400 1515.1200 1344.2200 ;
        RECT 1520.6800 1343.7400 1522.2800 1344.2200 ;
        RECT 1510.5600 1545.9300 1720.7800 1547.5300 ;
        RECT 1510.5600 1334.2300 1720.7800 1335.8300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1331.4000 1515.1200 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1549.4400 1515.1200 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1331.4000 1717.8200 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1549.4400 1717.8200 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1334.2300 1512.1600 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1334.2300 1720.7800 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1545.9300 1512.1600 1547.5300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1545.9300 1720.7800 1547.5300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 1104.5900 1702.2800 1317.8900 ;
        RECT 1655.6800 1104.5900 1657.2800 1317.8900 ;
        RECT 1610.6800 1104.5900 1612.2800 1317.8900 ;
        RECT 1565.6800 1104.5900 1567.2800 1317.8900 ;
        RECT 1520.6800 1104.5900 1522.2800 1317.8900 ;
        RECT 1716.2200 1101.7600 1717.8200 1321.4000 ;
        RECT 1513.5200 1101.7600 1515.1200 1321.4000 ;
      LAYER met3 ;
        RECT 1700.6800 1309.9400 1702.2800 1310.4200 ;
        RECT 1716.2200 1309.9400 1717.8200 1310.4200 ;
        RECT 1716.2200 1299.0600 1717.8200 1299.5400 ;
        RECT 1716.2200 1304.5000 1717.8200 1304.9800 ;
        RECT 1700.6800 1299.0600 1702.2800 1299.5400 ;
        RECT 1700.6800 1304.5000 1702.2800 1304.9800 ;
        RECT 1716.2200 1282.7400 1717.8200 1283.2200 ;
        RECT 1716.2200 1288.1800 1717.8200 1288.6600 ;
        RECT 1700.6800 1282.7400 1702.2800 1283.2200 ;
        RECT 1700.6800 1288.1800 1702.2800 1288.6600 ;
        RECT 1716.2200 1271.8600 1717.8200 1272.3400 ;
        RECT 1716.2200 1277.3000 1717.8200 1277.7800 ;
        RECT 1700.6800 1271.8600 1702.2800 1272.3400 ;
        RECT 1700.6800 1277.3000 1702.2800 1277.7800 ;
        RECT 1700.6800 1293.6200 1702.2800 1294.1000 ;
        RECT 1716.2200 1293.6200 1717.8200 1294.1000 ;
        RECT 1655.6800 1299.0600 1657.2800 1299.5400 ;
        RECT 1655.6800 1304.5000 1657.2800 1304.9800 ;
        RECT 1655.6800 1309.9400 1657.2800 1310.4200 ;
        RECT 1655.6800 1282.7400 1657.2800 1283.2200 ;
        RECT 1655.6800 1288.1800 1657.2800 1288.6600 ;
        RECT 1655.6800 1277.3000 1657.2800 1277.7800 ;
        RECT 1655.6800 1271.8600 1657.2800 1272.3400 ;
        RECT 1655.6800 1293.6200 1657.2800 1294.1000 ;
        RECT 1716.2200 1255.5400 1717.8200 1256.0200 ;
        RECT 1716.2200 1260.9800 1717.8200 1261.4600 ;
        RECT 1700.6800 1255.5400 1702.2800 1256.0200 ;
        RECT 1700.6800 1260.9800 1702.2800 1261.4600 ;
        RECT 1716.2200 1239.2200 1717.8200 1239.7000 ;
        RECT 1716.2200 1244.6600 1717.8200 1245.1400 ;
        RECT 1716.2200 1250.1000 1717.8200 1250.5800 ;
        RECT 1700.6800 1239.2200 1702.2800 1239.7000 ;
        RECT 1700.6800 1244.6600 1702.2800 1245.1400 ;
        RECT 1700.6800 1250.1000 1702.2800 1250.5800 ;
        RECT 1716.2200 1228.3400 1717.8200 1228.8200 ;
        RECT 1716.2200 1233.7800 1717.8200 1234.2600 ;
        RECT 1700.6800 1228.3400 1702.2800 1228.8200 ;
        RECT 1700.6800 1233.7800 1702.2800 1234.2600 ;
        RECT 1716.2200 1212.0200 1717.8200 1212.5000 ;
        RECT 1716.2200 1217.4600 1717.8200 1217.9400 ;
        RECT 1716.2200 1222.9000 1717.8200 1223.3800 ;
        RECT 1700.6800 1212.0200 1702.2800 1212.5000 ;
        RECT 1700.6800 1217.4600 1702.2800 1217.9400 ;
        RECT 1700.6800 1222.9000 1702.2800 1223.3800 ;
        RECT 1655.6800 1255.5400 1657.2800 1256.0200 ;
        RECT 1655.6800 1260.9800 1657.2800 1261.4600 ;
        RECT 1655.6800 1239.2200 1657.2800 1239.7000 ;
        RECT 1655.6800 1244.6600 1657.2800 1245.1400 ;
        RECT 1655.6800 1250.1000 1657.2800 1250.5800 ;
        RECT 1655.6800 1228.3400 1657.2800 1228.8200 ;
        RECT 1655.6800 1233.7800 1657.2800 1234.2600 ;
        RECT 1655.6800 1212.0200 1657.2800 1212.5000 ;
        RECT 1655.6800 1217.4600 1657.2800 1217.9400 ;
        RECT 1655.6800 1222.9000 1657.2800 1223.3800 ;
        RECT 1655.6800 1266.4200 1657.2800 1266.9000 ;
        RECT 1700.6800 1266.4200 1702.2800 1266.9000 ;
        RECT 1716.2200 1266.4200 1717.8200 1266.9000 ;
        RECT 1610.6800 1299.0600 1612.2800 1299.5400 ;
        RECT 1610.6800 1304.5000 1612.2800 1304.9800 ;
        RECT 1610.6800 1309.9400 1612.2800 1310.4200 ;
        RECT 1565.6800 1299.0600 1567.2800 1299.5400 ;
        RECT 1565.6800 1304.5000 1567.2800 1304.9800 ;
        RECT 1565.6800 1309.9400 1567.2800 1310.4200 ;
        RECT 1610.6800 1282.7400 1612.2800 1283.2200 ;
        RECT 1610.6800 1288.1800 1612.2800 1288.6600 ;
        RECT 1610.6800 1271.8600 1612.2800 1272.3400 ;
        RECT 1610.6800 1277.3000 1612.2800 1277.7800 ;
        RECT 1565.6800 1282.7400 1567.2800 1283.2200 ;
        RECT 1565.6800 1288.1800 1567.2800 1288.6600 ;
        RECT 1565.6800 1271.8600 1567.2800 1272.3400 ;
        RECT 1565.6800 1277.3000 1567.2800 1277.7800 ;
        RECT 1565.6800 1293.6200 1567.2800 1294.1000 ;
        RECT 1610.6800 1293.6200 1612.2800 1294.1000 ;
        RECT 1513.5200 1309.9400 1515.1200 1310.4200 ;
        RECT 1520.6800 1309.9400 1522.2800 1310.4200 ;
        RECT 1520.6800 1299.0600 1522.2800 1299.5400 ;
        RECT 1520.6800 1304.5000 1522.2800 1304.9800 ;
        RECT 1513.5200 1299.0600 1515.1200 1299.5400 ;
        RECT 1513.5200 1304.5000 1515.1200 1304.9800 ;
        RECT 1520.6800 1282.7400 1522.2800 1283.2200 ;
        RECT 1520.6800 1288.1800 1522.2800 1288.6600 ;
        RECT 1513.5200 1282.7400 1515.1200 1283.2200 ;
        RECT 1513.5200 1288.1800 1515.1200 1288.6600 ;
        RECT 1520.6800 1271.8600 1522.2800 1272.3400 ;
        RECT 1520.6800 1277.3000 1522.2800 1277.7800 ;
        RECT 1513.5200 1271.8600 1515.1200 1272.3400 ;
        RECT 1513.5200 1277.3000 1515.1200 1277.7800 ;
        RECT 1513.5200 1293.6200 1515.1200 1294.1000 ;
        RECT 1520.6800 1293.6200 1522.2800 1294.1000 ;
        RECT 1610.6800 1255.5400 1612.2800 1256.0200 ;
        RECT 1610.6800 1260.9800 1612.2800 1261.4600 ;
        RECT 1610.6800 1239.2200 1612.2800 1239.7000 ;
        RECT 1610.6800 1244.6600 1612.2800 1245.1400 ;
        RECT 1610.6800 1250.1000 1612.2800 1250.5800 ;
        RECT 1565.6800 1255.5400 1567.2800 1256.0200 ;
        RECT 1565.6800 1260.9800 1567.2800 1261.4600 ;
        RECT 1565.6800 1239.2200 1567.2800 1239.7000 ;
        RECT 1565.6800 1244.6600 1567.2800 1245.1400 ;
        RECT 1565.6800 1250.1000 1567.2800 1250.5800 ;
        RECT 1610.6800 1228.3400 1612.2800 1228.8200 ;
        RECT 1610.6800 1233.7800 1612.2800 1234.2600 ;
        RECT 1610.6800 1212.0200 1612.2800 1212.5000 ;
        RECT 1610.6800 1217.4600 1612.2800 1217.9400 ;
        RECT 1610.6800 1222.9000 1612.2800 1223.3800 ;
        RECT 1565.6800 1228.3400 1567.2800 1228.8200 ;
        RECT 1565.6800 1233.7800 1567.2800 1234.2600 ;
        RECT 1565.6800 1212.0200 1567.2800 1212.5000 ;
        RECT 1565.6800 1217.4600 1567.2800 1217.9400 ;
        RECT 1565.6800 1222.9000 1567.2800 1223.3800 ;
        RECT 1520.6800 1255.5400 1522.2800 1256.0200 ;
        RECT 1520.6800 1260.9800 1522.2800 1261.4600 ;
        RECT 1513.5200 1255.5400 1515.1200 1256.0200 ;
        RECT 1513.5200 1260.9800 1515.1200 1261.4600 ;
        RECT 1520.6800 1239.2200 1522.2800 1239.7000 ;
        RECT 1520.6800 1244.6600 1522.2800 1245.1400 ;
        RECT 1520.6800 1250.1000 1522.2800 1250.5800 ;
        RECT 1513.5200 1239.2200 1515.1200 1239.7000 ;
        RECT 1513.5200 1244.6600 1515.1200 1245.1400 ;
        RECT 1513.5200 1250.1000 1515.1200 1250.5800 ;
        RECT 1520.6800 1228.3400 1522.2800 1228.8200 ;
        RECT 1520.6800 1233.7800 1522.2800 1234.2600 ;
        RECT 1513.5200 1228.3400 1515.1200 1228.8200 ;
        RECT 1513.5200 1233.7800 1515.1200 1234.2600 ;
        RECT 1520.6800 1212.0200 1522.2800 1212.5000 ;
        RECT 1520.6800 1217.4600 1522.2800 1217.9400 ;
        RECT 1520.6800 1222.9000 1522.2800 1223.3800 ;
        RECT 1513.5200 1212.0200 1515.1200 1212.5000 ;
        RECT 1513.5200 1217.4600 1515.1200 1217.9400 ;
        RECT 1513.5200 1222.9000 1515.1200 1223.3800 ;
        RECT 1513.5200 1266.4200 1515.1200 1266.9000 ;
        RECT 1520.6800 1266.4200 1522.2800 1266.9000 ;
        RECT 1565.6800 1266.4200 1567.2800 1266.9000 ;
        RECT 1610.6800 1266.4200 1612.2800 1266.9000 ;
        RECT 1716.2200 1201.1400 1717.8200 1201.6200 ;
        RECT 1716.2200 1206.5800 1717.8200 1207.0600 ;
        RECT 1700.6800 1201.1400 1702.2800 1201.6200 ;
        RECT 1700.6800 1206.5800 1702.2800 1207.0600 ;
        RECT 1716.2200 1184.8200 1717.8200 1185.3000 ;
        RECT 1716.2200 1190.2600 1717.8200 1190.7400 ;
        RECT 1716.2200 1195.7000 1717.8200 1196.1800 ;
        RECT 1700.6800 1184.8200 1702.2800 1185.3000 ;
        RECT 1700.6800 1190.2600 1702.2800 1190.7400 ;
        RECT 1700.6800 1195.7000 1702.2800 1196.1800 ;
        RECT 1716.2200 1173.9400 1717.8200 1174.4200 ;
        RECT 1716.2200 1179.3800 1717.8200 1179.8600 ;
        RECT 1700.6800 1173.9400 1702.2800 1174.4200 ;
        RECT 1700.6800 1179.3800 1702.2800 1179.8600 ;
        RECT 1716.2200 1157.6200 1717.8200 1158.1000 ;
        RECT 1716.2200 1163.0600 1717.8200 1163.5400 ;
        RECT 1716.2200 1168.5000 1717.8200 1168.9800 ;
        RECT 1700.6800 1157.6200 1702.2800 1158.1000 ;
        RECT 1700.6800 1163.0600 1702.2800 1163.5400 ;
        RECT 1700.6800 1168.5000 1702.2800 1168.9800 ;
        RECT 1655.6800 1201.1400 1657.2800 1201.6200 ;
        RECT 1655.6800 1206.5800 1657.2800 1207.0600 ;
        RECT 1655.6800 1184.8200 1657.2800 1185.3000 ;
        RECT 1655.6800 1190.2600 1657.2800 1190.7400 ;
        RECT 1655.6800 1195.7000 1657.2800 1196.1800 ;
        RECT 1655.6800 1173.9400 1657.2800 1174.4200 ;
        RECT 1655.6800 1179.3800 1657.2800 1179.8600 ;
        RECT 1655.6800 1157.6200 1657.2800 1158.1000 ;
        RECT 1655.6800 1163.0600 1657.2800 1163.5400 ;
        RECT 1655.6800 1168.5000 1657.2800 1168.9800 ;
        RECT 1716.2200 1146.7400 1717.8200 1147.2200 ;
        RECT 1716.2200 1152.1800 1717.8200 1152.6600 ;
        RECT 1700.6800 1146.7400 1702.2800 1147.2200 ;
        RECT 1700.6800 1152.1800 1702.2800 1152.6600 ;
        RECT 1716.2200 1130.4200 1717.8200 1130.9000 ;
        RECT 1716.2200 1135.8600 1717.8200 1136.3400 ;
        RECT 1716.2200 1141.3000 1717.8200 1141.7800 ;
        RECT 1700.6800 1130.4200 1702.2800 1130.9000 ;
        RECT 1700.6800 1135.8600 1702.2800 1136.3400 ;
        RECT 1700.6800 1141.3000 1702.2800 1141.7800 ;
        RECT 1716.2200 1119.5400 1717.8200 1120.0200 ;
        RECT 1716.2200 1124.9800 1717.8200 1125.4600 ;
        RECT 1700.6800 1119.5400 1702.2800 1120.0200 ;
        RECT 1700.6800 1124.9800 1702.2800 1125.4600 ;
        RECT 1700.6800 1114.1000 1702.2800 1114.5800 ;
        RECT 1716.2200 1114.1000 1717.8200 1114.5800 ;
        RECT 1655.6800 1146.7400 1657.2800 1147.2200 ;
        RECT 1655.6800 1152.1800 1657.2800 1152.6600 ;
        RECT 1655.6800 1130.4200 1657.2800 1130.9000 ;
        RECT 1655.6800 1135.8600 1657.2800 1136.3400 ;
        RECT 1655.6800 1141.3000 1657.2800 1141.7800 ;
        RECT 1655.6800 1119.5400 1657.2800 1120.0200 ;
        RECT 1655.6800 1124.9800 1657.2800 1125.4600 ;
        RECT 1655.6800 1114.1000 1657.2800 1114.5800 ;
        RECT 1610.6800 1201.1400 1612.2800 1201.6200 ;
        RECT 1610.6800 1206.5800 1612.2800 1207.0600 ;
        RECT 1610.6800 1184.8200 1612.2800 1185.3000 ;
        RECT 1610.6800 1190.2600 1612.2800 1190.7400 ;
        RECT 1610.6800 1195.7000 1612.2800 1196.1800 ;
        RECT 1565.6800 1201.1400 1567.2800 1201.6200 ;
        RECT 1565.6800 1206.5800 1567.2800 1207.0600 ;
        RECT 1565.6800 1184.8200 1567.2800 1185.3000 ;
        RECT 1565.6800 1190.2600 1567.2800 1190.7400 ;
        RECT 1565.6800 1195.7000 1567.2800 1196.1800 ;
        RECT 1610.6800 1173.9400 1612.2800 1174.4200 ;
        RECT 1610.6800 1179.3800 1612.2800 1179.8600 ;
        RECT 1610.6800 1157.6200 1612.2800 1158.1000 ;
        RECT 1610.6800 1163.0600 1612.2800 1163.5400 ;
        RECT 1610.6800 1168.5000 1612.2800 1168.9800 ;
        RECT 1565.6800 1173.9400 1567.2800 1174.4200 ;
        RECT 1565.6800 1179.3800 1567.2800 1179.8600 ;
        RECT 1565.6800 1157.6200 1567.2800 1158.1000 ;
        RECT 1565.6800 1163.0600 1567.2800 1163.5400 ;
        RECT 1565.6800 1168.5000 1567.2800 1168.9800 ;
        RECT 1520.6800 1201.1400 1522.2800 1201.6200 ;
        RECT 1520.6800 1206.5800 1522.2800 1207.0600 ;
        RECT 1513.5200 1201.1400 1515.1200 1201.6200 ;
        RECT 1513.5200 1206.5800 1515.1200 1207.0600 ;
        RECT 1520.6800 1184.8200 1522.2800 1185.3000 ;
        RECT 1520.6800 1190.2600 1522.2800 1190.7400 ;
        RECT 1520.6800 1195.7000 1522.2800 1196.1800 ;
        RECT 1513.5200 1184.8200 1515.1200 1185.3000 ;
        RECT 1513.5200 1190.2600 1515.1200 1190.7400 ;
        RECT 1513.5200 1195.7000 1515.1200 1196.1800 ;
        RECT 1520.6800 1173.9400 1522.2800 1174.4200 ;
        RECT 1520.6800 1179.3800 1522.2800 1179.8600 ;
        RECT 1513.5200 1173.9400 1515.1200 1174.4200 ;
        RECT 1513.5200 1179.3800 1515.1200 1179.8600 ;
        RECT 1520.6800 1157.6200 1522.2800 1158.1000 ;
        RECT 1520.6800 1163.0600 1522.2800 1163.5400 ;
        RECT 1520.6800 1168.5000 1522.2800 1168.9800 ;
        RECT 1513.5200 1157.6200 1515.1200 1158.1000 ;
        RECT 1513.5200 1163.0600 1515.1200 1163.5400 ;
        RECT 1513.5200 1168.5000 1515.1200 1168.9800 ;
        RECT 1610.6800 1146.7400 1612.2800 1147.2200 ;
        RECT 1610.6800 1152.1800 1612.2800 1152.6600 ;
        RECT 1610.6800 1130.4200 1612.2800 1130.9000 ;
        RECT 1610.6800 1135.8600 1612.2800 1136.3400 ;
        RECT 1610.6800 1141.3000 1612.2800 1141.7800 ;
        RECT 1565.6800 1146.7400 1567.2800 1147.2200 ;
        RECT 1565.6800 1152.1800 1567.2800 1152.6600 ;
        RECT 1565.6800 1130.4200 1567.2800 1130.9000 ;
        RECT 1565.6800 1135.8600 1567.2800 1136.3400 ;
        RECT 1565.6800 1141.3000 1567.2800 1141.7800 ;
        RECT 1610.6800 1124.9800 1612.2800 1125.4600 ;
        RECT 1610.6800 1119.5400 1612.2800 1120.0200 ;
        RECT 1610.6800 1114.1000 1612.2800 1114.5800 ;
        RECT 1565.6800 1124.9800 1567.2800 1125.4600 ;
        RECT 1565.6800 1119.5400 1567.2800 1120.0200 ;
        RECT 1565.6800 1114.1000 1567.2800 1114.5800 ;
        RECT 1520.6800 1146.7400 1522.2800 1147.2200 ;
        RECT 1520.6800 1152.1800 1522.2800 1152.6600 ;
        RECT 1513.5200 1146.7400 1515.1200 1147.2200 ;
        RECT 1513.5200 1152.1800 1515.1200 1152.6600 ;
        RECT 1520.6800 1130.4200 1522.2800 1130.9000 ;
        RECT 1520.6800 1135.8600 1522.2800 1136.3400 ;
        RECT 1520.6800 1141.3000 1522.2800 1141.7800 ;
        RECT 1513.5200 1130.4200 1515.1200 1130.9000 ;
        RECT 1513.5200 1135.8600 1515.1200 1136.3400 ;
        RECT 1513.5200 1141.3000 1515.1200 1141.7800 ;
        RECT 1520.6800 1119.5400 1522.2800 1120.0200 ;
        RECT 1520.6800 1124.9800 1522.2800 1125.4600 ;
        RECT 1513.5200 1119.5400 1515.1200 1120.0200 ;
        RECT 1513.5200 1124.9800 1515.1200 1125.4600 ;
        RECT 1513.5200 1114.1000 1515.1200 1114.5800 ;
        RECT 1520.6800 1114.1000 1522.2800 1114.5800 ;
        RECT 1510.5600 1316.2900 1720.7800 1317.8900 ;
        RECT 1510.5600 1104.5900 1720.7800 1106.1900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1101.7600 1515.1200 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1319.8000 1515.1200 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1101.7600 1717.8200 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1319.8000 1717.8200 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1104.5900 1512.1600 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1104.5900 1720.7800 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1316.2900 1512.1600 1317.8900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1316.2900 1720.7800 1317.8900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 874.9500 1702.2800 1088.2500 ;
        RECT 1655.6800 874.9500 1657.2800 1088.2500 ;
        RECT 1610.6800 874.9500 1612.2800 1088.2500 ;
        RECT 1565.6800 874.9500 1567.2800 1088.2500 ;
        RECT 1520.6800 874.9500 1522.2800 1088.2500 ;
        RECT 1716.2200 872.1200 1717.8200 1091.7600 ;
        RECT 1513.5200 872.1200 1515.1200 1091.7600 ;
      LAYER met3 ;
        RECT 1700.6800 1080.3000 1702.2800 1080.7800 ;
        RECT 1716.2200 1080.3000 1717.8200 1080.7800 ;
        RECT 1716.2200 1069.4200 1717.8200 1069.9000 ;
        RECT 1716.2200 1074.8600 1717.8200 1075.3400 ;
        RECT 1700.6800 1069.4200 1702.2800 1069.9000 ;
        RECT 1700.6800 1074.8600 1702.2800 1075.3400 ;
        RECT 1716.2200 1053.1000 1717.8200 1053.5800 ;
        RECT 1716.2200 1058.5400 1717.8200 1059.0200 ;
        RECT 1700.6800 1053.1000 1702.2800 1053.5800 ;
        RECT 1700.6800 1058.5400 1702.2800 1059.0200 ;
        RECT 1716.2200 1042.2200 1717.8200 1042.7000 ;
        RECT 1716.2200 1047.6600 1717.8200 1048.1400 ;
        RECT 1700.6800 1042.2200 1702.2800 1042.7000 ;
        RECT 1700.6800 1047.6600 1702.2800 1048.1400 ;
        RECT 1700.6800 1063.9800 1702.2800 1064.4600 ;
        RECT 1716.2200 1063.9800 1717.8200 1064.4600 ;
        RECT 1655.6800 1069.4200 1657.2800 1069.9000 ;
        RECT 1655.6800 1074.8600 1657.2800 1075.3400 ;
        RECT 1655.6800 1080.3000 1657.2800 1080.7800 ;
        RECT 1655.6800 1053.1000 1657.2800 1053.5800 ;
        RECT 1655.6800 1058.5400 1657.2800 1059.0200 ;
        RECT 1655.6800 1047.6600 1657.2800 1048.1400 ;
        RECT 1655.6800 1042.2200 1657.2800 1042.7000 ;
        RECT 1655.6800 1063.9800 1657.2800 1064.4600 ;
        RECT 1716.2200 1025.9000 1717.8200 1026.3800 ;
        RECT 1716.2200 1031.3400 1717.8200 1031.8200 ;
        RECT 1700.6800 1025.9000 1702.2800 1026.3800 ;
        RECT 1700.6800 1031.3400 1702.2800 1031.8200 ;
        RECT 1716.2200 1009.5800 1717.8200 1010.0600 ;
        RECT 1716.2200 1015.0200 1717.8200 1015.5000 ;
        RECT 1716.2200 1020.4600 1717.8200 1020.9400 ;
        RECT 1700.6800 1009.5800 1702.2800 1010.0600 ;
        RECT 1700.6800 1015.0200 1702.2800 1015.5000 ;
        RECT 1700.6800 1020.4600 1702.2800 1020.9400 ;
        RECT 1716.2200 998.7000 1717.8200 999.1800 ;
        RECT 1716.2200 1004.1400 1717.8200 1004.6200 ;
        RECT 1700.6800 998.7000 1702.2800 999.1800 ;
        RECT 1700.6800 1004.1400 1702.2800 1004.6200 ;
        RECT 1716.2200 982.3800 1717.8200 982.8600 ;
        RECT 1716.2200 987.8200 1717.8200 988.3000 ;
        RECT 1716.2200 993.2600 1717.8200 993.7400 ;
        RECT 1700.6800 982.3800 1702.2800 982.8600 ;
        RECT 1700.6800 987.8200 1702.2800 988.3000 ;
        RECT 1700.6800 993.2600 1702.2800 993.7400 ;
        RECT 1655.6800 1025.9000 1657.2800 1026.3800 ;
        RECT 1655.6800 1031.3400 1657.2800 1031.8200 ;
        RECT 1655.6800 1009.5800 1657.2800 1010.0600 ;
        RECT 1655.6800 1015.0200 1657.2800 1015.5000 ;
        RECT 1655.6800 1020.4600 1657.2800 1020.9400 ;
        RECT 1655.6800 998.7000 1657.2800 999.1800 ;
        RECT 1655.6800 1004.1400 1657.2800 1004.6200 ;
        RECT 1655.6800 982.3800 1657.2800 982.8600 ;
        RECT 1655.6800 987.8200 1657.2800 988.3000 ;
        RECT 1655.6800 993.2600 1657.2800 993.7400 ;
        RECT 1655.6800 1036.7800 1657.2800 1037.2600 ;
        RECT 1700.6800 1036.7800 1702.2800 1037.2600 ;
        RECT 1716.2200 1036.7800 1717.8200 1037.2600 ;
        RECT 1610.6800 1069.4200 1612.2800 1069.9000 ;
        RECT 1610.6800 1074.8600 1612.2800 1075.3400 ;
        RECT 1610.6800 1080.3000 1612.2800 1080.7800 ;
        RECT 1565.6800 1069.4200 1567.2800 1069.9000 ;
        RECT 1565.6800 1074.8600 1567.2800 1075.3400 ;
        RECT 1565.6800 1080.3000 1567.2800 1080.7800 ;
        RECT 1610.6800 1053.1000 1612.2800 1053.5800 ;
        RECT 1610.6800 1058.5400 1612.2800 1059.0200 ;
        RECT 1610.6800 1042.2200 1612.2800 1042.7000 ;
        RECT 1610.6800 1047.6600 1612.2800 1048.1400 ;
        RECT 1565.6800 1053.1000 1567.2800 1053.5800 ;
        RECT 1565.6800 1058.5400 1567.2800 1059.0200 ;
        RECT 1565.6800 1042.2200 1567.2800 1042.7000 ;
        RECT 1565.6800 1047.6600 1567.2800 1048.1400 ;
        RECT 1565.6800 1063.9800 1567.2800 1064.4600 ;
        RECT 1610.6800 1063.9800 1612.2800 1064.4600 ;
        RECT 1513.5200 1080.3000 1515.1200 1080.7800 ;
        RECT 1520.6800 1080.3000 1522.2800 1080.7800 ;
        RECT 1520.6800 1069.4200 1522.2800 1069.9000 ;
        RECT 1520.6800 1074.8600 1522.2800 1075.3400 ;
        RECT 1513.5200 1069.4200 1515.1200 1069.9000 ;
        RECT 1513.5200 1074.8600 1515.1200 1075.3400 ;
        RECT 1520.6800 1053.1000 1522.2800 1053.5800 ;
        RECT 1520.6800 1058.5400 1522.2800 1059.0200 ;
        RECT 1513.5200 1053.1000 1515.1200 1053.5800 ;
        RECT 1513.5200 1058.5400 1515.1200 1059.0200 ;
        RECT 1520.6800 1042.2200 1522.2800 1042.7000 ;
        RECT 1520.6800 1047.6600 1522.2800 1048.1400 ;
        RECT 1513.5200 1042.2200 1515.1200 1042.7000 ;
        RECT 1513.5200 1047.6600 1515.1200 1048.1400 ;
        RECT 1513.5200 1063.9800 1515.1200 1064.4600 ;
        RECT 1520.6800 1063.9800 1522.2800 1064.4600 ;
        RECT 1610.6800 1025.9000 1612.2800 1026.3800 ;
        RECT 1610.6800 1031.3400 1612.2800 1031.8200 ;
        RECT 1610.6800 1009.5800 1612.2800 1010.0600 ;
        RECT 1610.6800 1015.0200 1612.2800 1015.5000 ;
        RECT 1610.6800 1020.4600 1612.2800 1020.9400 ;
        RECT 1565.6800 1025.9000 1567.2800 1026.3800 ;
        RECT 1565.6800 1031.3400 1567.2800 1031.8200 ;
        RECT 1565.6800 1009.5800 1567.2800 1010.0600 ;
        RECT 1565.6800 1015.0200 1567.2800 1015.5000 ;
        RECT 1565.6800 1020.4600 1567.2800 1020.9400 ;
        RECT 1610.6800 998.7000 1612.2800 999.1800 ;
        RECT 1610.6800 1004.1400 1612.2800 1004.6200 ;
        RECT 1610.6800 982.3800 1612.2800 982.8600 ;
        RECT 1610.6800 987.8200 1612.2800 988.3000 ;
        RECT 1610.6800 993.2600 1612.2800 993.7400 ;
        RECT 1565.6800 998.7000 1567.2800 999.1800 ;
        RECT 1565.6800 1004.1400 1567.2800 1004.6200 ;
        RECT 1565.6800 982.3800 1567.2800 982.8600 ;
        RECT 1565.6800 987.8200 1567.2800 988.3000 ;
        RECT 1565.6800 993.2600 1567.2800 993.7400 ;
        RECT 1520.6800 1025.9000 1522.2800 1026.3800 ;
        RECT 1520.6800 1031.3400 1522.2800 1031.8200 ;
        RECT 1513.5200 1025.9000 1515.1200 1026.3800 ;
        RECT 1513.5200 1031.3400 1515.1200 1031.8200 ;
        RECT 1520.6800 1009.5800 1522.2800 1010.0600 ;
        RECT 1520.6800 1015.0200 1522.2800 1015.5000 ;
        RECT 1520.6800 1020.4600 1522.2800 1020.9400 ;
        RECT 1513.5200 1009.5800 1515.1200 1010.0600 ;
        RECT 1513.5200 1015.0200 1515.1200 1015.5000 ;
        RECT 1513.5200 1020.4600 1515.1200 1020.9400 ;
        RECT 1520.6800 998.7000 1522.2800 999.1800 ;
        RECT 1520.6800 1004.1400 1522.2800 1004.6200 ;
        RECT 1513.5200 998.7000 1515.1200 999.1800 ;
        RECT 1513.5200 1004.1400 1515.1200 1004.6200 ;
        RECT 1520.6800 982.3800 1522.2800 982.8600 ;
        RECT 1520.6800 987.8200 1522.2800 988.3000 ;
        RECT 1520.6800 993.2600 1522.2800 993.7400 ;
        RECT 1513.5200 982.3800 1515.1200 982.8600 ;
        RECT 1513.5200 987.8200 1515.1200 988.3000 ;
        RECT 1513.5200 993.2600 1515.1200 993.7400 ;
        RECT 1513.5200 1036.7800 1515.1200 1037.2600 ;
        RECT 1520.6800 1036.7800 1522.2800 1037.2600 ;
        RECT 1565.6800 1036.7800 1567.2800 1037.2600 ;
        RECT 1610.6800 1036.7800 1612.2800 1037.2600 ;
        RECT 1716.2200 971.5000 1717.8200 971.9800 ;
        RECT 1716.2200 976.9400 1717.8200 977.4200 ;
        RECT 1700.6800 971.5000 1702.2800 971.9800 ;
        RECT 1700.6800 976.9400 1702.2800 977.4200 ;
        RECT 1716.2200 955.1800 1717.8200 955.6600 ;
        RECT 1716.2200 960.6200 1717.8200 961.1000 ;
        RECT 1716.2200 966.0600 1717.8200 966.5400 ;
        RECT 1700.6800 955.1800 1702.2800 955.6600 ;
        RECT 1700.6800 960.6200 1702.2800 961.1000 ;
        RECT 1700.6800 966.0600 1702.2800 966.5400 ;
        RECT 1716.2200 944.3000 1717.8200 944.7800 ;
        RECT 1716.2200 949.7400 1717.8200 950.2200 ;
        RECT 1700.6800 944.3000 1702.2800 944.7800 ;
        RECT 1700.6800 949.7400 1702.2800 950.2200 ;
        RECT 1716.2200 927.9800 1717.8200 928.4600 ;
        RECT 1716.2200 933.4200 1717.8200 933.9000 ;
        RECT 1716.2200 938.8600 1717.8200 939.3400 ;
        RECT 1700.6800 927.9800 1702.2800 928.4600 ;
        RECT 1700.6800 933.4200 1702.2800 933.9000 ;
        RECT 1700.6800 938.8600 1702.2800 939.3400 ;
        RECT 1655.6800 971.5000 1657.2800 971.9800 ;
        RECT 1655.6800 976.9400 1657.2800 977.4200 ;
        RECT 1655.6800 955.1800 1657.2800 955.6600 ;
        RECT 1655.6800 960.6200 1657.2800 961.1000 ;
        RECT 1655.6800 966.0600 1657.2800 966.5400 ;
        RECT 1655.6800 944.3000 1657.2800 944.7800 ;
        RECT 1655.6800 949.7400 1657.2800 950.2200 ;
        RECT 1655.6800 927.9800 1657.2800 928.4600 ;
        RECT 1655.6800 933.4200 1657.2800 933.9000 ;
        RECT 1655.6800 938.8600 1657.2800 939.3400 ;
        RECT 1716.2200 917.1000 1717.8200 917.5800 ;
        RECT 1716.2200 922.5400 1717.8200 923.0200 ;
        RECT 1700.6800 917.1000 1702.2800 917.5800 ;
        RECT 1700.6800 922.5400 1702.2800 923.0200 ;
        RECT 1716.2200 900.7800 1717.8200 901.2600 ;
        RECT 1716.2200 906.2200 1717.8200 906.7000 ;
        RECT 1716.2200 911.6600 1717.8200 912.1400 ;
        RECT 1700.6800 900.7800 1702.2800 901.2600 ;
        RECT 1700.6800 906.2200 1702.2800 906.7000 ;
        RECT 1700.6800 911.6600 1702.2800 912.1400 ;
        RECT 1716.2200 889.9000 1717.8200 890.3800 ;
        RECT 1716.2200 895.3400 1717.8200 895.8200 ;
        RECT 1700.6800 889.9000 1702.2800 890.3800 ;
        RECT 1700.6800 895.3400 1702.2800 895.8200 ;
        RECT 1700.6800 884.4600 1702.2800 884.9400 ;
        RECT 1716.2200 884.4600 1717.8200 884.9400 ;
        RECT 1655.6800 917.1000 1657.2800 917.5800 ;
        RECT 1655.6800 922.5400 1657.2800 923.0200 ;
        RECT 1655.6800 900.7800 1657.2800 901.2600 ;
        RECT 1655.6800 906.2200 1657.2800 906.7000 ;
        RECT 1655.6800 911.6600 1657.2800 912.1400 ;
        RECT 1655.6800 889.9000 1657.2800 890.3800 ;
        RECT 1655.6800 895.3400 1657.2800 895.8200 ;
        RECT 1655.6800 884.4600 1657.2800 884.9400 ;
        RECT 1610.6800 971.5000 1612.2800 971.9800 ;
        RECT 1610.6800 976.9400 1612.2800 977.4200 ;
        RECT 1610.6800 955.1800 1612.2800 955.6600 ;
        RECT 1610.6800 960.6200 1612.2800 961.1000 ;
        RECT 1610.6800 966.0600 1612.2800 966.5400 ;
        RECT 1565.6800 971.5000 1567.2800 971.9800 ;
        RECT 1565.6800 976.9400 1567.2800 977.4200 ;
        RECT 1565.6800 955.1800 1567.2800 955.6600 ;
        RECT 1565.6800 960.6200 1567.2800 961.1000 ;
        RECT 1565.6800 966.0600 1567.2800 966.5400 ;
        RECT 1610.6800 944.3000 1612.2800 944.7800 ;
        RECT 1610.6800 949.7400 1612.2800 950.2200 ;
        RECT 1610.6800 927.9800 1612.2800 928.4600 ;
        RECT 1610.6800 933.4200 1612.2800 933.9000 ;
        RECT 1610.6800 938.8600 1612.2800 939.3400 ;
        RECT 1565.6800 944.3000 1567.2800 944.7800 ;
        RECT 1565.6800 949.7400 1567.2800 950.2200 ;
        RECT 1565.6800 927.9800 1567.2800 928.4600 ;
        RECT 1565.6800 933.4200 1567.2800 933.9000 ;
        RECT 1565.6800 938.8600 1567.2800 939.3400 ;
        RECT 1520.6800 971.5000 1522.2800 971.9800 ;
        RECT 1520.6800 976.9400 1522.2800 977.4200 ;
        RECT 1513.5200 971.5000 1515.1200 971.9800 ;
        RECT 1513.5200 976.9400 1515.1200 977.4200 ;
        RECT 1520.6800 955.1800 1522.2800 955.6600 ;
        RECT 1520.6800 960.6200 1522.2800 961.1000 ;
        RECT 1520.6800 966.0600 1522.2800 966.5400 ;
        RECT 1513.5200 955.1800 1515.1200 955.6600 ;
        RECT 1513.5200 960.6200 1515.1200 961.1000 ;
        RECT 1513.5200 966.0600 1515.1200 966.5400 ;
        RECT 1520.6800 944.3000 1522.2800 944.7800 ;
        RECT 1520.6800 949.7400 1522.2800 950.2200 ;
        RECT 1513.5200 944.3000 1515.1200 944.7800 ;
        RECT 1513.5200 949.7400 1515.1200 950.2200 ;
        RECT 1520.6800 927.9800 1522.2800 928.4600 ;
        RECT 1520.6800 933.4200 1522.2800 933.9000 ;
        RECT 1520.6800 938.8600 1522.2800 939.3400 ;
        RECT 1513.5200 927.9800 1515.1200 928.4600 ;
        RECT 1513.5200 933.4200 1515.1200 933.9000 ;
        RECT 1513.5200 938.8600 1515.1200 939.3400 ;
        RECT 1610.6800 917.1000 1612.2800 917.5800 ;
        RECT 1610.6800 922.5400 1612.2800 923.0200 ;
        RECT 1610.6800 900.7800 1612.2800 901.2600 ;
        RECT 1610.6800 906.2200 1612.2800 906.7000 ;
        RECT 1610.6800 911.6600 1612.2800 912.1400 ;
        RECT 1565.6800 917.1000 1567.2800 917.5800 ;
        RECT 1565.6800 922.5400 1567.2800 923.0200 ;
        RECT 1565.6800 900.7800 1567.2800 901.2600 ;
        RECT 1565.6800 906.2200 1567.2800 906.7000 ;
        RECT 1565.6800 911.6600 1567.2800 912.1400 ;
        RECT 1610.6800 895.3400 1612.2800 895.8200 ;
        RECT 1610.6800 889.9000 1612.2800 890.3800 ;
        RECT 1610.6800 884.4600 1612.2800 884.9400 ;
        RECT 1565.6800 895.3400 1567.2800 895.8200 ;
        RECT 1565.6800 889.9000 1567.2800 890.3800 ;
        RECT 1565.6800 884.4600 1567.2800 884.9400 ;
        RECT 1520.6800 917.1000 1522.2800 917.5800 ;
        RECT 1520.6800 922.5400 1522.2800 923.0200 ;
        RECT 1513.5200 917.1000 1515.1200 917.5800 ;
        RECT 1513.5200 922.5400 1515.1200 923.0200 ;
        RECT 1520.6800 900.7800 1522.2800 901.2600 ;
        RECT 1520.6800 906.2200 1522.2800 906.7000 ;
        RECT 1520.6800 911.6600 1522.2800 912.1400 ;
        RECT 1513.5200 900.7800 1515.1200 901.2600 ;
        RECT 1513.5200 906.2200 1515.1200 906.7000 ;
        RECT 1513.5200 911.6600 1515.1200 912.1400 ;
        RECT 1520.6800 889.9000 1522.2800 890.3800 ;
        RECT 1520.6800 895.3400 1522.2800 895.8200 ;
        RECT 1513.5200 889.9000 1515.1200 890.3800 ;
        RECT 1513.5200 895.3400 1515.1200 895.8200 ;
        RECT 1513.5200 884.4600 1515.1200 884.9400 ;
        RECT 1520.6800 884.4600 1522.2800 884.9400 ;
        RECT 1510.5600 1086.6500 1720.7800 1088.2500 ;
        RECT 1510.5600 874.9500 1720.7800 876.5500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 872.1200 1515.1200 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 1090.1600 1515.1200 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 872.1200 1717.8200 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 1090.1600 1717.8200 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 874.9500 1512.1600 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 874.9500 1720.7800 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1086.6500 1512.1600 1088.2500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1086.6500 1720.7800 1088.2500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 645.3100 1702.2800 858.6100 ;
        RECT 1655.6800 645.3100 1657.2800 858.6100 ;
        RECT 1610.6800 645.3100 1612.2800 858.6100 ;
        RECT 1565.6800 645.3100 1567.2800 858.6100 ;
        RECT 1520.6800 645.3100 1522.2800 858.6100 ;
        RECT 1716.2200 642.4800 1717.8200 862.1200 ;
        RECT 1513.5200 642.4800 1515.1200 862.1200 ;
      LAYER met3 ;
        RECT 1700.6800 850.6600 1702.2800 851.1400 ;
        RECT 1716.2200 850.6600 1717.8200 851.1400 ;
        RECT 1716.2200 839.7800 1717.8200 840.2600 ;
        RECT 1716.2200 845.2200 1717.8200 845.7000 ;
        RECT 1700.6800 839.7800 1702.2800 840.2600 ;
        RECT 1700.6800 845.2200 1702.2800 845.7000 ;
        RECT 1716.2200 823.4600 1717.8200 823.9400 ;
        RECT 1716.2200 828.9000 1717.8200 829.3800 ;
        RECT 1700.6800 823.4600 1702.2800 823.9400 ;
        RECT 1700.6800 828.9000 1702.2800 829.3800 ;
        RECT 1716.2200 812.5800 1717.8200 813.0600 ;
        RECT 1716.2200 818.0200 1717.8200 818.5000 ;
        RECT 1700.6800 812.5800 1702.2800 813.0600 ;
        RECT 1700.6800 818.0200 1702.2800 818.5000 ;
        RECT 1700.6800 834.3400 1702.2800 834.8200 ;
        RECT 1716.2200 834.3400 1717.8200 834.8200 ;
        RECT 1655.6800 839.7800 1657.2800 840.2600 ;
        RECT 1655.6800 845.2200 1657.2800 845.7000 ;
        RECT 1655.6800 850.6600 1657.2800 851.1400 ;
        RECT 1655.6800 823.4600 1657.2800 823.9400 ;
        RECT 1655.6800 828.9000 1657.2800 829.3800 ;
        RECT 1655.6800 818.0200 1657.2800 818.5000 ;
        RECT 1655.6800 812.5800 1657.2800 813.0600 ;
        RECT 1655.6800 834.3400 1657.2800 834.8200 ;
        RECT 1716.2200 796.2600 1717.8200 796.7400 ;
        RECT 1716.2200 801.7000 1717.8200 802.1800 ;
        RECT 1700.6800 796.2600 1702.2800 796.7400 ;
        RECT 1700.6800 801.7000 1702.2800 802.1800 ;
        RECT 1716.2200 779.9400 1717.8200 780.4200 ;
        RECT 1716.2200 785.3800 1717.8200 785.8600 ;
        RECT 1716.2200 790.8200 1717.8200 791.3000 ;
        RECT 1700.6800 779.9400 1702.2800 780.4200 ;
        RECT 1700.6800 785.3800 1702.2800 785.8600 ;
        RECT 1700.6800 790.8200 1702.2800 791.3000 ;
        RECT 1716.2200 769.0600 1717.8200 769.5400 ;
        RECT 1716.2200 774.5000 1717.8200 774.9800 ;
        RECT 1700.6800 769.0600 1702.2800 769.5400 ;
        RECT 1700.6800 774.5000 1702.2800 774.9800 ;
        RECT 1716.2200 752.7400 1717.8200 753.2200 ;
        RECT 1716.2200 758.1800 1717.8200 758.6600 ;
        RECT 1716.2200 763.6200 1717.8200 764.1000 ;
        RECT 1700.6800 752.7400 1702.2800 753.2200 ;
        RECT 1700.6800 758.1800 1702.2800 758.6600 ;
        RECT 1700.6800 763.6200 1702.2800 764.1000 ;
        RECT 1655.6800 796.2600 1657.2800 796.7400 ;
        RECT 1655.6800 801.7000 1657.2800 802.1800 ;
        RECT 1655.6800 779.9400 1657.2800 780.4200 ;
        RECT 1655.6800 785.3800 1657.2800 785.8600 ;
        RECT 1655.6800 790.8200 1657.2800 791.3000 ;
        RECT 1655.6800 769.0600 1657.2800 769.5400 ;
        RECT 1655.6800 774.5000 1657.2800 774.9800 ;
        RECT 1655.6800 752.7400 1657.2800 753.2200 ;
        RECT 1655.6800 758.1800 1657.2800 758.6600 ;
        RECT 1655.6800 763.6200 1657.2800 764.1000 ;
        RECT 1655.6800 807.1400 1657.2800 807.6200 ;
        RECT 1700.6800 807.1400 1702.2800 807.6200 ;
        RECT 1716.2200 807.1400 1717.8200 807.6200 ;
        RECT 1610.6800 839.7800 1612.2800 840.2600 ;
        RECT 1610.6800 845.2200 1612.2800 845.7000 ;
        RECT 1610.6800 850.6600 1612.2800 851.1400 ;
        RECT 1565.6800 839.7800 1567.2800 840.2600 ;
        RECT 1565.6800 845.2200 1567.2800 845.7000 ;
        RECT 1565.6800 850.6600 1567.2800 851.1400 ;
        RECT 1610.6800 823.4600 1612.2800 823.9400 ;
        RECT 1610.6800 828.9000 1612.2800 829.3800 ;
        RECT 1610.6800 812.5800 1612.2800 813.0600 ;
        RECT 1610.6800 818.0200 1612.2800 818.5000 ;
        RECT 1565.6800 823.4600 1567.2800 823.9400 ;
        RECT 1565.6800 828.9000 1567.2800 829.3800 ;
        RECT 1565.6800 812.5800 1567.2800 813.0600 ;
        RECT 1565.6800 818.0200 1567.2800 818.5000 ;
        RECT 1565.6800 834.3400 1567.2800 834.8200 ;
        RECT 1610.6800 834.3400 1612.2800 834.8200 ;
        RECT 1513.5200 850.6600 1515.1200 851.1400 ;
        RECT 1520.6800 850.6600 1522.2800 851.1400 ;
        RECT 1520.6800 839.7800 1522.2800 840.2600 ;
        RECT 1520.6800 845.2200 1522.2800 845.7000 ;
        RECT 1513.5200 839.7800 1515.1200 840.2600 ;
        RECT 1513.5200 845.2200 1515.1200 845.7000 ;
        RECT 1520.6800 823.4600 1522.2800 823.9400 ;
        RECT 1520.6800 828.9000 1522.2800 829.3800 ;
        RECT 1513.5200 823.4600 1515.1200 823.9400 ;
        RECT 1513.5200 828.9000 1515.1200 829.3800 ;
        RECT 1520.6800 812.5800 1522.2800 813.0600 ;
        RECT 1520.6800 818.0200 1522.2800 818.5000 ;
        RECT 1513.5200 812.5800 1515.1200 813.0600 ;
        RECT 1513.5200 818.0200 1515.1200 818.5000 ;
        RECT 1513.5200 834.3400 1515.1200 834.8200 ;
        RECT 1520.6800 834.3400 1522.2800 834.8200 ;
        RECT 1610.6800 796.2600 1612.2800 796.7400 ;
        RECT 1610.6800 801.7000 1612.2800 802.1800 ;
        RECT 1610.6800 779.9400 1612.2800 780.4200 ;
        RECT 1610.6800 785.3800 1612.2800 785.8600 ;
        RECT 1610.6800 790.8200 1612.2800 791.3000 ;
        RECT 1565.6800 796.2600 1567.2800 796.7400 ;
        RECT 1565.6800 801.7000 1567.2800 802.1800 ;
        RECT 1565.6800 779.9400 1567.2800 780.4200 ;
        RECT 1565.6800 785.3800 1567.2800 785.8600 ;
        RECT 1565.6800 790.8200 1567.2800 791.3000 ;
        RECT 1610.6800 769.0600 1612.2800 769.5400 ;
        RECT 1610.6800 774.5000 1612.2800 774.9800 ;
        RECT 1610.6800 752.7400 1612.2800 753.2200 ;
        RECT 1610.6800 758.1800 1612.2800 758.6600 ;
        RECT 1610.6800 763.6200 1612.2800 764.1000 ;
        RECT 1565.6800 769.0600 1567.2800 769.5400 ;
        RECT 1565.6800 774.5000 1567.2800 774.9800 ;
        RECT 1565.6800 752.7400 1567.2800 753.2200 ;
        RECT 1565.6800 758.1800 1567.2800 758.6600 ;
        RECT 1565.6800 763.6200 1567.2800 764.1000 ;
        RECT 1520.6800 796.2600 1522.2800 796.7400 ;
        RECT 1520.6800 801.7000 1522.2800 802.1800 ;
        RECT 1513.5200 796.2600 1515.1200 796.7400 ;
        RECT 1513.5200 801.7000 1515.1200 802.1800 ;
        RECT 1520.6800 779.9400 1522.2800 780.4200 ;
        RECT 1520.6800 785.3800 1522.2800 785.8600 ;
        RECT 1520.6800 790.8200 1522.2800 791.3000 ;
        RECT 1513.5200 779.9400 1515.1200 780.4200 ;
        RECT 1513.5200 785.3800 1515.1200 785.8600 ;
        RECT 1513.5200 790.8200 1515.1200 791.3000 ;
        RECT 1520.6800 769.0600 1522.2800 769.5400 ;
        RECT 1520.6800 774.5000 1522.2800 774.9800 ;
        RECT 1513.5200 769.0600 1515.1200 769.5400 ;
        RECT 1513.5200 774.5000 1515.1200 774.9800 ;
        RECT 1520.6800 752.7400 1522.2800 753.2200 ;
        RECT 1520.6800 758.1800 1522.2800 758.6600 ;
        RECT 1520.6800 763.6200 1522.2800 764.1000 ;
        RECT 1513.5200 752.7400 1515.1200 753.2200 ;
        RECT 1513.5200 758.1800 1515.1200 758.6600 ;
        RECT 1513.5200 763.6200 1515.1200 764.1000 ;
        RECT 1513.5200 807.1400 1515.1200 807.6200 ;
        RECT 1520.6800 807.1400 1522.2800 807.6200 ;
        RECT 1565.6800 807.1400 1567.2800 807.6200 ;
        RECT 1610.6800 807.1400 1612.2800 807.6200 ;
        RECT 1716.2200 741.8600 1717.8200 742.3400 ;
        RECT 1716.2200 747.3000 1717.8200 747.7800 ;
        RECT 1700.6800 741.8600 1702.2800 742.3400 ;
        RECT 1700.6800 747.3000 1702.2800 747.7800 ;
        RECT 1716.2200 725.5400 1717.8200 726.0200 ;
        RECT 1716.2200 730.9800 1717.8200 731.4600 ;
        RECT 1716.2200 736.4200 1717.8200 736.9000 ;
        RECT 1700.6800 725.5400 1702.2800 726.0200 ;
        RECT 1700.6800 730.9800 1702.2800 731.4600 ;
        RECT 1700.6800 736.4200 1702.2800 736.9000 ;
        RECT 1716.2200 714.6600 1717.8200 715.1400 ;
        RECT 1716.2200 720.1000 1717.8200 720.5800 ;
        RECT 1700.6800 714.6600 1702.2800 715.1400 ;
        RECT 1700.6800 720.1000 1702.2800 720.5800 ;
        RECT 1716.2200 698.3400 1717.8200 698.8200 ;
        RECT 1716.2200 703.7800 1717.8200 704.2600 ;
        RECT 1716.2200 709.2200 1717.8200 709.7000 ;
        RECT 1700.6800 698.3400 1702.2800 698.8200 ;
        RECT 1700.6800 703.7800 1702.2800 704.2600 ;
        RECT 1700.6800 709.2200 1702.2800 709.7000 ;
        RECT 1655.6800 741.8600 1657.2800 742.3400 ;
        RECT 1655.6800 747.3000 1657.2800 747.7800 ;
        RECT 1655.6800 725.5400 1657.2800 726.0200 ;
        RECT 1655.6800 730.9800 1657.2800 731.4600 ;
        RECT 1655.6800 736.4200 1657.2800 736.9000 ;
        RECT 1655.6800 714.6600 1657.2800 715.1400 ;
        RECT 1655.6800 720.1000 1657.2800 720.5800 ;
        RECT 1655.6800 698.3400 1657.2800 698.8200 ;
        RECT 1655.6800 703.7800 1657.2800 704.2600 ;
        RECT 1655.6800 709.2200 1657.2800 709.7000 ;
        RECT 1716.2200 687.4600 1717.8200 687.9400 ;
        RECT 1716.2200 692.9000 1717.8200 693.3800 ;
        RECT 1700.6800 687.4600 1702.2800 687.9400 ;
        RECT 1700.6800 692.9000 1702.2800 693.3800 ;
        RECT 1716.2200 671.1400 1717.8200 671.6200 ;
        RECT 1716.2200 676.5800 1717.8200 677.0600 ;
        RECT 1716.2200 682.0200 1717.8200 682.5000 ;
        RECT 1700.6800 671.1400 1702.2800 671.6200 ;
        RECT 1700.6800 676.5800 1702.2800 677.0600 ;
        RECT 1700.6800 682.0200 1702.2800 682.5000 ;
        RECT 1716.2200 660.2600 1717.8200 660.7400 ;
        RECT 1716.2200 665.7000 1717.8200 666.1800 ;
        RECT 1700.6800 660.2600 1702.2800 660.7400 ;
        RECT 1700.6800 665.7000 1702.2800 666.1800 ;
        RECT 1700.6800 654.8200 1702.2800 655.3000 ;
        RECT 1716.2200 654.8200 1717.8200 655.3000 ;
        RECT 1655.6800 687.4600 1657.2800 687.9400 ;
        RECT 1655.6800 692.9000 1657.2800 693.3800 ;
        RECT 1655.6800 671.1400 1657.2800 671.6200 ;
        RECT 1655.6800 676.5800 1657.2800 677.0600 ;
        RECT 1655.6800 682.0200 1657.2800 682.5000 ;
        RECT 1655.6800 660.2600 1657.2800 660.7400 ;
        RECT 1655.6800 665.7000 1657.2800 666.1800 ;
        RECT 1655.6800 654.8200 1657.2800 655.3000 ;
        RECT 1610.6800 741.8600 1612.2800 742.3400 ;
        RECT 1610.6800 747.3000 1612.2800 747.7800 ;
        RECT 1610.6800 725.5400 1612.2800 726.0200 ;
        RECT 1610.6800 730.9800 1612.2800 731.4600 ;
        RECT 1610.6800 736.4200 1612.2800 736.9000 ;
        RECT 1565.6800 741.8600 1567.2800 742.3400 ;
        RECT 1565.6800 747.3000 1567.2800 747.7800 ;
        RECT 1565.6800 725.5400 1567.2800 726.0200 ;
        RECT 1565.6800 730.9800 1567.2800 731.4600 ;
        RECT 1565.6800 736.4200 1567.2800 736.9000 ;
        RECT 1610.6800 714.6600 1612.2800 715.1400 ;
        RECT 1610.6800 720.1000 1612.2800 720.5800 ;
        RECT 1610.6800 698.3400 1612.2800 698.8200 ;
        RECT 1610.6800 703.7800 1612.2800 704.2600 ;
        RECT 1610.6800 709.2200 1612.2800 709.7000 ;
        RECT 1565.6800 714.6600 1567.2800 715.1400 ;
        RECT 1565.6800 720.1000 1567.2800 720.5800 ;
        RECT 1565.6800 698.3400 1567.2800 698.8200 ;
        RECT 1565.6800 703.7800 1567.2800 704.2600 ;
        RECT 1565.6800 709.2200 1567.2800 709.7000 ;
        RECT 1520.6800 741.8600 1522.2800 742.3400 ;
        RECT 1520.6800 747.3000 1522.2800 747.7800 ;
        RECT 1513.5200 741.8600 1515.1200 742.3400 ;
        RECT 1513.5200 747.3000 1515.1200 747.7800 ;
        RECT 1520.6800 725.5400 1522.2800 726.0200 ;
        RECT 1520.6800 730.9800 1522.2800 731.4600 ;
        RECT 1520.6800 736.4200 1522.2800 736.9000 ;
        RECT 1513.5200 725.5400 1515.1200 726.0200 ;
        RECT 1513.5200 730.9800 1515.1200 731.4600 ;
        RECT 1513.5200 736.4200 1515.1200 736.9000 ;
        RECT 1520.6800 714.6600 1522.2800 715.1400 ;
        RECT 1520.6800 720.1000 1522.2800 720.5800 ;
        RECT 1513.5200 714.6600 1515.1200 715.1400 ;
        RECT 1513.5200 720.1000 1515.1200 720.5800 ;
        RECT 1520.6800 698.3400 1522.2800 698.8200 ;
        RECT 1520.6800 703.7800 1522.2800 704.2600 ;
        RECT 1520.6800 709.2200 1522.2800 709.7000 ;
        RECT 1513.5200 698.3400 1515.1200 698.8200 ;
        RECT 1513.5200 703.7800 1515.1200 704.2600 ;
        RECT 1513.5200 709.2200 1515.1200 709.7000 ;
        RECT 1610.6800 687.4600 1612.2800 687.9400 ;
        RECT 1610.6800 692.9000 1612.2800 693.3800 ;
        RECT 1610.6800 671.1400 1612.2800 671.6200 ;
        RECT 1610.6800 676.5800 1612.2800 677.0600 ;
        RECT 1610.6800 682.0200 1612.2800 682.5000 ;
        RECT 1565.6800 687.4600 1567.2800 687.9400 ;
        RECT 1565.6800 692.9000 1567.2800 693.3800 ;
        RECT 1565.6800 671.1400 1567.2800 671.6200 ;
        RECT 1565.6800 676.5800 1567.2800 677.0600 ;
        RECT 1565.6800 682.0200 1567.2800 682.5000 ;
        RECT 1610.6800 665.7000 1612.2800 666.1800 ;
        RECT 1610.6800 660.2600 1612.2800 660.7400 ;
        RECT 1610.6800 654.8200 1612.2800 655.3000 ;
        RECT 1565.6800 665.7000 1567.2800 666.1800 ;
        RECT 1565.6800 660.2600 1567.2800 660.7400 ;
        RECT 1565.6800 654.8200 1567.2800 655.3000 ;
        RECT 1520.6800 687.4600 1522.2800 687.9400 ;
        RECT 1520.6800 692.9000 1522.2800 693.3800 ;
        RECT 1513.5200 687.4600 1515.1200 687.9400 ;
        RECT 1513.5200 692.9000 1515.1200 693.3800 ;
        RECT 1520.6800 671.1400 1522.2800 671.6200 ;
        RECT 1520.6800 676.5800 1522.2800 677.0600 ;
        RECT 1520.6800 682.0200 1522.2800 682.5000 ;
        RECT 1513.5200 671.1400 1515.1200 671.6200 ;
        RECT 1513.5200 676.5800 1515.1200 677.0600 ;
        RECT 1513.5200 682.0200 1515.1200 682.5000 ;
        RECT 1520.6800 660.2600 1522.2800 660.7400 ;
        RECT 1520.6800 665.7000 1522.2800 666.1800 ;
        RECT 1513.5200 660.2600 1515.1200 660.7400 ;
        RECT 1513.5200 665.7000 1515.1200 666.1800 ;
        RECT 1513.5200 654.8200 1515.1200 655.3000 ;
        RECT 1520.6800 654.8200 1522.2800 655.3000 ;
        RECT 1510.5600 857.0100 1720.7800 858.6100 ;
        RECT 1510.5600 645.3100 1720.7800 646.9100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 642.4800 1515.1200 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 860.5200 1515.1200 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 642.4800 1717.8200 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 860.5200 1717.8200 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 645.3100 1512.1600 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 645.3100 1720.7800 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 857.0100 1512.1600 858.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 857.0100 1720.7800 858.6100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1700.6800 415.6700 1702.2800 628.9700 ;
        RECT 1655.6800 415.6700 1657.2800 628.9700 ;
        RECT 1610.6800 415.6700 1612.2800 628.9700 ;
        RECT 1565.6800 415.6700 1567.2800 628.9700 ;
        RECT 1520.6800 415.6700 1522.2800 628.9700 ;
        RECT 1716.2200 412.8400 1717.8200 632.4800 ;
        RECT 1513.5200 412.8400 1515.1200 632.4800 ;
      LAYER met3 ;
        RECT 1700.6800 621.0200 1702.2800 621.5000 ;
        RECT 1716.2200 621.0200 1717.8200 621.5000 ;
        RECT 1716.2200 610.1400 1717.8200 610.6200 ;
        RECT 1716.2200 615.5800 1717.8200 616.0600 ;
        RECT 1700.6800 610.1400 1702.2800 610.6200 ;
        RECT 1700.6800 615.5800 1702.2800 616.0600 ;
        RECT 1716.2200 593.8200 1717.8200 594.3000 ;
        RECT 1716.2200 599.2600 1717.8200 599.7400 ;
        RECT 1700.6800 593.8200 1702.2800 594.3000 ;
        RECT 1700.6800 599.2600 1702.2800 599.7400 ;
        RECT 1716.2200 582.9400 1717.8200 583.4200 ;
        RECT 1716.2200 588.3800 1717.8200 588.8600 ;
        RECT 1700.6800 582.9400 1702.2800 583.4200 ;
        RECT 1700.6800 588.3800 1702.2800 588.8600 ;
        RECT 1700.6800 604.7000 1702.2800 605.1800 ;
        RECT 1716.2200 604.7000 1717.8200 605.1800 ;
        RECT 1655.6800 610.1400 1657.2800 610.6200 ;
        RECT 1655.6800 615.5800 1657.2800 616.0600 ;
        RECT 1655.6800 621.0200 1657.2800 621.5000 ;
        RECT 1655.6800 593.8200 1657.2800 594.3000 ;
        RECT 1655.6800 599.2600 1657.2800 599.7400 ;
        RECT 1655.6800 588.3800 1657.2800 588.8600 ;
        RECT 1655.6800 582.9400 1657.2800 583.4200 ;
        RECT 1655.6800 604.7000 1657.2800 605.1800 ;
        RECT 1716.2200 566.6200 1717.8200 567.1000 ;
        RECT 1716.2200 572.0600 1717.8200 572.5400 ;
        RECT 1700.6800 566.6200 1702.2800 567.1000 ;
        RECT 1700.6800 572.0600 1702.2800 572.5400 ;
        RECT 1716.2200 550.3000 1717.8200 550.7800 ;
        RECT 1716.2200 555.7400 1717.8200 556.2200 ;
        RECT 1716.2200 561.1800 1717.8200 561.6600 ;
        RECT 1700.6800 550.3000 1702.2800 550.7800 ;
        RECT 1700.6800 555.7400 1702.2800 556.2200 ;
        RECT 1700.6800 561.1800 1702.2800 561.6600 ;
        RECT 1716.2200 539.4200 1717.8200 539.9000 ;
        RECT 1716.2200 544.8600 1717.8200 545.3400 ;
        RECT 1700.6800 539.4200 1702.2800 539.9000 ;
        RECT 1700.6800 544.8600 1702.2800 545.3400 ;
        RECT 1716.2200 523.1000 1717.8200 523.5800 ;
        RECT 1716.2200 528.5400 1717.8200 529.0200 ;
        RECT 1716.2200 533.9800 1717.8200 534.4600 ;
        RECT 1700.6800 523.1000 1702.2800 523.5800 ;
        RECT 1700.6800 528.5400 1702.2800 529.0200 ;
        RECT 1700.6800 533.9800 1702.2800 534.4600 ;
        RECT 1655.6800 566.6200 1657.2800 567.1000 ;
        RECT 1655.6800 572.0600 1657.2800 572.5400 ;
        RECT 1655.6800 550.3000 1657.2800 550.7800 ;
        RECT 1655.6800 555.7400 1657.2800 556.2200 ;
        RECT 1655.6800 561.1800 1657.2800 561.6600 ;
        RECT 1655.6800 539.4200 1657.2800 539.9000 ;
        RECT 1655.6800 544.8600 1657.2800 545.3400 ;
        RECT 1655.6800 523.1000 1657.2800 523.5800 ;
        RECT 1655.6800 528.5400 1657.2800 529.0200 ;
        RECT 1655.6800 533.9800 1657.2800 534.4600 ;
        RECT 1655.6800 577.5000 1657.2800 577.9800 ;
        RECT 1700.6800 577.5000 1702.2800 577.9800 ;
        RECT 1716.2200 577.5000 1717.8200 577.9800 ;
        RECT 1610.6800 610.1400 1612.2800 610.6200 ;
        RECT 1610.6800 615.5800 1612.2800 616.0600 ;
        RECT 1610.6800 621.0200 1612.2800 621.5000 ;
        RECT 1565.6800 610.1400 1567.2800 610.6200 ;
        RECT 1565.6800 615.5800 1567.2800 616.0600 ;
        RECT 1565.6800 621.0200 1567.2800 621.5000 ;
        RECT 1610.6800 593.8200 1612.2800 594.3000 ;
        RECT 1610.6800 599.2600 1612.2800 599.7400 ;
        RECT 1610.6800 582.9400 1612.2800 583.4200 ;
        RECT 1610.6800 588.3800 1612.2800 588.8600 ;
        RECT 1565.6800 593.8200 1567.2800 594.3000 ;
        RECT 1565.6800 599.2600 1567.2800 599.7400 ;
        RECT 1565.6800 582.9400 1567.2800 583.4200 ;
        RECT 1565.6800 588.3800 1567.2800 588.8600 ;
        RECT 1565.6800 604.7000 1567.2800 605.1800 ;
        RECT 1610.6800 604.7000 1612.2800 605.1800 ;
        RECT 1513.5200 621.0200 1515.1200 621.5000 ;
        RECT 1520.6800 621.0200 1522.2800 621.5000 ;
        RECT 1520.6800 610.1400 1522.2800 610.6200 ;
        RECT 1520.6800 615.5800 1522.2800 616.0600 ;
        RECT 1513.5200 610.1400 1515.1200 610.6200 ;
        RECT 1513.5200 615.5800 1515.1200 616.0600 ;
        RECT 1520.6800 593.8200 1522.2800 594.3000 ;
        RECT 1520.6800 599.2600 1522.2800 599.7400 ;
        RECT 1513.5200 593.8200 1515.1200 594.3000 ;
        RECT 1513.5200 599.2600 1515.1200 599.7400 ;
        RECT 1520.6800 582.9400 1522.2800 583.4200 ;
        RECT 1520.6800 588.3800 1522.2800 588.8600 ;
        RECT 1513.5200 582.9400 1515.1200 583.4200 ;
        RECT 1513.5200 588.3800 1515.1200 588.8600 ;
        RECT 1513.5200 604.7000 1515.1200 605.1800 ;
        RECT 1520.6800 604.7000 1522.2800 605.1800 ;
        RECT 1610.6800 566.6200 1612.2800 567.1000 ;
        RECT 1610.6800 572.0600 1612.2800 572.5400 ;
        RECT 1610.6800 550.3000 1612.2800 550.7800 ;
        RECT 1610.6800 555.7400 1612.2800 556.2200 ;
        RECT 1610.6800 561.1800 1612.2800 561.6600 ;
        RECT 1565.6800 566.6200 1567.2800 567.1000 ;
        RECT 1565.6800 572.0600 1567.2800 572.5400 ;
        RECT 1565.6800 550.3000 1567.2800 550.7800 ;
        RECT 1565.6800 555.7400 1567.2800 556.2200 ;
        RECT 1565.6800 561.1800 1567.2800 561.6600 ;
        RECT 1610.6800 539.4200 1612.2800 539.9000 ;
        RECT 1610.6800 544.8600 1612.2800 545.3400 ;
        RECT 1610.6800 523.1000 1612.2800 523.5800 ;
        RECT 1610.6800 528.5400 1612.2800 529.0200 ;
        RECT 1610.6800 533.9800 1612.2800 534.4600 ;
        RECT 1565.6800 539.4200 1567.2800 539.9000 ;
        RECT 1565.6800 544.8600 1567.2800 545.3400 ;
        RECT 1565.6800 523.1000 1567.2800 523.5800 ;
        RECT 1565.6800 528.5400 1567.2800 529.0200 ;
        RECT 1565.6800 533.9800 1567.2800 534.4600 ;
        RECT 1520.6800 566.6200 1522.2800 567.1000 ;
        RECT 1520.6800 572.0600 1522.2800 572.5400 ;
        RECT 1513.5200 566.6200 1515.1200 567.1000 ;
        RECT 1513.5200 572.0600 1515.1200 572.5400 ;
        RECT 1520.6800 550.3000 1522.2800 550.7800 ;
        RECT 1520.6800 555.7400 1522.2800 556.2200 ;
        RECT 1520.6800 561.1800 1522.2800 561.6600 ;
        RECT 1513.5200 550.3000 1515.1200 550.7800 ;
        RECT 1513.5200 555.7400 1515.1200 556.2200 ;
        RECT 1513.5200 561.1800 1515.1200 561.6600 ;
        RECT 1520.6800 539.4200 1522.2800 539.9000 ;
        RECT 1520.6800 544.8600 1522.2800 545.3400 ;
        RECT 1513.5200 539.4200 1515.1200 539.9000 ;
        RECT 1513.5200 544.8600 1515.1200 545.3400 ;
        RECT 1520.6800 523.1000 1522.2800 523.5800 ;
        RECT 1520.6800 528.5400 1522.2800 529.0200 ;
        RECT 1520.6800 533.9800 1522.2800 534.4600 ;
        RECT 1513.5200 523.1000 1515.1200 523.5800 ;
        RECT 1513.5200 528.5400 1515.1200 529.0200 ;
        RECT 1513.5200 533.9800 1515.1200 534.4600 ;
        RECT 1513.5200 577.5000 1515.1200 577.9800 ;
        RECT 1520.6800 577.5000 1522.2800 577.9800 ;
        RECT 1565.6800 577.5000 1567.2800 577.9800 ;
        RECT 1610.6800 577.5000 1612.2800 577.9800 ;
        RECT 1716.2200 512.2200 1717.8200 512.7000 ;
        RECT 1716.2200 517.6600 1717.8200 518.1400 ;
        RECT 1700.6800 512.2200 1702.2800 512.7000 ;
        RECT 1700.6800 517.6600 1702.2800 518.1400 ;
        RECT 1716.2200 495.9000 1717.8200 496.3800 ;
        RECT 1716.2200 501.3400 1717.8200 501.8200 ;
        RECT 1716.2200 506.7800 1717.8200 507.2600 ;
        RECT 1700.6800 495.9000 1702.2800 496.3800 ;
        RECT 1700.6800 501.3400 1702.2800 501.8200 ;
        RECT 1700.6800 506.7800 1702.2800 507.2600 ;
        RECT 1716.2200 485.0200 1717.8200 485.5000 ;
        RECT 1716.2200 490.4600 1717.8200 490.9400 ;
        RECT 1700.6800 485.0200 1702.2800 485.5000 ;
        RECT 1700.6800 490.4600 1702.2800 490.9400 ;
        RECT 1716.2200 468.7000 1717.8200 469.1800 ;
        RECT 1716.2200 474.1400 1717.8200 474.6200 ;
        RECT 1716.2200 479.5800 1717.8200 480.0600 ;
        RECT 1700.6800 468.7000 1702.2800 469.1800 ;
        RECT 1700.6800 474.1400 1702.2800 474.6200 ;
        RECT 1700.6800 479.5800 1702.2800 480.0600 ;
        RECT 1655.6800 512.2200 1657.2800 512.7000 ;
        RECT 1655.6800 517.6600 1657.2800 518.1400 ;
        RECT 1655.6800 495.9000 1657.2800 496.3800 ;
        RECT 1655.6800 501.3400 1657.2800 501.8200 ;
        RECT 1655.6800 506.7800 1657.2800 507.2600 ;
        RECT 1655.6800 485.0200 1657.2800 485.5000 ;
        RECT 1655.6800 490.4600 1657.2800 490.9400 ;
        RECT 1655.6800 468.7000 1657.2800 469.1800 ;
        RECT 1655.6800 474.1400 1657.2800 474.6200 ;
        RECT 1655.6800 479.5800 1657.2800 480.0600 ;
        RECT 1716.2200 457.8200 1717.8200 458.3000 ;
        RECT 1716.2200 463.2600 1717.8200 463.7400 ;
        RECT 1700.6800 457.8200 1702.2800 458.3000 ;
        RECT 1700.6800 463.2600 1702.2800 463.7400 ;
        RECT 1716.2200 441.5000 1717.8200 441.9800 ;
        RECT 1716.2200 446.9400 1717.8200 447.4200 ;
        RECT 1716.2200 452.3800 1717.8200 452.8600 ;
        RECT 1700.6800 441.5000 1702.2800 441.9800 ;
        RECT 1700.6800 446.9400 1702.2800 447.4200 ;
        RECT 1700.6800 452.3800 1702.2800 452.8600 ;
        RECT 1716.2200 430.6200 1717.8200 431.1000 ;
        RECT 1716.2200 436.0600 1717.8200 436.5400 ;
        RECT 1700.6800 430.6200 1702.2800 431.1000 ;
        RECT 1700.6800 436.0600 1702.2800 436.5400 ;
        RECT 1700.6800 425.1800 1702.2800 425.6600 ;
        RECT 1716.2200 425.1800 1717.8200 425.6600 ;
        RECT 1655.6800 457.8200 1657.2800 458.3000 ;
        RECT 1655.6800 463.2600 1657.2800 463.7400 ;
        RECT 1655.6800 441.5000 1657.2800 441.9800 ;
        RECT 1655.6800 446.9400 1657.2800 447.4200 ;
        RECT 1655.6800 452.3800 1657.2800 452.8600 ;
        RECT 1655.6800 430.6200 1657.2800 431.1000 ;
        RECT 1655.6800 436.0600 1657.2800 436.5400 ;
        RECT 1655.6800 425.1800 1657.2800 425.6600 ;
        RECT 1610.6800 512.2200 1612.2800 512.7000 ;
        RECT 1610.6800 517.6600 1612.2800 518.1400 ;
        RECT 1610.6800 495.9000 1612.2800 496.3800 ;
        RECT 1610.6800 501.3400 1612.2800 501.8200 ;
        RECT 1610.6800 506.7800 1612.2800 507.2600 ;
        RECT 1565.6800 512.2200 1567.2800 512.7000 ;
        RECT 1565.6800 517.6600 1567.2800 518.1400 ;
        RECT 1565.6800 495.9000 1567.2800 496.3800 ;
        RECT 1565.6800 501.3400 1567.2800 501.8200 ;
        RECT 1565.6800 506.7800 1567.2800 507.2600 ;
        RECT 1610.6800 485.0200 1612.2800 485.5000 ;
        RECT 1610.6800 490.4600 1612.2800 490.9400 ;
        RECT 1610.6800 468.7000 1612.2800 469.1800 ;
        RECT 1610.6800 474.1400 1612.2800 474.6200 ;
        RECT 1610.6800 479.5800 1612.2800 480.0600 ;
        RECT 1565.6800 485.0200 1567.2800 485.5000 ;
        RECT 1565.6800 490.4600 1567.2800 490.9400 ;
        RECT 1565.6800 468.7000 1567.2800 469.1800 ;
        RECT 1565.6800 474.1400 1567.2800 474.6200 ;
        RECT 1565.6800 479.5800 1567.2800 480.0600 ;
        RECT 1520.6800 512.2200 1522.2800 512.7000 ;
        RECT 1520.6800 517.6600 1522.2800 518.1400 ;
        RECT 1513.5200 512.2200 1515.1200 512.7000 ;
        RECT 1513.5200 517.6600 1515.1200 518.1400 ;
        RECT 1520.6800 495.9000 1522.2800 496.3800 ;
        RECT 1520.6800 501.3400 1522.2800 501.8200 ;
        RECT 1520.6800 506.7800 1522.2800 507.2600 ;
        RECT 1513.5200 495.9000 1515.1200 496.3800 ;
        RECT 1513.5200 501.3400 1515.1200 501.8200 ;
        RECT 1513.5200 506.7800 1515.1200 507.2600 ;
        RECT 1520.6800 485.0200 1522.2800 485.5000 ;
        RECT 1520.6800 490.4600 1522.2800 490.9400 ;
        RECT 1513.5200 485.0200 1515.1200 485.5000 ;
        RECT 1513.5200 490.4600 1515.1200 490.9400 ;
        RECT 1520.6800 468.7000 1522.2800 469.1800 ;
        RECT 1520.6800 474.1400 1522.2800 474.6200 ;
        RECT 1520.6800 479.5800 1522.2800 480.0600 ;
        RECT 1513.5200 468.7000 1515.1200 469.1800 ;
        RECT 1513.5200 474.1400 1515.1200 474.6200 ;
        RECT 1513.5200 479.5800 1515.1200 480.0600 ;
        RECT 1610.6800 457.8200 1612.2800 458.3000 ;
        RECT 1610.6800 463.2600 1612.2800 463.7400 ;
        RECT 1610.6800 441.5000 1612.2800 441.9800 ;
        RECT 1610.6800 446.9400 1612.2800 447.4200 ;
        RECT 1610.6800 452.3800 1612.2800 452.8600 ;
        RECT 1565.6800 457.8200 1567.2800 458.3000 ;
        RECT 1565.6800 463.2600 1567.2800 463.7400 ;
        RECT 1565.6800 441.5000 1567.2800 441.9800 ;
        RECT 1565.6800 446.9400 1567.2800 447.4200 ;
        RECT 1565.6800 452.3800 1567.2800 452.8600 ;
        RECT 1610.6800 436.0600 1612.2800 436.5400 ;
        RECT 1610.6800 430.6200 1612.2800 431.1000 ;
        RECT 1610.6800 425.1800 1612.2800 425.6600 ;
        RECT 1565.6800 436.0600 1567.2800 436.5400 ;
        RECT 1565.6800 430.6200 1567.2800 431.1000 ;
        RECT 1565.6800 425.1800 1567.2800 425.6600 ;
        RECT 1520.6800 457.8200 1522.2800 458.3000 ;
        RECT 1520.6800 463.2600 1522.2800 463.7400 ;
        RECT 1513.5200 457.8200 1515.1200 458.3000 ;
        RECT 1513.5200 463.2600 1515.1200 463.7400 ;
        RECT 1520.6800 441.5000 1522.2800 441.9800 ;
        RECT 1520.6800 446.9400 1522.2800 447.4200 ;
        RECT 1520.6800 452.3800 1522.2800 452.8600 ;
        RECT 1513.5200 441.5000 1515.1200 441.9800 ;
        RECT 1513.5200 446.9400 1515.1200 447.4200 ;
        RECT 1513.5200 452.3800 1515.1200 452.8600 ;
        RECT 1520.6800 430.6200 1522.2800 431.1000 ;
        RECT 1520.6800 436.0600 1522.2800 436.5400 ;
        RECT 1513.5200 430.6200 1515.1200 431.1000 ;
        RECT 1513.5200 436.0600 1515.1200 436.5400 ;
        RECT 1513.5200 425.1800 1515.1200 425.6600 ;
        RECT 1520.6800 425.1800 1522.2800 425.6600 ;
        RECT 1510.5600 627.3700 1720.7800 628.9700 ;
        RECT 1510.5600 415.6700 1720.7800 417.2700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 412.8400 1515.1200 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1513.5200 630.8800 1515.1200 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 412.8400 1717.8200 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1716.2200 630.8800 1717.8200 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 415.6700 1512.1600 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 415.6700 1720.7800 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 627.3700 1512.1600 628.9700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 627.3700 1720.7800 628.9700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1733.8400 2479.6000 1735.4400 2509.8600 ;
        RECT 1936.3400 2479.6000 1937.9400 2509.8600 ;
      LAYER met3 ;
        RECT 1936.3400 2500.1000 1937.9400 2500.5800 ;
        RECT 1733.8400 2500.1000 1735.4400 2500.5800 ;
        RECT 1936.3400 2489.2200 1937.9400 2489.7000 ;
        RECT 1733.8400 2489.2200 1735.4400 2489.7000 ;
        RECT 1936.3400 2494.6600 1937.9400 2495.1400 ;
        RECT 1733.8400 2494.6600 1735.4400 2495.1400 ;
        RECT 1730.7800 2505.5000 1941.0000 2507.1000 ;
        RECT 1730.7800 2481.1700 1941.0000 2482.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.8400 2479.6000 1735.4400 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.8400 2508.2600 1735.4400 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.3400 2479.6000 1937.9400 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.3400 2508.2600 1937.9400 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2481.1700 1732.3800 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2481.1700 1941.0000 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2505.5000 1732.3800 2507.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2505.5000 1941.0000 2507.1000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 186.0300 1922.5000 399.3300 ;
        RECT 1875.9000 186.0300 1877.5000 399.3300 ;
        RECT 1830.9000 186.0300 1832.5000 399.3300 ;
        RECT 1785.9000 186.0300 1787.5000 399.3300 ;
        RECT 1740.9000 186.0300 1742.5000 399.3300 ;
        RECT 1936.4400 183.2000 1938.0400 402.8400 ;
        RECT 1733.7400 183.2000 1735.3400 402.8400 ;
      LAYER met3 ;
        RECT 1920.9000 391.3800 1922.5000 391.8600 ;
        RECT 1936.4400 391.3800 1938.0400 391.8600 ;
        RECT 1936.4400 380.5000 1938.0400 380.9800 ;
        RECT 1936.4400 385.9400 1938.0400 386.4200 ;
        RECT 1920.9000 380.5000 1922.5000 380.9800 ;
        RECT 1920.9000 385.9400 1922.5000 386.4200 ;
        RECT 1936.4400 364.1800 1938.0400 364.6600 ;
        RECT 1936.4400 369.6200 1938.0400 370.1000 ;
        RECT 1920.9000 364.1800 1922.5000 364.6600 ;
        RECT 1920.9000 369.6200 1922.5000 370.1000 ;
        RECT 1936.4400 353.3000 1938.0400 353.7800 ;
        RECT 1936.4400 358.7400 1938.0400 359.2200 ;
        RECT 1920.9000 353.3000 1922.5000 353.7800 ;
        RECT 1920.9000 358.7400 1922.5000 359.2200 ;
        RECT 1920.9000 375.0600 1922.5000 375.5400 ;
        RECT 1936.4400 375.0600 1938.0400 375.5400 ;
        RECT 1875.9000 380.5000 1877.5000 380.9800 ;
        RECT 1875.9000 385.9400 1877.5000 386.4200 ;
        RECT 1875.9000 391.3800 1877.5000 391.8600 ;
        RECT 1875.9000 364.1800 1877.5000 364.6600 ;
        RECT 1875.9000 369.6200 1877.5000 370.1000 ;
        RECT 1875.9000 358.7400 1877.5000 359.2200 ;
        RECT 1875.9000 353.3000 1877.5000 353.7800 ;
        RECT 1875.9000 375.0600 1877.5000 375.5400 ;
        RECT 1936.4400 336.9800 1938.0400 337.4600 ;
        RECT 1936.4400 342.4200 1938.0400 342.9000 ;
        RECT 1920.9000 336.9800 1922.5000 337.4600 ;
        RECT 1920.9000 342.4200 1922.5000 342.9000 ;
        RECT 1936.4400 320.6600 1938.0400 321.1400 ;
        RECT 1936.4400 326.1000 1938.0400 326.5800 ;
        RECT 1936.4400 331.5400 1938.0400 332.0200 ;
        RECT 1920.9000 320.6600 1922.5000 321.1400 ;
        RECT 1920.9000 326.1000 1922.5000 326.5800 ;
        RECT 1920.9000 331.5400 1922.5000 332.0200 ;
        RECT 1936.4400 309.7800 1938.0400 310.2600 ;
        RECT 1936.4400 315.2200 1938.0400 315.7000 ;
        RECT 1920.9000 309.7800 1922.5000 310.2600 ;
        RECT 1920.9000 315.2200 1922.5000 315.7000 ;
        RECT 1936.4400 293.4600 1938.0400 293.9400 ;
        RECT 1936.4400 298.9000 1938.0400 299.3800 ;
        RECT 1936.4400 304.3400 1938.0400 304.8200 ;
        RECT 1920.9000 293.4600 1922.5000 293.9400 ;
        RECT 1920.9000 298.9000 1922.5000 299.3800 ;
        RECT 1920.9000 304.3400 1922.5000 304.8200 ;
        RECT 1875.9000 336.9800 1877.5000 337.4600 ;
        RECT 1875.9000 342.4200 1877.5000 342.9000 ;
        RECT 1875.9000 320.6600 1877.5000 321.1400 ;
        RECT 1875.9000 326.1000 1877.5000 326.5800 ;
        RECT 1875.9000 331.5400 1877.5000 332.0200 ;
        RECT 1875.9000 309.7800 1877.5000 310.2600 ;
        RECT 1875.9000 315.2200 1877.5000 315.7000 ;
        RECT 1875.9000 293.4600 1877.5000 293.9400 ;
        RECT 1875.9000 298.9000 1877.5000 299.3800 ;
        RECT 1875.9000 304.3400 1877.5000 304.8200 ;
        RECT 1875.9000 347.8600 1877.5000 348.3400 ;
        RECT 1920.9000 347.8600 1922.5000 348.3400 ;
        RECT 1936.4400 347.8600 1938.0400 348.3400 ;
        RECT 1830.9000 380.5000 1832.5000 380.9800 ;
        RECT 1830.9000 385.9400 1832.5000 386.4200 ;
        RECT 1830.9000 391.3800 1832.5000 391.8600 ;
        RECT 1785.9000 380.5000 1787.5000 380.9800 ;
        RECT 1785.9000 385.9400 1787.5000 386.4200 ;
        RECT 1785.9000 391.3800 1787.5000 391.8600 ;
        RECT 1830.9000 364.1800 1832.5000 364.6600 ;
        RECT 1830.9000 369.6200 1832.5000 370.1000 ;
        RECT 1830.9000 353.3000 1832.5000 353.7800 ;
        RECT 1830.9000 358.7400 1832.5000 359.2200 ;
        RECT 1785.9000 364.1800 1787.5000 364.6600 ;
        RECT 1785.9000 369.6200 1787.5000 370.1000 ;
        RECT 1785.9000 353.3000 1787.5000 353.7800 ;
        RECT 1785.9000 358.7400 1787.5000 359.2200 ;
        RECT 1785.9000 375.0600 1787.5000 375.5400 ;
        RECT 1830.9000 375.0600 1832.5000 375.5400 ;
        RECT 1733.7400 391.3800 1735.3400 391.8600 ;
        RECT 1740.9000 391.3800 1742.5000 391.8600 ;
        RECT 1740.9000 380.5000 1742.5000 380.9800 ;
        RECT 1740.9000 385.9400 1742.5000 386.4200 ;
        RECT 1733.7400 380.5000 1735.3400 380.9800 ;
        RECT 1733.7400 385.9400 1735.3400 386.4200 ;
        RECT 1740.9000 364.1800 1742.5000 364.6600 ;
        RECT 1740.9000 369.6200 1742.5000 370.1000 ;
        RECT 1733.7400 364.1800 1735.3400 364.6600 ;
        RECT 1733.7400 369.6200 1735.3400 370.1000 ;
        RECT 1740.9000 353.3000 1742.5000 353.7800 ;
        RECT 1740.9000 358.7400 1742.5000 359.2200 ;
        RECT 1733.7400 353.3000 1735.3400 353.7800 ;
        RECT 1733.7400 358.7400 1735.3400 359.2200 ;
        RECT 1733.7400 375.0600 1735.3400 375.5400 ;
        RECT 1740.9000 375.0600 1742.5000 375.5400 ;
        RECT 1830.9000 336.9800 1832.5000 337.4600 ;
        RECT 1830.9000 342.4200 1832.5000 342.9000 ;
        RECT 1830.9000 320.6600 1832.5000 321.1400 ;
        RECT 1830.9000 326.1000 1832.5000 326.5800 ;
        RECT 1830.9000 331.5400 1832.5000 332.0200 ;
        RECT 1785.9000 336.9800 1787.5000 337.4600 ;
        RECT 1785.9000 342.4200 1787.5000 342.9000 ;
        RECT 1785.9000 320.6600 1787.5000 321.1400 ;
        RECT 1785.9000 326.1000 1787.5000 326.5800 ;
        RECT 1785.9000 331.5400 1787.5000 332.0200 ;
        RECT 1830.9000 309.7800 1832.5000 310.2600 ;
        RECT 1830.9000 315.2200 1832.5000 315.7000 ;
        RECT 1830.9000 293.4600 1832.5000 293.9400 ;
        RECT 1830.9000 298.9000 1832.5000 299.3800 ;
        RECT 1830.9000 304.3400 1832.5000 304.8200 ;
        RECT 1785.9000 309.7800 1787.5000 310.2600 ;
        RECT 1785.9000 315.2200 1787.5000 315.7000 ;
        RECT 1785.9000 293.4600 1787.5000 293.9400 ;
        RECT 1785.9000 298.9000 1787.5000 299.3800 ;
        RECT 1785.9000 304.3400 1787.5000 304.8200 ;
        RECT 1740.9000 336.9800 1742.5000 337.4600 ;
        RECT 1740.9000 342.4200 1742.5000 342.9000 ;
        RECT 1733.7400 336.9800 1735.3400 337.4600 ;
        RECT 1733.7400 342.4200 1735.3400 342.9000 ;
        RECT 1740.9000 320.6600 1742.5000 321.1400 ;
        RECT 1740.9000 326.1000 1742.5000 326.5800 ;
        RECT 1740.9000 331.5400 1742.5000 332.0200 ;
        RECT 1733.7400 320.6600 1735.3400 321.1400 ;
        RECT 1733.7400 326.1000 1735.3400 326.5800 ;
        RECT 1733.7400 331.5400 1735.3400 332.0200 ;
        RECT 1740.9000 309.7800 1742.5000 310.2600 ;
        RECT 1740.9000 315.2200 1742.5000 315.7000 ;
        RECT 1733.7400 309.7800 1735.3400 310.2600 ;
        RECT 1733.7400 315.2200 1735.3400 315.7000 ;
        RECT 1740.9000 293.4600 1742.5000 293.9400 ;
        RECT 1740.9000 298.9000 1742.5000 299.3800 ;
        RECT 1740.9000 304.3400 1742.5000 304.8200 ;
        RECT 1733.7400 293.4600 1735.3400 293.9400 ;
        RECT 1733.7400 298.9000 1735.3400 299.3800 ;
        RECT 1733.7400 304.3400 1735.3400 304.8200 ;
        RECT 1733.7400 347.8600 1735.3400 348.3400 ;
        RECT 1740.9000 347.8600 1742.5000 348.3400 ;
        RECT 1785.9000 347.8600 1787.5000 348.3400 ;
        RECT 1830.9000 347.8600 1832.5000 348.3400 ;
        RECT 1936.4400 282.5800 1938.0400 283.0600 ;
        RECT 1936.4400 288.0200 1938.0400 288.5000 ;
        RECT 1920.9000 282.5800 1922.5000 283.0600 ;
        RECT 1920.9000 288.0200 1922.5000 288.5000 ;
        RECT 1936.4400 266.2600 1938.0400 266.7400 ;
        RECT 1936.4400 271.7000 1938.0400 272.1800 ;
        RECT 1936.4400 277.1400 1938.0400 277.6200 ;
        RECT 1920.9000 266.2600 1922.5000 266.7400 ;
        RECT 1920.9000 271.7000 1922.5000 272.1800 ;
        RECT 1920.9000 277.1400 1922.5000 277.6200 ;
        RECT 1936.4400 255.3800 1938.0400 255.8600 ;
        RECT 1936.4400 260.8200 1938.0400 261.3000 ;
        RECT 1920.9000 255.3800 1922.5000 255.8600 ;
        RECT 1920.9000 260.8200 1922.5000 261.3000 ;
        RECT 1936.4400 239.0600 1938.0400 239.5400 ;
        RECT 1936.4400 244.5000 1938.0400 244.9800 ;
        RECT 1936.4400 249.9400 1938.0400 250.4200 ;
        RECT 1920.9000 239.0600 1922.5000 239.5400 ;
        RECT 1920.9000 244.5000 1922.5000 244.9800 ;
        RECT 1920.9000 249.9400 1922.5000 250.4200 ;
        RECT 1875.9000 282.5800 1877.5000 283.0600 ;
        RECT 1875.9000 288.0200 1877.5000 288.5000 ;
        RECT 1875.9000 266.2600 1877.5000 266.7400 ;
        RECT 1875.9000 271.7000 1877.5000 272.1800 ;
        RECT 1875.9000 277.1400 1877.5000 277.6200 ;
        RECT 1875.9000 255.3800 1877.5000 255.8600 ;
        RECT 1875.9000 260.8200 1877.5000 261.3000 ;
        RECT 1875.9000 239.0600 1877.5000 239.5400 ;
        RECT 1875.9000 244.5000 1877.5000 244.9800 ;
        RECT 1875.9000 249.9400 1877.5000 250.4200 ;
        RECT 1936.4400 228.1800 1938.0400 228.6600 ;
        RECT 1936.4400 233.6200 1938.0400 234.1000 ;
        RECT 1920.9000 228.1800 1922.5000 228.6600 ;
        RECT 1920.9000 233.6200 1922.5000 234.1000 ;
        RECT 1936.4400 211.8600 1938.0400 212.3400 ;
        RECT 1936.4400 217.3000 1938.0400 217.7800 ;
        RECT 1936.4400 222.7400 1938.0400 223.2200 ;
        RECT 1920.9000 211.8600 1922.5000 212.3400 ;
        RECT 1920.9000 217.3000 1922.5000 217.7800 ;
        RECT 1920.9000 222.7400 1922.5000 223.2200 ;
        RECT 1936.4400 200.9800 1938.0400 201.4600 ;
        RECT 1936.4400 206.4200 1938.0400 206.9000 ;
        RECT 1920.9000 200.9800 1922.5000 201.4600 ;
        RECT 1920.9000 206.4200 1922.5000 206.9000 ;
        RECT 1920.9000 195.5400 1922.5000 196.0200 ;
        RECT 1936.4400 195.5400 1938.0400 196.0200 ;
        RECT 1875.9000 228.1800 1877.5000 228.6600 ;
        RECT 1875.9000 233.6200 1877.5000 234.1000 ;
        RECT 1875.9000 211.8600 1877.5000 212.3400 ;
        RECT 1875.9000 217.3000 1877.5000 217.7800 ;
        RECT 1875.9000 222.7400 1877.5000 223.2200 ;
        RECT 1875.9000 200.9800 1877.5000 201.4600 ;
        RECT 1875.9000 206.4200 1877.5000 206.9000 ;
        RECT 1875.9000 195.5400 1877.5000 196.0200 ;
        RECT 1830.9000 282.5800 1832.5000 283.0600 ;
        RECT 1830.9000 288.0200 1832.5000 288.5000 ;
        RECT 1830.9000 266.2600 1832.5000 266.7400 ;
        RECT 1830.9000 271.7000 1832.5000 272.1800 ;
        RECT 1830.9000 277.1400 1832.5000 277.6200 ;
        RECT 1785.9000 282.5800 1787.5000 283.0600 ;
        RECT 1785.9000 288.0200 1787.5000 288.5000 ;
        RECT 1785.9000 266.2600 1787.5000 266.7400 ;
        RECT 1785.9000 271.7000 1787.5000 272.1800 ;
        RECT 1785.9000 277.1400 1787.5000 277.6200 ;
        RECT 1830.9000 255.3800 1832.5000 255.8600 ;
        RECT 1830.9000 260.8200 1832.5000 261.3000 ;
        RECT 1830.9000 239.0600 1832.5000 239.5400 ;
        RECT 1830.9000 244.5000 1832.5000 244.9800 ;
        RECT 1830.9000 249.9400 1832.5000 250.4200 ;
        RECT 1785.9000 255.3800 1787.5000 255.8600 ;
        RECT 1785.9000 260.8200 1787.5000 261.3000 ;
        RECT 1785.9000 239.0600 1787.5000 239.5400 ;
        RECT 1785.9000 244.5000 1787.5000 244.9800 ;
        RECT 1785.9000 249.9400 1787.5000 250.4200 ;
        RECT 1740.9000 282.5800 1742.5000 283.0600 ;
        RECT 1740.9000 288.0200 1742.5000 288.5000 ;
        RECT 1733.7400 282.5800 1735.3400 283.0600 ;
        RECT 1733.7400 288.0200 1735.3400 288.5000 ;
        RECT 1740.9000 266.2600 1742.5000 266.7400 ;
        RECT 1740.9000 271.7000 1742.5000 272.1800 ;
        RECT 1740.9000 277.1400 1742.5000 277.6200 ;
        RECT 1733.7400 266.2600 1735.3400 266.7400 ;
        RECT 1733.7400 271.7000 1735.3400 272.1800 ;
        RECT 1733.7400 277.1400 1735.3400 277.6200 ;
        RECT 1740.9000 255.3800 1742.5000 255.8600 ;
        RECT 1740.9000 260.8200 1742.5000 261.3000 ;
        RECT 1733.7400 255.3800 1735.3400 255.8600 ;
        RECT 1733.7400 260.8200 1735.3400 261.3000 ;
        RECT 1740.9000 239.0600 1742.5000 239.5400 ;
        RECT 1740.9000 244.5000 1742.5000 244.9800 ;
        RECT 1740.9000 249.9400 1742.5000 250.4200 ;
        RECT 1733.7400 239.0600 1735.3400 239.5400 ;
        RECT 1733.7400 244.5000 1735.3400 244.9800 ;
        RECT 1733.7400 249.9400 1735.3400 250.4200 ;
        RECT 1830.9000 228.1800 1832.5000 228.6600 ;
        RECT 1830.9000 233.6200 1832.5000 234.1000 ;
        RECT 1830.9000 211.8600 1832.5000 212.3400 ;
        RECT 1830.9000 217.3000 1832.5000 217.7800 ;
        RECT 1830.9000 222.7400 1832.5000 223.2200 ;
        RECT 1785.9000 228.1800 1787.5000 228.6600 ;
        RECT 1785.9000 233.6200 1787.5000 234.1000 ;
        RECT 1785.9000 211.8600 1787.5000 212.3400 ;
        RECT 1785.9000 217.3000 1787.5000 217.7800 ;
        RECT 1785.9000 222.7400 1787.5000 223.2200 ;
        RECT 1830.9000 206.4200 1832.5000 206.9000 ;
        RECT 1830.9000 200.9800 1832.5000 201.4600 ;
        RECT 1830.9000 195.5400 1832.5000 196.0200 ;
        RECT 1785.9000 206.4200 1787.5000 206.9000 ;
        RECT 1785.9000 200.9800 1787.5000 201.4600 ;
        RECT 1785.9000 195.5400 1787.5000 196.0200 ;
        RECT 1740.9000 228.1800 1742.5000 228.6600 ;
        RECT 1740.9000 233.6200 1742.5000 234.1000 ;
        RECT 1733.7400 228.1800 1735.3400 228.6600 ;
        RECT 1733.7400 233.6200 1735.3400 234.1000 ;
        RECT 1740.9000 211.8600 1742.5000 212.3400 ;
        RECT 1740.9000 217.3000 1742.5000 217.7800 ;
        RECT 1740.9000 222.7400 1742.5000 223.2200 ;
        RECT 1733.7400 211.8600 1735.3400 212.3400 ;
        RECT 1733.7400 217.3000 1735.3400 217.7800 ;
        RECT 1733.7400 222.7400 1735.3400 223.2200 ;
        RECT 1740.9000 200.9800 1742.5000 201.4600 ;
        RECT 1740.9000 206.4200 1742.5000 206.9000 ;
        RECT 1733.7400 200.9800 1735.3400 201.4600 ;
        RECT 1733.7400 206.4200 1735.3400 206.9000 ;
        RECT 1733.7400 195.5400 1735.3400 196.0200 ;
        RECT 1740.9000 195.5400 1742.5000 196.0200 ;
        RECT 1730.7800 397.7300 1941.0000 399.3300 ;
        RECT 1730.7800 186.0300 1941.0000 187.6300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 183.2000 1735.3400 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 401.2400 1735.3400 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 183.2000 1938.0400 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 401.2400 1938.0400 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 186.0300 1732.3800 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 186.0300 1941.0000 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 397.7300 1732.3800 399.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 397.7300 1941.0000 399.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1733.8400 142.9400 1735.4400 173.2000 ;
        RECT 1936.3400 142.9400 1937.9400 173.2000 ;
      LAYER met3 ;
        RECT 1936.3400 163.4400 1937.9400 163.9200 ;
        RECT 1733.8400 163.4400 1735.4400 163.9200 ;
        RECT 1936.3400 152.5600 1937.9400 153.0400 ;
        RECT 1733.8400 152.5600 1735.4400 153.0400 ;
        RECT 1936.3400 158.0000 1937.9400 158.4800 ;
        RECT 1733.8400 158.0000 1735.4400 158.4800 ;
        RECT 1730.7800 168.8400 1941.0000 170.4400 ;
        RECT 1730.7800 144.5100 1941.0000 146.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.8400 142.9400 1735.4400 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.8400 171.6000 1735.4400 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.3400 142.9400 1937.9400 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.3400 171.6000 1937.9400 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 144.5100 1732.3800 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 144.5100 1941.0000 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 168.8400 1732.3800 170.4400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 168.8400 1941.0000 170.4400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 2252.7900 1922.5000 2466.0900 ;
        RECT 1875.9000 2252.7900 1877.5000 2466.0900 ;
        RECT 1830.9000 2252.7900 1832.5000 2466.0900 ;
        RECT 1785.9000 2252.7900 1787.5000 2466.0900 ;
        RECT 1740.9000 2252.7900 1742.5000 2466.0900 ;
        RECT 1936.4400 2249.9600 1938.0400 2469.6000 ;
        RECT 1733.7400 2249.9600 1735.3400 2469.6000 ;
      LAYER met3 ;
        RECT 1920.9000 2458.1400 1922.5000 2458.6200 ;
        RECT 1936.4400 2458.1400 1938.0400 2458.6200 ;
        RECT 1936.4400 2447.2600 1938.0400 2447.7400 ;
        RECT 1936.4400 2452.7000 1938.0400 2453.1800 ;
        RECT 1920.9000 2447.2600 1922.5000 2447.7400 ;
        RECT 1920.9000 2452.7000 1922.5000 2453.1800 ;
        RECT 1936.4400 2430.9400 1938.0400 2431.4200 ;
        RECT 1936.4400 2436.3800 1938.0400 2436.8600 ;
        RECT 1920.9000 2430.9400 1922.5000 2431.4200 ;
        RECT 1920.9000 2436.3800 1922.5000 2436.8600 ;
        RECT 1936.4400 2420.0600 1938.0400 2420.5400 ;
        RECT 1936.4400 2425.5000 1938.0400 2425.9800 ;
        RECT 1920.9000 2420.0600 1922.5000 2420.5400 ;
        RECT 1920.9000 2425.5000 1922.5000 2425.9800 ;
        RECT 1920.9000 2441.8200 1922.5000 2442.3000 ;
        RECT 1936.4400 2441.8200 1938.0400 2442.3000 ;
        RECT 1875.9000 2447.2600 1877.5000 2447.7400 ;
        RECT 1875.9000 2452.7000 1877.5000 2453.1800 ;
        RECT 1875.9000 2458.1400 1877.5000 2458.6200 ;
        RECT 1875.9000 2430.9400 1877.5000 2431.4200 ;
        RECT 1875.9000 2436.3800 1877.5000 2436.8600 ;
        RECT 1875.9000 2425.5000 1877.5000 2425.9800 ;
        RECT 1875.9000 2420.0600 1877.5000 2420.5400 ;
        RECT 1875.9000 2441.8200 1877.5000 2442.3000 ;
        RECT 1936.4400 2403.7400 1938.0400 2404.2200 ;
        RECT 1936.4400 2409.1800 1938.0400 2409.6600 ;
        RECT 1920.9000 2403.7400 1922.5000 2404.2200 ;
        RECT 1920.9000 2409.1800 1922.5000 2409.6600 ;
        RECT 1936.4400 2387.4200 1938.0400 2387.9000 ;
        RECT 1936.4400 2392.8600 1938.0400 2393.3400 ;
        RECT 1936.4400 2398.3000 1938.0400 2398.7800 ;
        RECT 1920.9000 2387.4200 1922.5000 2387.9000 ;
        RECT 1920.9000 2392.8600 1922.5000 2393.3400 ;
        RECT 1920.9000 2398.3000 1922.5000 2398.7800 ;
        RECT 1936.4400 2376.5400 1938.0400 2377.0200 ;
        RECT 1936.4400 2381.9800 1938.0400 2382.4600 ;
        RECT 1920.9000 2376.5400 1922.5000 2377.0200 ;
        RECT 1920.9000 2381.9800 1922.5000 2382.4600 ;
        RECT 1936.4400 2360.2200 1938.0400 2360.7000 ;
        RECT 1936.4400 2365.6600 1938.0400 2366.1400 ;
        RECT 1936.4400 2371.1000 1938.0400 2371.5800 ;
        RECT 1920.9000 2360.2200 1922.5000 2360.7000 ;
        RECT 1920.9000 2365.6600 1922.5000 2366.1400 ;
        RECT 1920.9000 2371.1000 1922.5000 2371.5800 ;
        RECT 1875.9000 2403.7400 1877.5000 2404.2200 ;
        RECT 1875.9000 2409.1800 1877.5000 2409.6600 ;
        RECT 1875.9000 2387.4200 1877.5000 2387.9000 ;
        RECT 1875.9000 2392.8600 1877.5000 2393.3400 ;
        RECT 1875.9000 2398.3000 1877.5000 2398.7800 ;
        RECT 1875.9000 2376.5400 1877.5000 2377.0200 ;
        RECT 1875.9000 2381.9800 1877.5000 2382.4600 ;
        RECT 1875.9000 2360.2200 1877.5000 2360.7000 ;
        RECT 1875.9000 2365.6600 1877.5000 2366.1400 ;
        RECT 1875.9000 2371.1000 1877.5000 2371.5800 ;
        RECT 1875.9000 2414.6200 1877.5000 2415.1000 ;
        RECT 1920.9000 2414.6200 1922.5000 2415.1000 ;
        RECT 1936.4400 2414.6200 1938.0400 2415.1000 ;
        RECT 1830.9000 2447.2600 1832.5000 2447.7400 ;
        RECT 1830.9000 2452.7000 1832.5000 2453.1800 ;
        RECT 1830.9000 2458.1400 1832.5000 2458.6200 ;
        RECT 1785.9000 2447.2600 1787.5000 2447.7400 ;
        RECT 1785.9000 2452.7000 1787.5000 2453.1800 ;
        RECT 1785.9000 2458.1400 1787.5000 2458.6200 ;
        RECT 1830.9000 2430.9400 1832.5000 2431.4200 ;
        RECT 1830.9000 2436.3800 1832.5000 2436.8600 ;
        RECT 1830.9000 2420.0600 1832.5000 2420.5400 ;
        RECT 1830.9000 2425.5000 1832.5000 2425.9800 ;
        RECT 1785.9000 2430.9400 1787.5000 2431.4200 ;
        RECT 1785.9000 2436.3800 1787.5000 2436.8600 ;
        RECT 1785.9000 2420.0600 1787.5000 2420.5400 ;
        RECT 1785.9000 2425.5000 1787.5000 2425.9800 ;
        RECT 1785.9000 2441.8200 1787.5000 2442.3000 ;
        RECT 1830.9000 2441.8200 1832.5000 2442.3000 ;
        RECT 1733.7400 2458.1400 1735.3400 2458.6200 ;
        RECT 1740.9000 2458.1400 1742.5000 2458.6200 ;
        RECT 1740.9000 2447.2600 1742.5000 2447.7400 ;
        RECT 1740.9000 2452.7000 1742.5000 2453.1800 ;
        RECT 1733.7400 2447.2600 1735.3400 2447.7400 ;
        RECT 1733.7400 2452.7000 1735.3400 2453.1800 ;
        RECT 1740.9000 2430.9400 1742.5000 2431.4200 ;
        RECT 1740.9000 2436.3800 1742.5000 2436.8600 ;
        RECT 1733.7400 2430.9400 1735.3400 2431.4200 ;
        RECT 1733.7400 2436.3800 1735.3400 2436.8600 ;
        RECT 1740.9000 2420.0600 1742.5000 2420.5400 ;
        RECT 1740.9000 2425.5000 1742.5000 2425.9800 ;
        RECT 1733.7400 2420.0600 1735.3400 2420.5400 ;
        RECT 1733.7400 2425.5000 1735.3400 2425.9800 ;
        RECT 1733.7400 2441.8200 1735.3400 2442.3000 ;
        RECT 1740.9000 2441.8200 1742.5000 2442.3000 ;
        RECT 1830.9000 2403.7400 1832.5000 2404.2200 ;
        RECT 1830.9000 2409.1800 1832.5000 2409.6600 ;
        RECT 1830.9000 2387.4200 1832.5000 2387.9000 ;
        RECT 1830.9000 2392.8600 1832.5000 2393.3400 ;
        RECT 1830.9000 2398.3000 1832.5000 2398.7800 ;
        RECT 1785.9000 2403.7400 1787.5000 2404.2200 ;
        RECT 1785.9000 2409.1800 1787.5000 2409.6600 ;
        RECT 1785.9000 2387.4200 1787.5000 2387.9000 ;
        RECT 1785.9000 2392.8600 1787.5000 2393.3400 ;
        RECT 1785.9000 2398.3000 1787.5000 2398.7800 ;
        RECT 1830.9000 2376.5400 1832.5000 2377.0200 ;
        RECT 1830.9000 2381.9800 1832.5000 2382.4600 ;
        RECT 1830.9000 2360.2200 1832.5000 2360.7000 ;
        RECT 1830.9000 2365.6600 1832.5000 2366.1400 ;
        RECT 1830.9000 2371.1000 1832.5000 2371.5800 ;
        RECT 1785.9000 2376.5400 1787.5000 2377.0200 ;
        RECT 1785.9000 2381.9800 1787.5000 2382.4600 ;
        RECT 1785.9000 2360.2200 1787.5000 2360.7000 ;
        RECT 1785.9000 2365.6600 1787.5000 2366.1400 ;
        RECT 1785.9000 2371.1000 1787.5000 2371.5800 ;
        RECT 1740.9000 2403.7400 1742.5000 2404.2200 ;
        RECT 1740.9000 2409.1800 1742.5000 2409.6600 ;
        RECT 1733.7400 2403.7400 1735.3400 2404.2200 ;
        RECT 1733.7400 2409.1800 1735.3400 2409.6600 ;
        RECT 1740.9000 2387.4200 1742.5000 2387.9000 ;
        RECT 1740.9000 2392.8600 1742.5000 2393.3400 ;
        RECT 1740.9000 2398.3000 1742.5000 2398.7800 ;
        RECT 1733.7400 2387.4200 1735.3400 2387.9000 ;
        RECT 1733.7400 2392.8600 1735.3400 2393.3400 ;
        RECT 1733.7400 2398.3000 1735.3400 2398.7800 ;
        RECT 1740.9000 2376.5400 1742.5000 2377.0200 ;
        RECT 1740.9000 2381.9800 1742.5000 2382.4600 ;
        RECT 1733.7400 2376.5400 1735.3400 2377.0200 ;
        RECT 1733.7400 2381.9800 1735.3400 2382.4600 ;
        RECT 1740.9000 2360.2200 1742.5000 2360.7000 ;
        RECT 1740.9000 2365.6600 1742.5000 2366.1400 ;
        RECT 1740.9000 2371.1000 1742.5000 2371.5800 ;
        RECT 1733.7400 2360.2200 1735.3400 2360.7000 ;
        RECT 1733.7400 2365.6600 1735.3400 2366.1400 ;
        RECT 1733.7400 2371.1000 1735.3400 2371.5800 ;
        RECT 1733.7400 2414.6200 1735.3400 2415.1000 ;
        RECT 1740.9000 2414.6200 1742.5000 2415.1000 ;
        RECT 1785.9000 2414.6200 1787.5000 2415.1000 ;
        RECT 1830.9000 2414.6200 1832.5000 2415.1000 ;
        RECT 1936.4400 2349.3400 1938.0400 2349.8200 ;
        RECT 1936.4400 2354.7800 1938.0400 2355.2600 ;
        RECT 1920.9000 2349.3400 1922.5000 2349.8200 ;
        RECT 1920.9000 2354.7800 1922.5000 2355.2600 ;
        RECT 1936.4400 2333.0200 1938.0400 2333.5000 ;
        RECT 1936.4400 2338.4600 1938.0400 2338.9400 ;
        RECT 1936.4400 2343.9000 1938.0400 2344.3800 ;
        RECT 1920.9000 2333.0200 1922.5000 2333.5000 ;
        RECT 1920.9000 2338.4600 1922.5000 2338.9400 ;
        RECT 1920.9000 2343.9000 1922.5000 2344.3800 ;
        RECT 1936.4400 2322.1400 1938.0400 2322.6200 ;
        RECT 1936.4400 2327.5800 1938.0400 2328.0600 ;
        RECT 1920.9000 2322.1400 1922.5000 2322.6200 ;
        RECT 1920.9000 2327.5800 1922.5000 2328.0600 ;
        RECT 1936.4400 2305.8200 1938.0400 2306.3000 ;
        RECT 1936.4400 2311.2600 1938.0400 2311.7400 ;
        RECT 1936.4400 2316.7000 1938.0400 2317.1800 ;
        RECT 1920.9000 2305.8200 1922.5000 2306.3000 ;
        RECT 1920.9000 2311.2600 1922.5000 2311.7400 ;
        RECT 1920.9000 2316.7000 1922.5000 2317.1800 ;
        RECT 1875.9000 2349.3400 1877.5000 2349.8200 ;
        RECT 1875.9000 2354.7800 1877.5000 2355.2600 ;
        RECT 1875.9000 2333.0200 1877.5000 2333.5000 ;
        RECT 1875.9000 2338.4600 1877.5000 2338.9400 ;
        RECT 1875.9000 2343.9000 1877.5000 2344.3800 ;
        RECT 1875.9000 2322.1400 1877.5000 2322.6200 ;
        RECT 1875.9000 2327.5800 1877.5000 2328.0600 ;
        RECT 1875.9000 2305.8200 1877.5000 2306.3000 ;
        RECT 1875.9000 2311.2600 1877.5000 2311.7400 ;
        RECT 1875.9000 2316.7000 1877.5000 2317.1800 ;
        RECT 1936.4400 2294.9400 1938.0400 2295.4200 ;
        RECT 1936.4400 2300.3800 1938.0400 2300.8600 ;
        RECT 1920.9000 2294.9400 1922.5000 2295.4200 ;
        RECT 1920.9000 2300.3800 1922.5000 2300.8600 ;
        RECT 1936.4400 2278.6200 1938.0400 2279.1000 ;
        RECT 1936.4400 2284.0600 1938.0400 2284.5400 ;
        RECT 1936.4400 2289.5000 1938.0400 2289.9800 ;
        RECT 1920.9000 2278.6200 1922.5000 2279.1000 ;
        RECT 1920.9000 2284.0600 1922.5000 2284.5400 ;
        RECT 1920.9000 2289.5000 1922.5000 2289.9800 ;
        RECT 1936.4400 2267.7400 1938.0400 2268.2200 ;
        RECT 1936.4400 2273.1800 1938.0400 2273.6600 ;
        RECT 1920.9000 2267.7400 1922.5000 2268.2200 ;
        RECT 1920.9000 2273.1800 1922.5000 2273.6600 ;
        RECT 1920.9000 2262.3000 1922.5000 2262.7800 ;
        RECT 1936.4400 2262.3000 1938.0400 2262.7800 ;
        RECT 1875.9000 2294.9400 1877.5000 2295.4200 ;
        RECT 1875.9000 2300.3800 1877.5000 2300.8600 ;
        RECT 1875.9000 2278.6200 1877.5000 2279.1000 ;
        RECT 1875.9000 2284.0600 1877.5000 2284.5400 ;
        RECT 1875.9000 2289.5000 1877.5000 2289.9800 ;
        RECT 1875.9000 2267.7400 1877.5000 2268.2200 ;
        RECT 1875.9000 2273.1800 1877.5000 2273.6600 ;
        RECT 1875.9000 2262.3000 1877.5000 2262.7800 ;
        RECT 1830.9000 2349.3400 1832.5000 2349.8200 ;
        RECT 1830.9000 2354.7800 1832.5000 2355.2600 ;
        RECT 1830.9000 2333.0200 1832.5000 2333.5000 ;
        RECT 1830.9000 2338.4600 1832.5000 2338.9400 ;
        RECT 1830.9000 2343.9000 1832.5000 2344.3800 ;
        RECT 1785.9000 2349.3400 1787.5000 2349.8200 ;
        RECT 1785.9000 2354.7800 1787.5000 2355.2600 ;
        RECT 1785.9000 2333.0200 1787.5000 2333.5000 ;
        RECT 1785.9000 2338.4600 1787.5000 2338.9400 ;
        RECT 1785.9000 2343.9000 1787.5000 2344.3800 ;
        RECT 1830.9000 2322.1400 1832.5000 2322.6200 ;
        RECT 1830.9000 2327.5800 1832.5000 2328.0600 ;
        RECT 1830.9000 2305.8200 1832.5000 2306.3000 ;
        RECT 1830.9000 2311.2600 1832.5000 2311.7400 ;
        RECT 1830.9000 2316.7000 1832.5000 2317.1800 ;
        RECT 1785.9000 2322.1400 1787.5000 2322.6200 ;
        RECT 1785.9000 2327.5800 1787.5000 2328.0600 ;
        RECT 1785.9000 2305.8200 1787.5000 2306.3000 ;
        RECT 1785.9000 2311.2600 1787.5000 2311.7400 ;
        RECT 1785.9000 2316.7000 1787.5000 2317.1800 ;
        RECT 1740.9000 2349.3400 1742.5000 2349.8200 ;
        RECT 1740.9000 2354.7800 1742.5000 2355.2600 ;
        RECT 1733.7400 2349.3400 1735.3400 2349.8200 ;
        RECT 1733.7400 2354.7800 1735.3400 2355.2600 ;
        RECT 1740.9000 2333.0200 1742.5000 2333.5000 ;
        RECT 1740.9000 2338.4600 1742.5000 2338.9400 ;
        RECT 1740.9000 2343.9000 1742.5000 2344.3800 ;
        RECT 1733.7400 2333.0200 1735.3400 2333.5000 ;
        RECT 1733.7400 2338.4600 1735.3400 2338.9400 ;
        RECT 1733.7400 2343.9000 1735.3400 2344.3800 ;
        RECT 1740.9000 2322.1400 1742.5000 2322.6200 ;
        RECT 1740.9000 2327.5800 1742.5000 2328.0600 ;
        RECT 1733.7400 2322.1400 1735.3400 2322.6200 ;
        RECT 1733.7400 2327.5800 1735.3400 2328.0600 ;
        RECT 1740.9000 2305.8200 1742.5000 2306.3000 ;
        RECT 1740.9000 2311.2600 1742.5000 2311.7400 ;
        RECT 1740.9000 2316.7000 1742.5000 2317.1800 ;
        RECT 1733.7400 2305.8200 1735.3400 2306.3000 ;
        RECT 1733.7400 2311.2600 1735.3400 2311.7400 ;
        RECT 1733.7400 2316.7000 1735.3400 2317.1800 ;
        RECT 1830.9000 2294.9400 1832.5000 2295.4200 ;
        RECT 1830.9000 2300.3800 1832.5000 2300.8600 ;
        RECT 1830.9000 2278.6200 1832.5000 2279.1000 ;
        RECT 1830.9000 2284.0600 1832.5000 2284.5400 ;
        RECT 1830.9000 2289.5000 1832.5000 2289.9800 ;
        RECT 1785.9000 2294.9400 1787.5000 2295.4200 ;
        RECT 1785.9000 2300.3800 1787.5000 2300.8600 ;
        RECT 1785.9000 2278.6200 1787.5000 2279.1000 ;
        RECT 1785.9000 2284.0600 1787.5000 2284.5400 ;
        RECT 1785.9000 2289.5000 1787.5000 2289.9800 ;
        RECT 1830.9000 2273.1800 1832.5000 2273.6600 ;
        RECT 1830.9000 2267.7400 1832.5000 2268.2200 ;
        RECT 1830.9000 2262.3000 1832.5000 2262.7800 ;
        RECT 1785.9000 2273.1800 1787.5000 2273.6600 ;
        RECT 1785.9000 2267.7400 1787.5000 2268.2200 ;
        RECT 1785.9000 2262.3000 1787.5000 2262.7800 ;
        RECT 1740.9000 2294.9400 1742.5000 2295.4200 ;
        RECT 1740.9000 2300.3800 1742.5000 2300.8600 ;
        RECT 1733.7400 2294.9400 1735.3400 2295.4200 ;
        RECT 1733.7400 2300.3800 1735.3400 2300.8600 ;
        RECT 1740.9000 2278.6200 1742.5000 2279.1000 ;
        RECT 1740.9000 2284.0600 1742.5000 2284.5400 ;
        RECT 1740.9000 2289.5000 1742.5000 2289.9800 ;
        RECT 1733.7400 2278.6200 1735.3400 2279.1000 ;
        RECT 1733.7400 2284.0600 1735.3400 2284.5400 ;
        RECT 1733.7400 2289.5000 1735.3400 2289.9800 ;
        RECT 1740.9000 2267.7400 1742.5000 2268.2200 ;
        RECT 1740.9000 2273.1800 1742.5000 2273.6600 ;
        RECT 1733.7400 2267.7400 1735.3400 2268.2200 ;
        RECT 1733.7400 2273.1800 1735.3400 2273.6600 ;
        RECT 1733.7400 2262.3000 1735.3400 2262.7800 ;
        RECT 1740.9000 2262.3000 1742.5000 2262.7800 ;
        RECT 1730.7800 2464.4900 1941.0000 2466.0900 ;
        RECT 1730.7800 2252.7900 1941.0000 2254.3900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 2249.9600 1735.3400 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 2468.0000 1735.3400 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 2249.9600 1938.0400 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 2468.0000 1938.0400 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2252.7900 1732.3800 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2252.7900 1941.0000 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2464.4900 1732.3800 2466.0900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2464.4900 1941.0000 2466.0900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 2023.1500 1922.5000 2236.4500 ;
        RECT 1875.9000 2023.1500 1877.5000 2236.4500 ;
        RECT 1830.9000 2023.1500 1832.5000 2236.4500 ;
        RECT 1785.9000 2023.1500 1787.5000 2236.4500 ;
        RECT 1740.9000 2023.1500 1742.5000 2236.4500 ;
        RECT 1936.4400 2020.3200 1938.0400 2239.9600 ;
        RECT 1733.7400 2020.3200 1735.3400 2239.9600 ;
      LAYER met3 ;
        RECT 1920.9000 2228.5000 1922.5000 2228.9800 ;
        RECT 1936.4400 2228.5000 1938.0400 2228.9800 ;
        RECT 1936.4400 2217.6200 1938.0400 2218.1000 ;
        RECT 1936.4400 2223.0600 1938.0400 2223.5400 ;
        RECT 1920.9000 2217.6200 1922.5000 2218.1000 ;
        RECT 1920.9000 2223.0600 1922.5000 2223.5400 ;
        RECT 1936.4400 2201.3000 1938.0400 2201.7800 ;
        RECT 1936.4400 2206.7400 1938.0400 2207.2200 ;
        RECT 1920.9000 2201.3000 1922.5000 2201.7800 ;
        RECT 1920.9000 2206.7400 1922.5000 2207.2200 ;
        RECT 1936.4400 2190.4200 1938.0400 2190.9000 ;
        RECT 1936.4400 2195.8600 1938.0400 2196.3400 ;
        RECT 1920.9000 2190.4200 1922.5000 2190.9000 ;
        RECT 1920.9000 2195.8600 1922.5000 2196.3400 ;
        RECT 1920.9000 2212.1800 1922.5000 2212.6600 ;
        RECT 1936.4400 2212.1800 1938.0400 2212.6600 ;
        RECT 1875.9000 2217.6200 1877.5000 2218.1000 ;
        RECT 1875.9000 2223.0600 1877.5000 2223.5400 ;
        RECT 1875.9000 2228.5000 1877.5000 2228.9800 ;
        RECT 1875.9000 2201.3000 1877.5000 2201.7800 ;
        RECT 1875.9000 2206.7400 1877.5000 2207.2200 ;
        RECT 1875.9000 2195.8600 1877.5000 2196.3400 ;
        RECT 1875.9000 2190.4200 1877.5000 2190.9000 ;
        RECT 1875.9000 2212.1800 1877.5000 2212.6600 ;
        RECT 1936.4400 2174.1000 1938.0400 2174.5800 ;
        RECT 1936.4400 2179.5400 1938.0400 2180.0200 ;
        RECT 1920.9000 2174.1000 1922.5000 2174.5800 ;
        RECT 1920.9000 2179.5400 1922.5000 2180.0200 ;
        RECT 1936.4400 2157.7800 1938.0400 2158.2600 ;
        RECT 1936.4400 2163.2200 1938.0400 2163.7000 ;
        RECT 1936.4400 2168.6600 1938.0400 2169.1400 ;
        RECT 1920.9000 2157.7800 1922.5000 2158.2600 ;
        RECT 1920.9000 2163.2200 1922.5000 2163.7000 ;
        RECT 1920.9000 2168.6600 1922.5000 2169.1400 ;
        RECT 1936.4400 2146.9000 1938.0400 2147.3800 ;
        RECT 1936.4400 2152.3400 1938.0400 2152.8200 ;
        RECT 1920.9000 2146.9000 1922.5000 2147.3800 ;
        RECT 1920.9000 2152.3400 1922.5000 2152.8200 ;
        RECT 1936.4400 2130.5800 1938.0400 2131.0600 ;
        RECT 1936.4400 2136.0200 1938.0400 2136.5000 ;
        RECT 1936.4400 2141.4600 1938.0400 2141.9400 ;
        RECT 1920.9000 2130.5800 1922.5000 2131.0600 ;
        RECT 1920.9000 2136.0200 1922.5000 2136.5000 ;
        RECT 1920.9000 2141.4600 1922.5000 2141.9400 ;
        RECT 1875.9000 2174.1000 1877.5000 2174.5800 ;
        RECT 1875.9000 2179.5400 1877.5000 2180.0200 ;
        RECT 1875.9000 2157.7800 1877.5000 2158.2600 ;
        RECT 1875.9000 2163.2200 1877.5000 2163.7000 ;
        RECT 1875.9000 2168.6600 1877.5000 2169.1400 ;
        RECT 1875.9000 2146.9000 1877.5000 2147.3800 ;
        RECT 1875.9000 2152.3400 1877.5000 2152.8200 ;
        RECT 1875.9000 2130.5800 1877.5000 2131.0600 ;
        RECT 1875.9000 2136.0200 1877.5000 2136.5000 ;
        RECT 1875.9000 2141.4600 1877.5000 2141.9400 ;
        RECT 1875.9000 2184.9800 1877.5000 2185.4600 ;
        RECT 1920.9000 2184.9800 1922.5000 2185.4600 ;
        RECT 1936.4400 2184.9800 1938.0400 2185.4600 ;
        RECT 1830.9000 2217.6200 1832.5000 2218.1000 ;
        RECT 1830.9000 2223.0600 1832.5000 2223.5400 ;
        RECT 1830.9000 2228.5000 1832.5000 2228.9800 ;
        RECT 1785.9000 2217.6200 1787.5000 2218.1000 ;
        RECT 1785.9000 2223.0600 1787.5000 2223.5400 ;
        RECT 1785.9000 2228.5000 1787.5000 2228.9800 ;
        RECT 1830.9000 2201.3000 1832.5000 2201.7800 ;
        RECT 1830.9000 2206.7400 1832.5000 2207.2200 ;
        RECT 1830.9000 2190.4200 1832.5000 2190.9000 ;
        RECT 1830.9000 2195.8600 1832.5000 2196.3400 ;
        RECT 1785.9000 2201.3000 1787.5000 2201.7800 ;
        RECT 1785.9000 2206.7400 1787.5000 2207.2200 ;
        RECT 1785.9000 2190.4200 1787.5000 2190.9000 ;
        RECT 1785.9000 2195.8600 1787.5000 2196.3400 ;
        RECT 1785.9000 2212.1800 1787.5000 2212.6600 ;
        RECT 1830.9000 2212.1800 1832.5000 2212.6600 ;
        RECT 1733.7400 2228.5000 1735.3400 2228.9800 ;
        RECT 1740.9000 2228.5000 1742.5000 2228.9800 ;
        RECT 1740.9000 2217.6200 1742.5000 2218.1000 ;
        RECT 1740.9000 2223.0600 1742.5000 2223.5400 ;
        RECT 1733.7400 2217.6200 1735.3400 2218.1000 ;
        RECT 1733.7400 2223.0600 1735.3400 2223.5400 ;
        RECT 1740.9000 2201.3000 1742.5000 2201.7800 ;
        RECT 1740.9000 2206.7400 1742.5000 2207.2200 ;
        RECT 1733.7400 2201.3000 1735.3400 2201.7800 ;
        RECT 1733.7400 2206.7400 1735.3400 2207.2200 ;
        RECT 1740.9000 2190.4200 1742.5000 2190.9000 ;
        RECT 1740.9000 2195.8600 1742.5000 2196.3400 ;
        RECT 1733.7400 2190.4200 1735.3400 2190.9000 ;
        RECT 1733.7400 2195.8600 1735.3400 2196.3400 ;
        RECT 1733.7400 2212.1800 1735.3400 2212.6600 ;
        RECT 1740.9000 2212.1800 1742.5000 2212.6600 ;
        RECT 1830.9000 2174.1000 1832.5000 2174.5800 ;
        RECT 1830.9000 2179.5400 1832.5000 2180.0200 ;
        RECT 1830.9000 2157.7800 1832.5000 2158.2600 ;
        RECT 1830.9000 2163.2200 1832.5000 2163.7000 ;
        RECT 1830.9000 2168.6600 1832.5000 2169.1400 ;
        RECT 1785.9000 2174.1000 1787.5000 2174.5800 ;
        RECT 1785.9000 2179.5400 1787.5000 2180.0200 ;
        RECT 1785.9000 2157.7800 1787.5000 2158.2600 ;
        RECT 1785.9000 2163.2200 1787.5000 2163.7000 ;
        RECT 1785.9000 2168.6600 1787.5000 2169.1400 ;
        RECT 1830.9000 2146.9000 1832.5000 2147.3800 ;
        RECT 1830.9000 2152.3400 1832.5000 2152.8200 ;
        RECT 1830.9000 2130.5800 1832.5000 2131.0600 ;
        RECT 1830.9000 2136.0200 1832.5000 2136.5000 ;
        RECT 1830.9000 2141.4600 1832.5000 2141.9400 ;
        RECT 1785.9000 2146.9000 1787.5000 2147.3800 ;
        RECT 1785.9000 2152.3400 1787.5000 2152.8200 ;
        RECT 1785.9000 2130.5800 1787.5000 2131.0600 ;
        RECT 1785.9000 2136.0200 1787.5000 2136.5000 ;
        RECT 1785.9000 2141.4600 1787.5000 2141.9400 ;
        RECT 1740.9000 2174.1000 1742.5000 2174.5800 ;
        RECT 1740.9000 2179.5400 1742.5000 2180.0200 ;
        RECT 1733.7400 2174.1000 1735.3400 2174.5800 ;
        RECT 1733.7400 2179.5400 1735.3400 2180.0200 ;
        RECT 1740.9000 2157.7800 1742.5000 2158.2600 ;
        RECT 1740.9000 2163.2200 1742.5000 2163.7000 ;
        RECT 1740.9000 2168.6600 1742.5000 2169.1400 ;
        RECT 1733.7400 2157.7800 1735.3400 2158.2600 ;
        RECT 1733.7400 2163.2200 1735.3400 2163.7000 ;
        RECT 1733.7400 2168.6600 1735.3400 2169.1400 ;
        RECT 1740.9000 2146.9000 1742.5000 2147.3800 ;
        RECT 1740.9000 2152.3400 1742.5000 2152.8200 ;
        RECT 1733.7400 2146.9000 1735.3400 2147.3800 ;
        RECT 1733.7400 2152.3400 1735.3400 2152.8200 ;
        RECT 1740.9000 2130.5800 1742.5000 2131.0600 ;
        RECT 1740.9000 2136.0200 1742.5000 2136.5000 ;
        RECT 1740.9000 2141.4600 1742.5000 2141.9400 ;
        RECT 1733.7400 2130.5800 1735.3400 2131.0600 ;
        RECT 1733.7400 2136.0200 1735.3400 2136.5000 ;
        RECT 1733.7400 2141.4600 1735.3400 2141.9400 ;
        RECT 1733.7400 2184.9800 1735.3400 2185.4600 ;
        RECT 1740.9000 2184.9800 1742.5000 2185.4600 ;
        RECT 1785.9000 2184.9800 1787.5000 2185.4600 ;
        RECT 1830.9000 2184.9800 1832.5000 2185.4600 ;
        RECT 1936.4400 2119.7000 1938.0400 2120.1800 ;
        RECT 1936.4400 2125.1400 1938.0400 2125.6200 ;
        RECT 1920.9000 2119.7000 1922.5000 2120.1800 ;
        RECT 1920.9000 2125.1400 1922.5000 2125.6200 ;
        RECT 1936.4400 2103.3800 1938.0400 2103.8600 ;
        RECT 1936.4400 2108.8200 1938.0400 2109.3000 ;
        RECT 1936.4400 2114.2600 1938.0400 2114.7400 ;
        RECT 1920.9000 2103.3800 1922.5000 2103.8600 ;
        RECT 1920.9000 2108.8200 1922.5000 2109.3000 ;
        RECT 1920.9000 2114.2600 1922.5000 2114.7400 ;
        RECT 1936.4400 2092.5000 1938.0400 2092.9800 ;
        RECT 1936.4400 2097.9400 1938.0400 2098.4200 ;
        RECT 1920.9000 2092.5000 1922.5000 2092.9800 ;
        RECT 1920.9000 2097.9400 1922.5000 2098.4200 ;
        RECT 1936.4400 2076.1800 1938.0400 2076.6600 ;
        RECT 1936.4400 2081.6200 1938.0400 2082.1000 ;
        RECT 1936.4400 2087.0600 1938.0400 2087.5400 ;
        RECT 1920.9000 2076.1800 1922.5000 2076.6600 ;
        RECT 1920.9000 2081.6200 1922.5000 2082.1000 ;
        RECT 1920.9000 2087.0600 1922.5000 2087.5400 ;
        RECT 1875.9000 2119.7000 1877.5000 2120.1800 ;
        RECT 1875.9000 2125.1400 1877.5000 2125.6200 ;
        RECT 1875.9000 2103.3800 1877.5000 2103.8600 ;
        RECT 1875.9000 2108.8200 1877.5000 2109.3000 ;
        RECT 1875.9000 2114.2600 1877.5000 2114.7400 ;
        RECT 1875.9000 2092.5000 1877.5000 2092.9800 ;
        RECT 1875.9000 2097.9400 1877.5000 2098.4200 ;
        RECT 1875.9000 2076.1800 1877.5000 2076.6600 ;
        RECT 1875.9000 2081.6200 1877.5000 2082.1000 ;
        RECT 1875.9000 2087.0600 1877.5000 2087.5400 ;
        RECT 1936.4400 2065.3000 1938.0400 2065.7800 ;
        RECT 1936.4400 2070.7400 1938.0400 2071.2200 ;
        RECT 1920.9000 2065.3000 1922.5000 2065.7800 ;
        RECT 1920.9000 2070.7400 1922.5000 2071.2200 ;
        RECT 1936.4400 2048.9800 1938.0400 2049.4600 ;
        RECT 1936.4400 2054.4200 1938.0400 2054.9000 ;
        RECT 1936.4400 2059.8600 1938.0400 2060.3400 ;
        RECT 1920.9000 2048.9800 1922.5000 2049.4600 ;
        RECT 1920.9000 2054.4200 1922.5000 2054.9000 ;
        RECT 1920.9000 2059.8600 1922.5000 2060.3400 ;
        RECT 1936.4400 2038.1000 1938.0400 2038.5800 ;
        RECT 1936.4400 2043.5400 1938.0400 2044.0200 ;
        RECT 1920.9000 2038.1000 1922.5000 2038.5800 ;
        RECT 1920.9000 2043.5400 1922.5000 2044.0200 ;
        RECT 1920.9000 2032.6600 1922.5000 2033.1400 ;
        RECT 1936.4400 2032.6600 1938.0400 2033.1400 ;
        RECT 1875.9000 2065.3000 1877.5000 2065.7800 ;
        RECT 1875.9000 2070.7400 1877.5000 2071.2200 ;
        RECT 1875.9000 2048.9800 1877.5000 2049.4600 ;
        RECT 1875.9000 2054.4200 1877.5000 2054.9000 ;
        RECT 1875.9000 2059.8600 1877.5000 2060.3400 ;
        RECT 1875.9000 2038.1000 1877.5000 2038.5800 ;
        RECT 1875.9000 2043.5400 1877.5000 2044.0200 ;
        RECT 1875.9000 2032.6600 1877.5000 2033.1400 ;
        RECT 1830.9000 2119.7000 1832.5000 2120.1800 ;
        RECT 1830.9000 2125.1400 1832.5000 2125.6200 ;
        RECT 1830.9000 2103.3800 1832.5000 2103.8600 ;
        RECT 1830.9000 2108.8200 1832.5000 2109.3000 ;
        RECT 1830.9000 2114.2600 1832.5000 2114.7400 ;
        RECT 1785.9000 2119.7000 1787.5000 2120.1800 ;
        RECT 1785.9000 2125.1400 1787.5000 2125.6200 ;
        RECT 1785.9000 2103.3800 1787.5000 2103.8600 ;
        RECT 1785.9000 2108.8200 1787.5000 2109.3000 ;
        RECT 1785.9000 2114.2600 1787.5000 2114.7400 ;
        RECT 1830.9000 2092.5000 1832.5000 2092.9800 ;
        RECT 1830.9000 2097.9400 1832.5000 2098.4200 ;
        RECT 1830.9000 2076.1800 1832.5000 2076.6600 ;
        RECT 1830.9000 2081.6200 1832.5000 2082.1000 ;
        RECT 1830.9000 2087.0600 1832.5000 2087.5400 ;
        RECT 1785.9000 2092.5000 1787.5000 2092.9800 ;
        RECT 1785.9000 2097.9400 1787.5000 2098.4200 ;
        RECT 1785.9000 2076.1800 1787.5000 2076.6600 ;
        RECT 1785.9000 2081.6200 1787.5000 2082.1000 ;
        RECT 1785.9000 2087.0600 1787.5000 2087.5400 ;
        RECT 1740.9000 2119.7000 1742.5000 2120.1800 ;
        RECT 1740.9000 2125.1400 1742.5000 2125.6200 ;
        RECT 1733.7400 2119.7000 1735.3400 2120.1800 ;
        RECT 1733.7400 2125.1400 1735.3400 2125.6200 ;
        RECT 1740.9000 2103.3800 1742.5000 2103.8600 ;
        RECT 1740.9000 2108.8200 1742.5000 2109.3000 ;
        RECT 1740.9000 2114.2600 1742.5000 2114.7400 ;
        RECT 1733.7400 2103.3800 1735.3400 2103.8600 ;
        RECT 1733.7400 2108.8200 1735.3400 2109.3000 ;
        RECT 1733.7400 2114.2600 1735.3400 2114.7400 ;
        RECT 1740.9000 2092.5000 1742.5000 2092.9800 ;
        RECT 1740.9000 2097.9400 1742.5000 2098.4200 ;
        RECT 1733.7400 2092.5000 1735.3400 2092.9800 ;
        RECT 1733.7400 2097.9400 1735.3400 2098.4200 ;
        RECT 1740.9000 2076.1800 1742.5000 2076.6600 ;
        RECT 1740.9000 2081.6200 1742.5000 2082.1000 ;
        RECT 1740.9000 2087.0600 1742.5000 2087.5400 ;
        RECT 1733.7400 2076.1800 1735.3400 2076.6600 ;
        RECT 1733.7400 2081.6200 1735.3400 2082.1000 ;
        RECT 1733.7400 2087.0600 1735.3400 2087.5400 ;
        RECT 1830.9000 2065.3000 1832.5000 2065.7800 ;
        RECT 1830.9000 2070.7400 1832.5000 2071.2200 ;
        RECT 1830.9000 2048.9800 1832.5000 2049.4600 ;
        RECT 1830.9000 2054.4200 1832.5000 2054.9000 ;
        RECT 1830.9000 2059.8600 1832.5000 2060.3400 ;
        RECT 1785.9000 2065.3000 1787.5000 2065.7800 ;
        RECT 1785.9000 2070.7400 1787.5000 2071.2200 ;
        RECT 1785.9000 2048.9800 1787.5000 2049.4600 ;
        RECT 1785.9000 2054.4200 1787.5000 2054.9000 ;
        RECT 1785.9000 2059.8600 1787.5000 2060.3400 ;
        RECT 1830.9000 2043.5400 1832.5000 2044.0200 ;
        RECT 1830.9000 2038.1000 1832.5000 2038.5800 ;
        RECT 1830.9000 2032.6600 1832.5000 2033.1400 ;
        RECT 1785.9000 2043.5400 1787.5000 2044.0200 ;
        RECT 1785.9000 2038.1000 1787.5000 2038.5800 ;
        RECT 1785.9000 2032.6600 1787.5000 2033.1400 ;
        RECT 1740.9000 2065.3000 1742.5000 2065.7800 ;
        RECT 1740.9000 2070.7400 1742.5000 2071.2200 ;
        RECT 1733.7400 2065.3000 1735.3400 2065.7800 ;
        RECT 1733.7400 2070.7400 1735.3400 2071.2200 ;
        RECT 1740.9000 2048.9800 1742.5000 2049.4600 ;
        RECT 1740.9000 2054.4200 1742.5000 2054.9000 ;
        RECT 1740.9000 2059.8600 1742.5000 2060.3400 ;
        RECT 1733.7400 2048.9800 1735.3400 2049.4600 ;
        RECT 1733.7400 2054.4200 1735.3400 2054.9000 ;
        RECT 1733.7400 2059.8600 1735.3400 2060.3400 ;
        RECT 1740.9000 2038.1000 1742.5000 2038.5800 ;
        RECT 1740.9000 2043.5400 1742.5000 2044.0200 ;
        RECT 1733.7400 2038.1000 1735.3400 2038.5800 ;
        RECT 1733.7400 2043.5400 1735.3400 2044.0200 ;
        RECT 1733.7400 2032.6600 1735.3400 2033.1400 ;
        RECT 1740.9000 2032.6600 1742.5000 2033.1400 ;
        RECT 1730.7800 2234.8500 1941.0000 2236.4500 ;
        RECT 1730.7800 2023.1500 1941.0000 2024.7500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 2020.3200 1735.3400 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 2238.3600 1735.3400 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 2020.3200 1938.0400 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 2238.3600 1938.0400 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2023.1500 1732.3800 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2023.1500 1941.0000 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2234.8500 1732.3800 2236.4500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2234.8500 1941.0000 2236.4500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 1793.5100 1922.5000 2006.8100 ;
        RECT 1875.9000 1793.5100 1877.5000 2006.8100 ;
        RECT 1830.9000 1793.5100 1832.5000 2006.8100 ;
        RECT 1785.9000 1793.5100 1787.5000 2006.8100 ;
        RECT 1740.9000 1793.5100 1742.5000 2006.8100 ;
        RECT 1936.4400 1790.6800 1938.0400 2010.3200 ;
        RECT 1733.7400 1790.6800 1735.3400 2010.3200 ;
      LAYER met3 ;
        RECT 1920.9000 1998.8600 1922.5000 1999.3400 ;
        RECT 1936.4400 1998.8600 1938.0400 1999.3400 ;
        RECT 1936.4400 1987.9800 1938.0400 1988.4600 ;
        RECT 1936.4400 1993.4200 1938.0400 1993.9000 ;
        RECT 1920.9000 1987.9800 1922.5000 1988.4600 ;
        RECT 1920.9000 1993.4200 1922.5000 1993.9000 ;
        RECT 1936.4400 1971.6600 1938.0400 1972.1400 ;
        RECT 1936.4400 1977.1000 1938.0400 1977.5800 ;
        RECT 1920.9000 1971.6600 1922.5000 1972.1400 ;
        RECT 1920.9000 1977.1000 1922.5000 1977.5800 ;
        RECT 1936.4400 1960.7800 1938.0400 1961.2600 ;
        RECT 1936.4400 1966.2200 1938.0400 1966.7000 ;
        RECT 1920.9000 1960.7800 1922.5000 1961.2600 ;
        RECT 1920.9000 1966.2200 1922.5000 1966.7000 ;
        RECT 1920.9000 1982.5400 1922.5000 1983.0200 ;
        RECT 1936.4400 1982.5400 1938.0400 1983.0200 ;
        RECT 1875.9000 1987.9800 1877.5000 1988.4600 ;
        RECT 1875.9000 1993.4200 1877.5000 1993.9000 ;
        RECT 1875.9000 1998.8600 1877.5000 1999.3400 ;
        RECT 1875.9000 1971.6600 1877.5000 1972.1400 ;
        RECT 1875.9000 1977.1000 1877.5000 1977.5800 ;
        RECT 1875.9000 1966.2200 1877.5000 1966.7000 ;
        RECT 1875.9000 1960.7800 1877.5000 1961.2600 ;
        RECT 1875.9000 1982.5400 1877.5000 1983.0200 ;
        RECT 1936.4400 1944.4600 1938.0400 1944.9400 ;
        RECT 1936.4400 1949.9000 1938.0400 1950.3800 ;
        RECT 1920.9000 1944.4600 1922.5000 1944.9400 ;
        RECT 1920.9000 1949.9000 1922.5000 1950.3800 ;
        RECT 1936.4400 1928.1400 1938.0400 1928.6200 ;
        RECT 1936.4400 1933.5800 1938.0400 1934.0600 ;
        RECT 1936.4400 1939.0200 1938.0400 1939.5000 ;
        RECT 1920.9000 1928.1400 1922.5000 1928.6200 ;
        RECT 1920.9000 1933.5800 1922.5000 1934.0600 ;
        RECT 1920.9000 1939.0200 1922.5000 1939.5000 ;
        RECT 1936.4400 1917.2600 1938.0400 1917.7400 ;
        RECT 1936.4400 1922.7000 1938.0400 1923.1800 ;
        RECT 1920.9000 1917.2600 1922.5000 1917.7400 ;
        RECT 1920.9000 1922.7000 1922.5000 1923.1800 ;
        RECT 1936.4400 1900.9400 1938.0400 1901.4200 ;
        RECT 1936.4400 1906.3800 1938.0400 1906.8600 ;
        RECT 1936.4400 1911.8200 1938.0400 1912.3000 ;
        RECT 1920.9000 1900.9400 1922.5000 1901.4200 ;
        RECT 1920.9000 1906.3800 1922.5000 1906.8600 ;
        RECT 1920.9000 1911.8200 1922.5000 1912.3000 ;
        RECT 1875.9000 1944.4600 1877.5000 1944.9400 ;
        RECT 1875.9000 1949.9000 1877.5000 1950.3800 ;
        RECT 1875.9000 1928.1400 1877.5000 1928.6200 ;
        RECT 1875.9000 1933.5800 1877.5000 1934.0600 ;
        RECT 1875.9000 1939.0200 1877.5000 1939.5000 ;
        RECT 1875.9000 1917.2600 1877.5000 1917.7400 ;
        RECT 1875.9000 1922.7000 1877.5000 1923.1800 ;
        RECT 1875.9000 1900.9400 1877.5000 1901.4200 ;
        RECT 1875.9000 1906.3800 1877.5000 1906.8600 ;
        RECT 1875.9000 1911.8200 1877.5000 1912.3000 ;
        RECT 1875.9000 1955.3400 1877.5000 1955.8200 ;
        RECT 1920.9000 1955.3400 1922.5000 1955.8200 ;
        RECT 1936.4400 1955.3400 1938.0400 1955.8200 ;
        RECT 1830.9000 1987.9800 1832.5000 1988.4600 ;
        RECT 1830.9000 1993.4200 1832.5000 1993.9000 ;
        RECT 1830.9000 1998.8600 1832.5000 1999.3400 ;
        RECT 1785.9000 1987.9800 1787.5000 1988.4600 ;
        RECT 1785.9000 1993.4200 1787.5000 1993.9000 ;
        RECT 1785.9000 1998.8600 1787.5000 1999.3400 ;
        RECT 1830.9000 1971.6600 1832.5000 1972.1400 ;
        RECT 1830.9000 1977.1000 1832.5000 1977.5800 ;
        RECT 1830.9000 1960.7800 1832.5000 1961.2600 ;
        RECT 1830.9000 1966.2200 1832.5000 1966.7000 ;
        RECT 1785.9000 1971.6600 1787.5000 1972.1400 ;
        RECT 1785.9000 1977.1000 1787.5000 1977.5800 ;
        RECT 1785.9000 1960.7800 1787.5000 1961.2600 ;
        RECT 1785.9000 1966.2200 1787.5000 1966.7000 ;
        RECT 1785.9000 1982.5400 1787.5000 1983.0200 ;
        RECT 1830.9000 1982.5400 1832.5000 1983.0200 ;
        RECT 1733.7400 1998.8600 1735.3400 1999.3400 ;
        RECT 1740.9000 1998.8600 1742.5000 1999.3400 ;
        RECT 1740.9000 1987.9800 1742.5000 1988.4600 ;
        RECT 1740.9000 1993.4200 1742.5000 1993.9000 ;
        RECT 1733.7400 1987.9800 1735.3400 1988.4600 ;
        RECT 1733.7400 1993.4200 1735.3400 1993.9000 ;
        RECT 1740.9000 1971.6600 1742.5000 1972.1400 ;
        RECT 1740.9000 1977.1000 1742.5000 1977.5800 ;
        RECT 1733.7400 1971.6600 1735.3400 1972.1400 ;
        RECT 1733.7400 1977.1000 1735.3400 1977.5800 ;
        RECT 1740.9000 1960.7800 1742.5000 1961.2600 ;
        RECT 1740.9000 1966.2200 1742.5000 1966.7000 ;
        RECT 1733.7400 1960.7800 1735.3400 1961.2600 ;
        RECT 1733.7400 1966.2200 1735.3400 1966.7000 ;
        RECT 1733.7400 1982.5400 1735.3400 1983.0200 ;
        RECT 1740.9000 1982.5400 1742.5000 1983.0200 ;
        RECT 1830.9000 1944.4600 1832.5000 1944.9400 ;
        RECT 1830.9000 1949.9000 1832.5000 1950.3800 ;
        RECT 1830.9000 1928.1400 1832.5000 1928.6200 ;
        RECT 1830.9000 1933.5800 1832.5000 1934.0600 ;
        RECT 1830.9000 1939.0200 1832.5000 1939.5000 ;
        RECT 1785.9000 1944.4600 1787.5000 1944.9400 ;
        RECT 1785.9000 1949.9000 1787.5000 1950.3800 ;
        RECT 1785.9000 1928.1400 1787.5000 1928.6200 ;
        RECT 1785.9000 1933.5800 1787.5000 1934.0600 ;
        RECT 1785.9000 1939.0200 1787.5000 1939.5000 ;
        RECT 1830.9000 1917.2600 1832.5000 1917.7400 ;
        RECT 1830.9000 1922.7000 1832.5000 1923.1800 ;
        RECT 1830.9000 1900.9400 1832.5000 1901.4200 ;
        RECT 1830.9000 1906.3800 1832.5000 1906.8600 ;
        RECT 1830.9000 1911.8200 1832.5000 1912.3000 ;
        RECT 1785.9000 1917.2600 1787.5000 1917.7400 ;
        RECT 1785.9000 1922.7000 1787.5000 1923.1800 ;
        RECT 1785.9000 1900.9400 1787.5000 1901.4200 ;
        RECT 1785.9000 1906.3800 1787.5000 1906.8600 ;
        RECT 1785.9000 1911.8200 1787.5000 1912.3000 ;
        RECT 1740.9000 1944.4600 1742.5000 1944.9400 ;
        RECT 1740.9000 1949.9000 1742.5000 1950.3800 ;
        RECT 1733.7400 1944.4600 1735.3400 1944.9400 ;
        RECT 1733.7400 1949.9000 1735.3400 1950.3800 ;
        RECT 1740.9000 1928.1400 1742.5000 1928.6200 ;
        RECT 1740.9000 1933.5800 1742.5000 1934.0600 ;
        RECT 1740.9000 1939.0200 1742.5000 1939.5000 ;
        RECT 1733.7400 1928.1400 1735.3400 1928.6200 ;
        RECT 1733.7400 1933.5800 1735.3400 1934.0600 ;
        RECT 1733.7400 1939.0200 1735.3400 1939.5000 ;
        RECT 1740.9000 1917.2600 1742.5000 1917.7400 ;
        RECT 1740.9000 1922.7000 1742.5000 1923.1800 ;
        RECT 1733.7400 1917.2600 1735.3400 1917.7400 ;
        RECT 1733.7400 1922.7000 1735.3400 1923.1800 ;
        RECT 1740.9000 1900.9400 1742.5000 1901.4200 ;
        RECT 1740.9000 1906.3800 1742.5000 1906.8600 ;
        RECT 1740.9000 1911.8200 1742.5000 1912.3000 ;
        RECT 1733.7400 1900.9400 1735.3400 1901.4200 ;
        RECT 1733.7400 1906.3800 1735.3400 1906.8600 ;
        RECT 1733.7400 1911.8200 1735.3400 1912.3000 ;
        RECT 1733.7400 1955.3400 1735.3400 1955.8200 ;
        RECT 1740.9000 1955.3400 1742.5000 1955.8200 ;
        RECT 1785.9000 1955.3400 1787.5000 1955.8200 ;
        RECT 1830.9000 1955.3400 1832.5000 1955.8200 ;
        RECT 1936.4400 1890.0600 1938.0400 1890.5400 ;
        RECT 1936.4400 1895.5000 1938.0400 1895.9800 ;
        RECT 1920.9000 1890.0600 1922.5000 1890.5400 ;
        RECT 1920.9000 1895.5000 1922.5000 1895.9800 ;
        RECT 1936.4400 1873.7400 1938.0400 1874.2200 ;
        RECT 1936.4400 1879.1800 1938.0400 1879.6600 ;
        RECT 1936.4400 1884.6200 1938.0400 1885.1000 ;
        RECT 1920.9000 1873.7400 1922.5000 1874.2200 ;
        RECT 1920.9000 1879.1800 1922.5000 1879.6600 ;
        RECT 1920.9000 1884.6200 1922.5000 1885.1000 ;
        RECT 1936.4400 1862.8600 1938.0400 1863.3400 ;
        RECT 1936.4400 1868.3000 1938.0400 1868.7800 ;
        RECT 1920.9000 1862.8600 1922.5000 1863.3400 ;
        RECT 1920.9000 1868.3000 1922.5000 1868.7800 ;
        RECT 1936.4400 1846.5400 1938.0400 1847.0200 ;
        RECT 1936.4400 1851.9800 1938.0400 1852.4600 ;
        RECT 1936.4400 1857.4200 1938.0400 1857.9000 ;
        RECT 1920.9000 1846.5400 1922.5000 1847.0200 ;
        RECT 1920.9000 1851.9800 1922.5000 1852.4600 ;
        RECT 1920.9000 1857.4200 1922.5000 1857.9000 ;
        RECT 1875.9000 1890.0600 1877.5000 1890.5400 ;
        RECT 1875.9000 1895.5000 1877.5000 1895.9800 ;
        RECT 1875.9000 1873.7400 1877.5000 1874.2200 ;
        RECT 1875.9000 1879.1800 1877.5000 1879.6600 ;
        RECT 1875.9000 1884.6200 1877.5000 1885.1000 ;
        RECT 1875.9000 1862.8600 1877.5000 1863.3400 ;
        RECT 1875.9000 1868.3000 1877.5000 1868.7800 ;
        RECT 1875.9000 1846.5400 1877.5000 1847.0200 ;
        RECT 1875.9000 1851.9800 1877.5000 1852.4600 ;
        RECT 1875.9000 1857.4200 1877.5000 1857.9000 ;
        RECT 1936.4400 1835.6600 1938.0400 1836.1400 ;
        RECT 1936.4400 1841.1000 1938.0400 1841.5800 ;
        RECT 1920.9000 1835.6600 1922.5000 1836.1400 ;
        RECT 1920.9000 1841.1000 1922.5000 1841.5800 ;
        RECT 1936.4400 1819.3400 1938.0400 1819.8200 ;
        RECT 1936.4400 1824.7800 1938.0400 1825.2600 ;
        RECT 1936.4400 1830.2200 1938.0400 1830.7000 ;
        RECT 1920.9000 1819.3400 1922.5000 1819.8200 ;
        RECT 1920.9000 1824.7800 1922.5000 1825.2600 ;
        RECT 1920.9000 1830.2200 1922.5000 1830.7000 ;
        RECT 1936.4400 1808.4600 1938.0400 1808.9400 ;
        RECT 1936.4400 1813.9000 1938.0400 1814.3800 ;
        RECT 1920.9000 1808.4600 1922.5000 1808.9400 ;
        RECT 1920.9000 1813.9000 1922.5000 1814.3800 ;
        RECT 1920.9000 1803.0200 1922.5000 1803.5000 ;
        RECT 1936.4400 1803.0200 1938.0400 1803.5000 ;
        RECT 1875.9000 1835.6600 1877.5000 1836.1400 ;
        RECT 1875.9000 1841.1000 1877.5000 1841.5800 ;
        RECT 1875.9000 1819.3400 1877.5000 1819.8200 ;
        RECT 1875.9000 1824.7800 1877.5000 1825.2600 ;
        RECT 1875.9000 1830.2200 1877.5000 1830.7000 ;
        RECT 1875.9000 1808.4600 1877.5000 1808.9400 ;
        RECT 1875.9000 1813.9000 1877.5000 1814.3800 ;
        RECT 1875.9000 1803.0200 1877.5000 1803.5000 ;
        RECT 1830.9000 1890.0600 1832.5000 1890.5400 ;
        RECT 1830.9000 1895.5000 1832.5000 1895.9800 ;
        RECT 1830.9000 1873.7400 1832.5000 1874.2200 ;
        RECT 1830.9000 1879.1800 1832.5000 1879.6600 ;
        RECT 1830.9000 1884.6200 1832.5000 1885.1000 ;
        RECT 1785.9000 1890.0600 1787.5000 1890.5400 ;
        RECT 1785.9000 1895.5000 1787.5000 1895.9800 ;
        RECT 1785.9000 1873.7400 1787.5000 1874.2200 ;
        RECT 1785.9000 1879.1800 1787.5000 1879.6600 ;
        RECT 1785.9000 1884.6200 1787.5000 1885.1000 ;
        RECT 1830.9000 1862.8600 1832.5000 1863.3400 ;
        RECT 1830.9000 1868.3000 1832.5000 1868.7800 ;
        RECT 1830.9000 1846.5400 1832.5000 1847.0200 ;
        RECT 1830.9000 1851.9800 1832.5000 1852.4600 ;
        RECT 1830.9000 1857.4200 1832.5000 1857.9000 ;
        RECT 1785.9000 1862.8600 1787.5000 1863.3400 ;
        RECT 1785.9000 1868.3000 1787.5000 1868.7800 ;
        RECT 1785.9000 1846.5400 1787.5000 1847.0200 ;
        RECT 1785.9000 1851.9800 1787.5000 1852.4600 ;
        RECT 1785.9000 1857.4200 1787.5000 1857.9000 ;
        RECT 1740.9000 1890.0600 1742.5000 1890.5400 ;
        RECT 1740.9000 1895.5000 1742.5000 1895.9800 ;
        RECT 1733.7400 1890.0600 1735.3400 1890.5400 ;
        RECT 1733.7400 1895.5000 1735.3400 1895.9800 ;
        RECT 1740.9000 1873.7400 1742.5000 1874.2200 ;
        RECT 1740.9000 1879.1800 1742.5000 1879.6600 ;
        RECT 1740.9000 1884.6200 1742.5000 1885.1000 ;
        RECT 1733.7400 1873.7400 1735.3400 1874.2200 ;
        RECT 1733.7400 1879.1800 1735.3400 1879.6600 ;
        RECT 1733.7400 1884.6200 1735.3400 1885.1000 ;
        RECT 1740.9000 1862.8600 1742.5000 1863.3400 ;
        RECT 1740.9000 1868.3000 1742.5000 1868.7800 ;
        RECT 1733.7400 1862.8600 1735.3400 1863.3400 ;
        RECT 1733.7400 1868.3000 1735.3400 1868.7800 ;
        RECT 1740.9000 1846.5400 1742.5000 1847.0200 ;
        RECT 1740.9000 1851.9800 1742.5000 1852.4600 ;
        RECT 1740.9000 1857.4200 1742.5000 1857.9000 ;
        RECT 1733.7400 1846.5400 1735.3400 1847.0200 ;
        RECT 1733.7400 1851.9800 1735.3400 1852.4600 ;
        RECT 1733.7400 1857.4200 1735.3400 1857.9000 ;
        RECT 1830.9000 1835.6600 1832.5000 1836.1400 ;
        RECT 1830.9000 1841.1000 1832.5000 1841.5800 ;
        RECT 1830.9000 1819.3400 1832.5000 1819.8200 ;
        RECT 1830.9000 1824.7800 1832.5000 1825.2600 ;
        RECT 1830.9000 1830.2200 1832.5000 1830.7000 ;
        RECT 1785.9000 1835.6600 1787.5000 1836.1400 ;
        RECT 1785.9000 1841.1000 1787.5000 1841.5800 ;
        RECT 1785.9000 1819.3400 1787.5000 1819.8200 ;
        RECT 1785.9000 1824.7800 1787.5000 1825.2600 ;
        RECT 1785.9000 1830.2200 1787.5000 1830.7000 ;
        RECT 1830.9000 1813.9000 1832.5000 1814.3800 ;
        RECT 1830.9000 1808.4600 1832.5000 1808.9400 ;
        RECT 1830.9000 1803.0200 1832.5000 1803.5000 ;
        RECT 1785.9000 1813.9000 1787.5000 1814.3800 ;
        RECT 1785.9000 1808.4600 1787.5000 1808.9400 ;
        RECT 1785.9000 1803.0200 1787.5000 1803.5000 ;
        RECT 1740.9000 1835.6600 1742.5000 1836.1400 ;
        RECT 1740.9000 1841.1000 1742.5000 1841.5800 ;
        RECT 1733.7400 1835.6600 1735.3400 1836.1400 ;
        RECT 1733.7400 1841.1000 1735.3400 1841.5800 ;
        RECT 1740.9000 1819.3400 1742.5000 1819.8200 ;
        RECT 1740.9000 1824.7800 1742.5000 1825.2600 ;
        RECT 1740.9000 1830.2200 1742.5000 1830.7000 ;
        RECT 1733.7400 1819.3400 1735.3400 1819.8200 ;
        RECT 1733.7400 1824.7800 1735.3400 1825.2600 ;
        RECT 1733.7400 1830.2200 1735.3400 1830.7000 ;
        RECT 1740.9000 1808.4600 1742.5000 1808.9400 ;
        RECT 1740.9000 1813.9000 1742.5000 1814.3800 ;
        RECT 1733.7400 1808.4600 1735.3400 1808.9400 ;
        RECT 1733.7400 1813.9000 1735.3400 1814.3800 ;
        RECT 1733.7400 1803.0200 1735.3400 1803.5000 ;
        RECT 1740.9000 1803.0200 1742.5000 1803.5000 ;
        RECT 1730.7800 2005.2100 1941.0000 2006.8100 ;
        RECT 1730.7800 1793.5100 1941.0000 1795.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1790.6800 1735.3400 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 2008.7200 1735.3400 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1790.6800 1938.0400 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 2008.7200 1938.0400 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1793.5100 1732.3800 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1793.5100 1941.0000 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2005.2100 1732.3800 2006.8100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2005.2100 1941.0000 2006.8100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 1563.8700 1922.5000 1777.1700 ;
        RECT 1875.9000 1563.8700 1877.5000 1777.1700 ;
        RECT 1830.9000 1563.8700 1832.5000 1777.1700 ;
        RECT 1785.9000 1563.8700 1787.5000 1777.1700 ;
        RECT 1740.9000 1563.8700 1742.5000 1777.1700 ;
        RECT 1936.4400 1561.0400 1938.0400 1780.6800 ;
        RECT 1733.7400 1561.0400 1735.3400 1780.6800 ;
      LAYER met3 ;
        RECT 1920.9000 1769.2200 1922.5000 1769.7000 ;
        RECT 1936.4400 1769.2200 1938.0400 1769.7000 ;
        RECT 1936.4400 1758.3400 1938.0400 1758.8200 ;
        RECT 1936.4400 1763.7800 1938.0400 1764.2600 ;
        RECT 1920.9000 1758.3400 1922.5000 1758.8200 ;
        RECT 1920.9000 1763.7800 1922.5000 1764.2600 ;
        RECT 1936.4400 1742.0200 1938.0400 1742.5000 ;
        RECT 1936.4400 1747.4600 1938.0400 1747.9400 ;
        RECT 1920.9000 1742.0200 1922.5000 1742.5000 ;
        RECT 1920.9000 1747.4600 1922.5000 1747.9400 ;
        RECT 1936.4400 1731.1400 1938.0400 1731.6200 ;
        RECT 1936.4400 1736.5800 1938.0400 1737.0600 ;
        RECT 1920.9000 1731.1400 1922.5000 1731.6200 ;
        RECT 1920.9000 1736.5800 1922.5000 1737.0600 ;
        RECT 1920.9000 1752.9000 1922.5000 1753.3800 ;
        RECT 1936.4400 1752.9000 1938.0400 1753.3800 ;
        RECT 1875.9000 1758.3400 1877.5000 1758.8200 ;
        RECT 1875.9000 1763.7800 1877.5000 1764.2600 ;
        RECT 1875.9000 1769.2200 1877.5000 1769.7000 ;
        RECT 1875.9000 1742.0200 1877.5000 1742.5000 ;
        RECT 1875.9000 1747.4600 1877.5000 1747.9400 ;
        RECT 1875.9000 1736.5800 1877.5000 1737.0600 ;
        RECT 1875.9000 1731.1400 1877.5000 1731.6200 ;
        RECT 1875.9000 1752.9000 1877.5000 1753.3800 ;
        RECT 1936.4400 1714.8200 1938.0400 1715.3000 ;
        RECT 1936.4400 1720.2600 1938.0400 1720.7400 ;
        RECT 1920.9000 1714.8200 1922.5000 1715.3000 ;
        RECT 1920.9000 1720.2600 1922.5000 1720.7400 ;
        RECT 1936.4400 1698.5000 1938.0400 1698.9800 ;
        RECT 1936.4400 1703.9400 1938.0400 1704.4200 ;
        RECT 1936.4400 1709.3800 1938.0400 1709.8600 ;
        RECT 1920.9000 1698.5000 1922.5000 1698.9800 ;
        RECT 1920.9000 1703.9400 1922.5000 1704.4200 ;
        RECT 1920.9000 1709.3800 1922.5000 1709.8600 ;
        RECT 1936.4400 1687.6200 1938.0400 1688.1000 ;
        RECT 1936.4400 1693.0600 1938.0400 1693.5400 ;
        RECT 1920.9000 1687.6200 1922.5000 1688.1000 ;
        RECT 1920.9000 1693.0600 1922.5000 1693.5400 ;
        RECT 1936.4400 1671.3000 1938.0400 1671.7800 ;
        RECT 1936.4400 1676.7400 1938.0400 1677.2200 ;
        RECT 1936.4400 1682.1800 1938.0400 1682.6600 ;
        RECT 1920.9000 1671.3000 1922.5000 1671.7800 ;
        RECT 1920.9000 1676.7400 1922.5000 1677.2200 ;
        RECT 1920.9000 1682.1800 1922.5000 1682.6600 ;
        RECT 1875.9000 1714.8200 1877.5000 1715.3000 ;
        RECT 1875.9000 1720.2600 1877.5000 1720.7400 ;
        RECT 1875.9000 1698.5000 1877.5000 1698.9800 ;
        RECT 1875.9000 1703.9400 1877.5000 1704.4200 ;
        RECT 1875.9000 1709.3800 1877.5000 1709.8600 ;
        RECT 1875.9000 1687.6200 1877.5000 1688.1000 ;
        RECT 1875.9000 1693.0600 1877.5000 1693.5400 ;
        RECT 1875.9000 1671.3000 1877.5000 1671.7800 ;
        RECT 1875.9000 1676.7400 1877.5000 1677.2200 ;
        RECT 1875.9000 1682.1800 1877.5000 1682.6600 ;
        RECT 1875.9000 1725.7000 1877.5000 1726.1800 ;
        RECT 1920.9000 1725.7000 1922.5000 1726.1800 ;
        RECT 1936.4400 1725.7000 1938.0400 1726.1800 ;
        RECT 1830.9000 1758.3400 1832.5000 1758.8200 ;
        RECT 1830.9000 1763.7800 1832.5000 1764.2600 ;
        RECT 1830.9000 1769.2200 1832.5000 1769.7000 ;
        RECT 1785.9000 1758.3400 1787.5000 1758.8200 ;
        RECT 1785.9000 1763.7800 1787.5000 1764.2600 ;
        RECT 1785.9000 1769.2200 1787.5000 1769.7000 ;
        RECT 1830.9000 1742.0200 1832.5000 1742.5000 ;
        RECT 1830.9000 1747.4600 1832.5000 1747.9400 ;
        RECT 1830.9000 1731.1400 1832.5000 1731.6200 ;
        RECT 1830.9000 1736.5800 1832.5000 1737.0600 ;
        RECT 1785.9000 1742.0200 1787.5000 1742.5000 ;
        RECT 1785.9000 1747.4600 1787.5000 1747.9400 ;
        RECT 1785.9000 1731.1400 1787.5000 1731.6200 ;
        RECT 1785.9000 1736.5800 1787.5000 1737.0600 ;
        RECT 1785.9000 1752.9000 1787.5000 1753.3800 ;
        RECT 1830.9000 1752.9000 1832.5000 1753.3800 ;
        RECT 1733.7400 1769.2200 1735.3400 1769.7000 ;
        RECT 1740.9000 1769.2200 1742.5000 1769.7000 ;
        RECT 1740.9000 1758.3400 1742.5000 1758.8200 ;
        RECT 1740.9000 1763.7800 1742.5000 1764.2600 ;
        RECT 1733.7400 1758.3400 1735.3400 1758.8200 ;
        RECT 1733.7400 1763.7800 1735.3400 1764.2600 ;
        RECT 1740.9000 1742.0200 1742.5000 1742.5000 ;
        RECT 1740.9000 1747.4600 1742.5000 1747.9400 ;
        RECT 1733.7400 1742.0200 1735.3400 1742.5000 ;
        RECT 1733.7400 1747.4600 1735.3400 1747.9400 ;
        RECT 1740.9000 1731.1400 1742.5000 1731.6200 ;
        RECT 1740.9000 1736.5800 1742.5000 1737.0600 ;
        RECT 1733.7400 1731.1400 1735.3400 1731.6200 ;
        RECT 1733.7400 1736.5800 1735.3400 1737.0600 ;
        RECT 1733.7400 1752.9000 1735.3400 1753.3800 ;
        RECT 1740.9000 1752.9000 1742.5000 1753.3800 ;
        RECT 1830.9000 1714.8200 1832.5000 1715.3000 ;
        RECT 1830.9000 1720.2600 1832.5000 1720.7400 ;
        RECT 1830.9000 1698.5000 1832.5000 1698.9800 ;
        RECT 1830.9000 1703.9400 1832.5000 1704.4200 ;
        RECT 1830.9000 1709.3800 1832.5000 1709.8600 ;
        RECT 1785.9000 1714.8200 1787.5000 1715.3000 ;
        RECT 1785.9000 1720.2600 1787.5000 1720.7400 ;
        RECT 1785.9000 1698.5000 1787.5000 1698.9800 ;
        RECT 1785.9000 1703.9400 1787.5000 1704.4200 ;
        RECT 1785.9000 1709.3800 1787.5000 1709.8600 ;
        RECT 1830.9000 1687.6200 1832.5000 1688.1000 ;
        RECT 1830.9000 1693.0600 1832.5000 1693.5400 ;
        RECT 1830.9000 1671.3000 1832.5000 1671.7800 ;
        RECT 1830.9000 1676.7400 1832.5000 1677.2200 ;
        RECT 1830.9000 1682.1800 1832.5000 1682.6600 ;
        RECT 1785.9000 1687.6200 1787.5000 1688.1000 ;
        RECT 1785.9000 1693.0600 1787.5000 1693.5400 ;
        RECT 1785.9000 1671.3000 1787.5000 1671.7800 ;
        RECT 1785.9000 1676.7400 1787.5000 1677.2200 ;
        RECT 1785.9000 1682.1800 1787.5000 1682.6600 ;
        RECT 1740.9000 1714.8200 1742.5000 1715.3000 ;
        RECT 1740.9000 1720.2600 1742.5000 1720.7400 ;
        RECT 1733.7400 1714.8200 1735.3400 1715.3000 ;
        RECT 1733.7400 1720.2600 1735.3400 1720.7400 ;
        RECT 1740.9000 1698.5000 1742.5000 1698.9800 ;
        RECT 1740.9000 1703.9400 1742.5000 1704.4200 ;
        RECT 1740.9000 1709.3800 1742.5000 1709.8600 ;
        RECT 1733.7400 1698.5000 1735.3400 1698.9800 ;
        RECT 1733.7400 1703.9400 1735.3400 1704.4200 ;
        RECT 1733.7400 1709.3800 1735.3400 1709.8600 ;
        RECT 1740.9000 1687.6200 1742.5000 1688.1000 ;
        RECT 1740.9000 1693.0600 1742.5000 1693.5400 ;
        RECT 1733.7400 1687.6200 1735.3400 1688.1000 ;
        RECT 1733.7400 1693.0600 1735.3400 1693.5400 ;
        RECT 1740.9000 1671.3000 1742.5000 1671.7800 ;
        RECT 1740.9000 1676.7400 1742.5000 1677.2200 ;
        RECT 1740.9000 1682.1800 1742.5000 1682.6600 ;
        RECT 1733.7400 1671.3000 1735.3400 1671.7800 ;
        RECT 1733.7400 1676.7400 1735.3400 1677.2200 ;
        RECT 1733.7400 1682.1800 1735.3400 1682.6600 ;
        RECT 1733.7400 1725.7000 1735.3400 1726.1800 ;
        RECT 1740.9000 1725.7000 1742.5000 1726.1800 ;
        RECT 1785.9000 1725.7000 1787.5000 1726.1800 ;
        RECT 1830.9000 1725.7000 1832.5000 1726.1800 ;
        RECT 1936.4400 1660.4200 1938.0400 1660.9000 ;
        RECT 1936.4400 1665.8600 1938.0400 1666.3400 ;
        RECT 1920.9000 1660.4200 1922.5000 1660.9000 ;
        RECT 1920.9000 1665.8600 1922.5000 1666.3400 ;
        RECT 1936.4400 1644.1000 1938.0400 1644.5800 ;
        RECT 1936.4400 1649.5400 1938.0400 1650.0200 ;
        RECT 1936.4400 1654.9800 1938.0400 1655.4600 ;
        RECT 1920.9000 1644.1000 1922.5000 1644.5800 ;
        RECT 1920.9000 1649.5400 1922.5000 1650.0200 ;
        RECT 1920.9000 1654.9800 1922.5000 1655.4600 ;
        RECT 1936.4400 1633.2200 1938.0400 1633.7000 ;
        RECT 1936.4400 1638.6600 1938.0400 1639.1400 ;
        RECT 1920.9000 1633.2200 1922.5000 1633.7000 ;
        RECT 1920.9000 1638.6600 1922.5000 1639.1400 ;
        RECT 1936.4400 1616.9000 1938.0400 1617.3800 ;
        RECT 1936.4400 1622.3400 1938.0400 1622.8200 ;
        RECT 1936.4400 1627.7800 1938.0400 1628.2600 ;
        RECT 1920.9000 1616.9000 1922.5000 1617.3800 ;
        RECT 1920.9000 1622.3400 1922.5000 1622.8200 ;
        RECT 1920.9000 1627.7800 1922.5000 1628.2600 ;
        RECT 1875.9000 1660.4200 1877.5000 1660.9000 ;
        RECT 1875.9000 1665.8600 1877.5000 1666.3400 ;
        RECT 1875.9000 1644.1000 1877.5000 1644.5800 ;
        RECT 1875.9000 1649.5400 1877.5000 1650.0200 ;
        RECT 1875.9000 1654.9800 1877.5000 1655.4600 ;
        RECT 1875.9000 1633.2200 1877.5000 1633.7000 ;
        RECT 1875.9000 1638.6600 1877.5000 1639.1400 ;
        RECT 1875.9000 1616.9000 1877.5000 1617.3800 ;
        RECT 1875.9000 1622.3400 1877.5000 1622.8200 ;
        RECT 1875.9000 1627.7800 1877.5000 1628.2600 ;
        RECT 1936.4400 1606.0200 1938.0400 1606.5000 ;
        RECT 1936.4400 1611.4600 1938.0400 1611.9400 ;
        RECT 1920.9000 1606.0200 1922.5000 1606.5000 ;
        RECT 1920.9000 1611.4600 1922.5000 1611.9400 ;
        RECT 1936.4400 1589.7000 1938.0400 1590.1800 ;
        RECT 1936.4400 1595.1400 1938.0400 1595.6200 ;
        RECT 1936.4400 1600.5800 1938.0400 1601.0600 ;
        RECT 1920.9000 1589.7000 1922.5000 1590.1800 ;
        RECT 1920.9000 1595.1400 1922.5000 1595.6200 ;
        RECT 1920.9000 1600.5800 1922.5000 1601.0600 ;
        RECT 1936.4400 1578.8200 1938.0400 1579.3000 ;
        RECT 1936.4400 1584.2600 1938.0400 1584.7400 ;
        RECT 1920.9000 1578.8200 1922.5000 1579.3000 ;
        RECT 1920.9000 1584.2600 1922.5000 1584.7400 ;
        RECT 1920.9000 1573.3800 1922.5000 1573.8600 ;
        RECT 1936.4400 1573.3800 1938.0400 1573.8600 ;
        RECT 1875.9000 1606.0200 1877.5000 1606.5000 ;
        RECT 1875.9000 1611.4600 1877.5000 1611.9400 ;
        RECT 1875.9000 1589.7000 1877.5000 1590.1800 ;
        RECT 1875.9000 1595.1400 1877.5000 1595.6200 ;
        RECT 1875.9000 1600.5800 1877.5000 1601.0600 ;
        RECT 1875.9000 1578.8200 1877.5000 1579.3000 ;
        RECT 1875.9000 1584.2600 1877.5000 1584.7400 ;
        RECT 1875.9000 1573.3800 1877.5000 1573.8600 ;
        RECT 1830.9000 1660.4200 1832.5000 1660.9000 ;
        RECT 1830.9000 1665.8600 1832.5000 1666.3400 ;
        RECT 1830.9000 1644.1000 1832.5000 1644.5800 ;
        RECT 1830.9000 1649.5400 1832.5000 1650.0200 ;
        RECT 1830.9000 1654.9800 1832.5000 1655.4600 ;
        RECT 1785.9000 1660.4200 1787.5000 1660.9000 ;
        RECT 1785.9000 1665.8600 1787.5000 1666.3400 ;
        RECT 1785.9000 1644.1000 1787.5000 1644.5800 ;
        RECT 1785.9000 1649.5400 1787.5000 1650.0200 ;
        RECT 1785.9000 1654.9800 1787.5000 1655.4600 ;
        RECT 1830.9000 1633.2200 1832.5000 1633.7000 ;
        RECT 1830.9000 1638.6600 1832.5000 1639.1400 ;
        RECT 1830.9000 1616.9000 1832.5000 1617.3800 ;
        RECT 1830.9000 1622.3400 1832.5000 1622.8200 ;
        RECT 1830.9000 1627.7800 1832.5000 1628.2600 ;
        RECT 1785.9000 1633.2200 1787.5000 1633.7000 ;
        RECT 1785.9000 1638.6600 1787.5000 1639.1400 ;
        RECT 1785.9000 1616.9000 1787.5000 1617.3800 ;
        RECT 1785.9000 1622.3400 1787.5000 1622.8200 ;
        RECT 1785.9000 1627.7800 1787.5000 1628.2600 ;
        RECT 1740.9000 1660.4200 1742.5000 1660.9000 ;
        RECT 1740.9000 1665.8600 1742.5000 1666.3400 ;
        RECT 1733.7400 1660.4200 1735.3400 1660.9000 ;
        RECT 1733.7400 1665.8600 1735.3400 1666.3400 ;
        RECT 1740.9000 1644.1000 1742.5000 1644.5800 ;
        RECT 1740.9000 1649.5400 1742.5000 1650.0200 ;
        RECT 1740.9000 1654.9800 1742.5000 1655.4600 ;
        RECT 1733.7400 1644.1000 1735.3400 1644.5800 ;
        RECT 1733.7400 1649.5400 1735.3400 1650.0200 ;
        RECT 1733.7400 1654.9800 1735.3400 1655.4600 ;
        RECT 1740.9000 1633.2200 1742.5000 1633.7000 ;
        RECT 1740.9000 1638.6600 1742.5000 1639.1400 ;
        RECT 1733.7400 1633.2200 1735.3400 1633.7000 ;
        RECT 1733.7400 1638.6600 1735.3400 1639.1400 ;
        RECT 1740.9000 1616.9000 1742.5000 1617.3800 ;
        RECT 1740.9000 1622.3400 1742.5000 1622.8200 ;
        RECT 1740.9000 1627.7800 1742.5000 1628.2600 ;
        RECT 1733.7400 1616.9000 1735.3400 1617.3800 ;
        RECT 1733.7400 1622.3400 1735.3400 1622.8200 ;
        RECT 1733.7400 1627.7800 1735.3400 1628.2600 ;
        RECT 1830.9000 1606.0200 1832.5000 1606.5000 ;
        RECT 1830.9000 1611.4600 1832.5000 1611.9400 ;
        RECT 1830.9000 1589.7000 1832.5000 1590.1800 ;
        RECT 1830.9000 1595.1400 1832.5000 1595.6200 ;
        RECT 1830.9000 1600.5800 1832.5000 1601.0600 ;
        RECT 1785.9000 1606.0200 1787.5000 1606.5000 ;
        RECT 1785.9000 1611.4600 1787.5000 1611.9400 ;
        RECT 1785.9000 1589.7000 1787.5000 1590.1800 ;
        RECT 1785.9000 1595.1400 1787.5000 1595.6200 ;
        RECT 1785.9000 1600.5800 1787.5000 1601.0600 ;
        RECT 1830.9000 1584.2600 1832.5000 1584.7400 ;
        RECT 1830.9000 1578.8200 1832.5000 1579.3000 ;
        RECT 1830.9000 1573.3800 1832.5000 1573.8600 ;
        RECT 1785.9000 1584.2600 1787.5000 1584.7400 ;
        RECT 1785.9000 1578.8200 1787.5000 1579.3000 ;
        RECT 1785.9000 1573.3800 1787.5000 1573.8600 ;
        RECT 1740.9000 1606.0200 1742.5000 1606.5000 ;
        RECT 1740.9000 1611.4600 1742.5000 1611.9400 ;
        RECT 1733.7400 1606.0200 1735.3400 1606.5000 ;
        RECT 1733.7400 1611.4600 1735.3400 1611.9400 ;
        RECT 1740.9000 1589.7000 1742.5000 1590.1800 ;
        RECT 1740.9000 1595.1400 1742.5000 1595.6200 ;
        RECT 1740.9000 1600.5800 1742.5000 1601.0600 ;
        RECT 1733.7400 1589.7000 1735.3400 1590.1800 ;
        RECT 1733.7400 1595.1400 1735.3400 1595.6200 ;
        RECT 1733.7400 1600.5800 1735.3400 1601.0600 ;
        RECT 1740.9000 1578.8200 1742.5000 1579.3000 ;
        RECT 1740.9000 1584.2600 1742.5000 1584.7400 ;
        RECT 1733.7400 1578.8200 1735.3400 1579.3000 ;
        RECT 1733.7400 1584.2600 1735.3400 1584.7400 ;
        RECT 1733.7400 1573.3800 1735.3400 1573.8600 ;
        RECT 1740.9000 1573.3800 1742.5000 1573.8600 ;
        RECT 1730.7800 1775.5700 1941.0000 1777.1700 ;
        RECT 1730.7800 1563.8700 1941.0000 1565.4700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1561.0400 1735.3400 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1779.0800 1735.3400 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1561.0400 1938.0400 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1779.0800 1938.0400 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1563.8700 1732.3800 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1563.8700 1941.0000 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1775.5700 1732.3800 1777.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1775.5700 1941.0000 1777.1700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 1334.2300 1922.5000 1547.5300 ;
        RECT 1875.9000 1334.2300 1877.5000 1547.5300 ;
        RECT 1830.9000 1334.2300 1832.5000 1547.5300 ;
        RECT 1785.9000 1334.2300 1787.5000 1547.5300 ;
        RECT 1740.9000 1334.2300 1742.5000 1547.5300 ;
        RECT 1936.4400 1331.4000 1938.0400 1551.0400 ;
        RECT 1733.7400 1331.4000 1735.3400 1551.0400 ;
      LAYER met3 ;
        RECT 1920.9000 1539.5800 1922.5000 1540.0600 ;
        RECT 1936.4400 1539.5800 1938.0400 1540.0600 ;
        RECT 1936.4400 1528.7000 1938.0400 1529.1800 ;
        RECT 1936.4400 1534.1400 1938.0400 1534.6200 ;
        RECT 1920.9000 1528.7000 1922.5000 1529.1800 ;
        RECT 1920.9000 1534.1400 1922.5000 1534.6200 ;
        RECT 1936.4400 1512.3800 1938.0400 1512.8600 ;
        RECT 1936.4400 1517.8200 1938.0400 1518.3000 ;
        RECT 1920.9000 1512.3800 1922.5000 1512.8600 ;
        RECT 1920.9000 1517.8200 1922.5000 1518.3000 ;
        RECT 1936.4400 1501.5000 1938.0400 1501.9800 ;
        RECT 1936.4400 1506.9400 1938.0400 1507.4200 ;
        RECT 1920.9000 1501.5000 1922.5000 1501.9800 ;
        RECT 1920.9000 1506.9400 1922.5000 1507.4200 ;
        RECT 1920.9000 1523.2600 1922.5000 1523.7400 ;
        RECT 1936.4400 1523.2600 1938.0400 1523.7400 ;
        RECT 1875.9000 1528.7000 1877.5000 1529.1800 ;
        RECT 1875.9000 1534.1400 1877.5000 1534.6200 ;
        RECT 1875.9000 1539.5800 1877.5000 1540.0600 ;
        RECT 1875.9000 1512.3800 1877.5000 1512.8600 ;
        RECT 1875.9000 1517.8200 1877.5000 1518.3000 ;
        RECT 1875.9000 1506.9400 1877.5000 1507.4200 ;
        RECT 1875.9000 1501.5000 1877.5000 1501.9800 ;
        RECT 1875.9000 1523.2600 1877.5000 1523.7400 ;
        RECT 1936.4400 1485.1800 1938.0400 1485.6600 ;
        RECT 1936.4400 1490.6200 1938.0400 1491.1000 ;
        RECT 1920.9000 1485.1800 1922.5000 1485.6600 ;
        RECT 1920.9000 1490.6200 1922.5000 1491.1000 ;
        RECT 1936.4400 1468.8600 1938.0400 1469.3400 ;
        RECT 1936.4400 1474.3000 1938.0400 1474.7800 ;
        RECT 1936.4400 1479.7400 1938.0400 1480.2200 ;
        RECT 1920.9000 1468.8600 1922.5000 1469.3400 ;
        RECT 1920.9000 1474.3000 1922.5000 1474.7800 ;
        RECT 1920.9000 1479.7400 1922.5000 1480.2200 ;
        RECT 1936.4400 1457.9800 1938.0400 1458.4600 ;
        RECT 1936.4400 1463.4200 1938.0400 1463.9000 ;
        RECT 1920.9000 1457.9800 1922.5000 1458.4600 ;
        RECT 1920.9000 1463.4200 1922.5000 1463.9000 ;
        RECT 1936.4400 1441.6600 1938.0400 1442.1400 ;
        RECT 1936.4400 1447.1000 1938.0400 1447.5800 ;
        RECT 1936.4400 1452.5400 1938.0400 1453.0200 ;
        RECT 1920.9000 1441.6600 1922.5000 1442.1400 ;
        RECT 1920.9000 1447.1000 1922.5000 1447.5800 ;
        RECT 1920.9000 1452.5400 1922.5000 1453.0200 ;
        RECT 1875.9000 1485.1800 1877.5000 1485.6600 ;
        RECT 1875.9000 1490.6200 1877.5000 1491.1000 ;
        RECT 1875.9000 1468.8600 1877.5000 1469.3400 ;
        RECT 1875.9000 1474.3000 1877.5000 1474.7800 ;
        RECT 1875.9000 1479.7400 1877.5000 1480.2200 ;
        RECT 1875.9000 1457.9800 1877.5000 1458.4600 ;
        RECT 1875.9000 1463.4200 1877.5000 1463.9000 ;
        RECT 1875.9000 1441.6600 1877.5000 1442.1400 ;
        RECT 1875.9000 1447.1000 1877.5000 1447.5800 ;
        RECT 1875.9000 1452.5400 1877.5000 1453.0200 ;
        RECT 1875.9000 1496.0600 1877.5000 1496.5400 ;
        RECT 1920.9000 1496.0600 1922.5000 1496.5400 ;
        RECT 1936.4400 1496.0600 1938.0400 1496.5400 ;
        RECT 1830.9000 1528.7000 1832.5000 1529.1800 ;
        RECT 1830.9000 1534.1400 1832.5000 1534.6200 ;
        RECT 1830.9000 1539.5800 1832.5000 1540.0600 ;
        RECT 1785.9000 1528.7000 1787.5000 1529.1800 ;
        RECT 1785.9000 1534.1400 1787.5000 1534.6200 ;
        RECT 1785.9000 1539.5800 1787.5000 1540.0600 ;
        RECT 1830.9000 1512.3800 1832.5000 1512.8600 ;
        RECT 1830.9000 1517.8200 1832.5000 1518.3000 ;
        RECT 1830.9000 1501.5000 1832.5000 1501.9800 ;
        RECT 1830.9000 1506.9400 1832.5000 1507.4200 ;
        RECT 1785.9000 1512.3800 1787.5000 1512.8600 ;
        RECT 1785.9000 1517.8200 1787.5000 1518.3000 ;
        RECT 1785.9000 1501.5000 1787.5000 1501.9800 ;
        RECT 1785.9000 1506.9400 1787.5000 1507.4200 ;
        RECT 1785.9000 1523.2600 1787.5000 1523.7400 ;
        RECT 1830.9000 1523.2600 1832.5000 1523.7400 ;
        RECT 1733.7400 1539.5800 1735.3400 1540.0600 ;
        RECT 1740.9000 1539.5800 1742.5000 1540.0600 ;
        RECT 1740.9000 1528.7000 1742.5000 1529.1800 ;
        RECT 1740.9000 1534.1400 1742.5000 1534.6200 ;
        RECT 1733.7400 1528.7000 1735.3400 1529.1800 ;
        RECT 1733.7400 1534.1400 1735.3400 1534.6200 ;
        RECT 1740.9000 1512.3800 1742.5000 1512.8600 ;
        RECT 1740.9000 1517.8200 1742.5000 1518.3000 ;
        RECT 1733.7400 1512.3800 1735.3400 1512.8600 ;
        RECT 1733.7400 1517.8200 1735.3400 1518.3000 ;
        RECT 1740.9000 1501.5000 1742.5000 1501.9800 ;
        RECT 1740.9000 1506.9400 1742.5000 1507.4200 ;
        RECT 1733.7400 1501.5000 1735.3400 1501.9800 ;
        RECT 1733.7400 1506.9400 1735.3400 1507.4200 ;
        RECT 1733.7400 1523.2600 1735.3400 1523.7400 ;
        RECT 1740.9000 1523.2600 1742.5000 1523.7400 ;
        RECT 1830.9000 1485.1800 1832.5000 1485.6600 ;
        RECT 1830.9000 1490.6200 1832.5000 1491.1000 ;
        RECT 1830.9000 1468.8600 1832.5000 1469.3400 ;
        RECT 1830.9000 1474.3000 1832.5000 1474.7800 ;
        RECT 1830.9000 1479.7400 1832.5000 1480.2200 ;
        RECT 1785.9000 1485.1800 1787.5000 1485.6600 ;
        RECT 1785.9000 1490.6200 1787.5000 1491.1000 ;
        RECT 1785.9000 1468.8600 1787.5000 1469.3400 ;
        RECT 1785.9000 1474.3000 1787.5000 1474.7800 ;
        RECT 1785.9000 1479.7400 1787.5000 1480.2200 ;
        RECT 1830.9000 1457.9800 1832.5000 1458.4600 ;
        RECT 1830.9000 1463.4200 1832.5000 1463.9000 ;
        RECT 1830.9000 1441.6600 1832.5000 1442.1400 ;
        RECT 1830.9000 1447.1000 1832.5000 1447.5800 ;
        RECT 1830.9000 1452.5400 1832.5000 1453.0200 ;
        RECT 1785.9000 1457.9800 1787.5000 1458.4600 ;
        RECT 1785.9000 1463.4200 1787.5000 1463.9000 ;
        RECT 1785.9000 1441.6600 1787.5000 1442.1400 ;
        RECT 1785.9000 1447.1000 1787.5000 1447.5800 ;
        RECT 1785.9000 1452.5400 1787.5000 1453.0200 ;
        RECT 1740.9000 1485.1800 1742.5000 1485.6600 ;
        RECT 1740.9000 1490.6200 1742.5000 1491.1000 ;
        RECT 1733.7400 1485.1800 1735.3400 1485.6600 ;
        RECT 1733.7400 1490.6200 1735.3400 1491.1000 ;
        RECT 1740.9000 1468.8600 1742.5000 1469.3400 ;
        RECT 1740.9000 1474.3000 1742.5000 1474.7800 ;
        RECT 1740.9000 1479.7400 1742.5000 1480.2200 ;
        RECT 1733.7400 1468.8600 1735.3400 1469.3400 ;
        RECT 1733.7400 1474.3000 1735.3400 1474.7800 ;
        RECT 1733.7400 1479.7400 1735.3400 1480.2200 ;
        RECT 1740.9000 1457.9800 1742.5000 1458.4600 ;
        RECT 1740.9000 1463.4200 1742.5000 1463.9000 ;
        RECT 1733.7400 1457.9800 1735.3400 1458.4600 ;
        RECT 1733.7400 1463.4200 1735.3400 1463.9000 ;
        RECT 1740.9000 1441.6600 1742.5000 1442.1400 ;
        RECT 1740.9000 1447.1000 1742.5000 1447.5800 ;
        RECT 1740.9000 1452.5400 1742.5000 1453.0200 ;
        RECT 1733.7400 1441.6600 1735.3400 1442.1400 ;
        RECT 1733.7400 1447.1000 1735.3400 1447.5800 ;
        RECT 1733.7400 1452.5400 1735.3400 1453.0200 ;
        RECT 1733.7400 1496.0600 1735.3400 1496.5400 ;
        RECT 1740.9000 1496.0600 1742.5000 1496.5400 ;
        RECT 1785.9000 1496.0600 1787.5000 1496.5400 ;
        RECT 1830.9000 1496.0600 1832.5000 1496.5400 ;
        RECT 1936.4400 1430.7800 1938.0400 1431.2600 ;
        RECT 1936.4400 1436.2200 1938.0400 1436.7000 ;
        RECT 1920.9000 1430.7800 1922.5000 1431.2600 ;
        RECT 1920.9000 1436.2200 1922.5000 1436.7000 ;
        RECT 1936.4400 1414.4600 1938.0400 1414.9400 ;
        RECT 1936.4400 1419.9000 1938.0400 1420.3800 ;
        RECT 1936.4400 1425.3400 1938.0400 1425.8200 ;
        RECT 1920.9000 1414.4600 1922.5000 1414.9400 ;
        RECT 1920.9000 1419.9000 1922.5000 1420.3800 ;
        RECT 1920.9000 1425.3400 1922.5000 1425.8200 ;
        RECT 1936.4400 1403.5800 1938.0400 1404.0600 ;
        RECT 1936.4400 1409.0200 1938.0400 1409.5000 ;
        RECT 1920.9000 1403.5800 1922.5000 1404.0600 ;
        RECT 1920.9000 1409.0200 1922.5000 1409.5000 ;
        RECT 1936.4400 1387.2600 1938.0400 1387.7400 ;
        RECT 1936.4400 1392.7000 1938.0400 1393.1800 ;
        RECT 1936.4400 1398.1400 1938.0400 1398.6200 ;
        RECT 1920.9000 1387.2600 1922.5000 1387.7400 ;
        RECT 1920.9000 1392.7000 1922.5000 1393.1800 ;
        RECT 1920.9000 1398.1400 1922.5000 1398.6200 ;
        RECT 1875.9000 1430.7800 1877.5000 1431.2600 ;
        RECT 1875.9000 1436.2200 1877.5000 1436.7000 ;
        RECT 1875.9000 1414.4600 1877.5000 1414.9400 ;
        RECT 1875.9000 1419.9000 1877.5000 1420.3800 ;
        RECT 1875.9000 1425.3400 1877.5000 1425.8200 ;
        RECT 1875.9000 1403.5800 1877.5000 1404.0600 ;
        RECT 1875.9000 1409.0200 1877.5000 1409.5000 ;
        RECT 1875.9000 1387.2600 1877.5000 1387.7400 ;
        RECT 1875.9000 1392.7000 1877.5000 1393.1800 ;
        RECT 1875.9000 1398.1400 1877.5000 1398.6200 ;
        RECT 1936.4400 1376.3800 1938.0400 1376.8600 ;
        RECT 1936.4400 1381.8200 1938.0400 1382.3000 ;
        RECT 1920.9000 1376.3800 1922.5000 1376.8600 ;
        RECT 1920.9000 1381.8200 1922.5000 1382.3000 ;
        RECT 1936.4400 1360.0600 1938.0400 1360.5400 ;
        RECT 1936.4400 1365.5000 1938.0400 1365.9800 ;
        RECT 1936.4400 1370.9400 1938.0400 1371.4200 ;
        RECT 1920.9000 1360.0600 1922.5000 1360.5400 ;
        RECT 1920.9000 1365.5000 1922.5000 1365.9800 ;
        RECT 1920.9000 1370.9400 1922.5000 1371.4200 ;
        RECT 1936.4400 1349.1800 1938.0400 1349.6600 ;
        RECT 1936.4400 1354.6200 1938.0400 1355.1000 ;
        RECT 1920.9000 1349.1800 1922.5000 1349.6600 ;
        RECT 1920.9000 1354.6200 1922.5000 1355.1000 ;
        RECT 1920.9000 1343.7400 1922.5000 1344.2200 ;
        RECT 1936.4400 1343.7400 1938.0400 1344.2200 ;
        RECT 1875.9000 1376.3800 1877.5000 1376.8600 ;
        RECT 1875.9000 1381.8200 1877.5000 1382.3000 ;
        RECT 1875.9000 1360.0600 1877.5000 1360.5400 ;
        RECT 1875.9000 1365.5000 1877.5000 1365.9800 ;
        RECT 1875.9000 1370.9400 1877.5000 1371.4200 ;
        RECT 1875.9000 1349.1800 1877.5000 1349.6600 ;
        RECT 1875.9000 1354.6200 1877.5000 1355.1000 ;
        RECT 1875.9000 1343.7400 1877.5000 1344.2200 ;
        RECT 1830.9000 1430.7800 1832.5000 1431.2600 ;
        RECT 1830.9000 1436.2200 1832.5000 1436.7000 ;
        RECT 1830.9000 1414.4600 1832.5000 1414.9400 ;
        RECT 1830.9000 1419.9000 1832.5000 1420.3800 ;
        RECT 1830.9000 1425.3400 1832.5000 1425.8200 ;
        RECT 1785.9000 1430.7800 1787.5000 1431.2600 ;
        RECT 1785.9000 1436.2200 1787.5000 1436.7000 ;
        RECT 1785.9000 1414.4600 1787.5000 1414.9400 ;
        RECT 1785.9000 1419.9000 1787.5000 1420.3800 ;
        RECT 1785.9000 1425.3400 1787.5000 1425.8200 ;
        RECT 1830.9000 1403.5800 1832.5000 1404.0600 ;
        RECT 1830.9000 1409.0200 1832.5000 1409.5000 ;
        RECT 1830.9000 1387.2600 1832.5000 1387.7400 ;
        RECT 1830.9000 1392.7000 1832.5000 1393.1800 ;
        RECT 1830.9000 1398.1400 1832.5000 1398.6200 ;
        RECT 1785.9000 1403.5800 1787.5000 1404.0600 ;
        RECT 1785.9000 1409.0200 1787.5000 1409.5000 ;
        RECT 1785.9000 1387.2600 1787.5000 1387.7400 ;
        RECT 1785.9000 1392.7000 1787.5000 1393.1800 ;
        RECT 1785.9000 1398.1400 1787.5000 1398.6200 ;
        RECT 1740.9000 1430.7800 1742.5000 1431.2600 ;
        RECT 1740.9000 1436.2200 1742.5000 1436.7000 ;
        RECT 1733.7400 1430.7800 1735.3400 1431.2600 ;
        RECT 1733.7400 1436.2200 1735.3400 1436.7000 ;
        RECT 1740.9000 1414.4600 1742.5000 1414.9400 ;
        RECT 1740.9000 1419.9000 1742.5000 1420.3800 ;
        RECT 1740.9000 1425.3400 1742.5000 1425.8200 ;
        RECT 1733.7400 1414.4600 1735.3400 1414.9400 ;
        RECT 1733.7400 1419.9000 1735.3400 1420.3800 ;
        RECT 1733.7400 1425.3400 1735.3400 1425.8200 ;
        RECT 1740.9000 1403.5800 1742.5000 1404.0600 ;
        RECT 1740.9000 1409.0200 1742.5000 1409.5000 ;
        RECT 1733.7400 1403.5800 1735.3400 1404.0600 ;
        RECT 1733.7400 1409.0200 1735.3400 1409.5000 ;
        RECT 1740.9000 1387.2600 1742.5000 1387.7400 ;
        RECT 1740.9000 1392.7000 1742.5000 1393.1800 ;
        RECT 1740.9000 1398.1400 1742.5000 1398.6200 ;
        RECT 1733.7400 1387.2600 1735.3400 1387.7400 ;
        RECT 1733.7400 1392.7000 1735.3400 1393.1800 ;
        RECT 1733.7400 1398.1400 1735.3400 1398.6200 ;
        RECT 1830.9000 1376.3800 1832.5000 1376.8600 ;
        RECT 1830.9000 1381.8200 1832.5000 1382.3000 ;
        RECT 1830.9000 1360.0600 1832.5000 1360.5400 ;
        RECT 1830.9000 1365.5000 1832.5000 1365.9800 ;
        RECT 1830.9000 1370.9400 1832.5000 1371.4200 ;
        RECT 1785.9000 1376.3800 1787.5000 1376.8600 ;
        RECT 1785.9000 1381.8200 1787.5000 1382.3000 ;
        RECT 1785.9000 1360.0600 1787.5000 1360.5400 ;
        RECT 1785.9000 1365.5000 1787.5000 1365.9800 ;
        RECT 1785.9000 1370.9400 1787.5000 1371.4200 ;
        RECT 1830.9000 1354.6200 1832.5000 1355.1000 ;
        RECT 1830.9000 1349.1800 1832.5000 1349.6600 ;
        RECT 1830.9000 1343.7400 1832.5000 1344.2200 ;
        RECT 1785.9000 1354.6200 1787.5000 1355.1000 ;
        RECT 1785.9000 1349.1800 1787.5000 1349.6600 ;
        RECT 1785.9000 1343.7400 1787.5000 1344.2200 ;
        RECT 1740.9000 1376.3800 1742.5000 1376.8600 ;
        RECT 1740.9000 1381.8200 1742.5000 1382.3000 ;
        RECT 1733.7400 1376.3800 1735.3400 1376.8600 ;
        RECT 1733.7400 1381.8200 1735.3400 1382.3000 ;
        RECT 1740.9000 1360.0600 1742.5000 1360.5400 ;
        RECT 1740.9000 1365.5000 1742.5000 1365.9800 ;
        RECT 1740.9000 1370.9400 1742.5000 1371.4200 ;
        RECT 1733.7400 1360.0600 1735.3400 1360.5400 ;
        RECT 1733.7400 1365.5000 1735.3400 1365.9800 ;
        RECT 1733.7400 1370.9400 1735.3400 1371.4200 ;
        RECT 1740.9000 1349.1800 1742.5000 1349.6600 ;
        RECT 1740.9000 1354.6200 1742.5000 1355.1000 ;
        RECT 1733.7400 1349.1800 1735.3400 1349.6600 ;
        RECT 1733.7400 1354.6200 1735.3400 1355.1000 ;
        RECT 1733.7400 1343.7400 1735.3400 1344.2200 ;
        RECT 1740.9000 1343.7400 1742.5000 1344.2200 ;
        RECT 1730.7800 1545.9300 1941.0000 1547.5300 ;
        RECT 1730.7800 1334.2300 1941.0000 1335.8300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1331.4000 1735.3400 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1549.4400 1735.3400 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1331.4000 1938.0400 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1549.4400 1938.0400 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1334.2300 1732.3800 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1334.2300 1941.0000 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1545.9300 1732.3800 1547.5300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1545.9300 1941.0000 1547.5300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 1104.5900 1922.5000 1317.8900 ;
        RECT 1875.9000 1104.5900 1877.5000 1317.8900 ;
        RECT 1830.9000 1104.5900 1832.5000 1317.8900 ;
        RECT 1785.9000 1104.5900 1787.5000 1317.8900 ;
        RECT 1740.9000 1104.5900 1742.5000 1317.8900 ;
        RECT 1936.4400 1101.7600 1938.0400 1321.4000 ;
        RECT 1733.7400 1101.7600 1735.3400 1321.4000 ;
      LAYER met3 ;
        RECT 1920.9000 1309.9400 1922.5000 1310.4200 ;
        RECT 1936.4400 1309.9400 1938.0400 1310.4200 ;
        RECT 1936.4400 1299.0600 1938.0400 1299.5400 ;
        RECT 1936.4400 1304.5000 1938.0400 1304.9800 ;
        RECT 1920.9000 1299.0600 1922.5000 1299.5400 ;
        RECT 1920.9000 1304.5000 1922.5000 1304.9800 ;
        RECT 1936.4400 1282.7400 1938.0400 1283.2200 ;
        RECT 1936.4400 1288.1800 1938.0400 1288.6600 ;
        RECT 1920.9000 1282.7400 1922.5000 1283.2200 ;
        RECT 1920.9000 1288.1800 1922.5000 1288.6600 ;
        RECT 1936.4400 1271.8600 1938.0400 1272.3400 ;
        RECT 1936.4400 1277.3000 1938.0400 1277.7800 ;
        RECT 1920.9000 1271.8600 1922.5000 1272.3400 ;
        RECT 1920.9000 1277.3000 1922.5000 1277.7800 ;
        RECT 1920.9000 1293.6200 1922.5000 1294.1000 ;
        RECT 1936.4400 1293.6200 1938.0400 1294.1000 ;
        RECT 1875.9000 1299.0600 1877.5000 1299.5400 ;
        RECT 1875.9000 1304.5000 1877.5000 1304.9800 ;
        RECT 1875.9000 1309.9400 1877.5000 1310.4200 ;
        RECT 1875.9000 1282.7400 1877.5000 1283.2200 ;
        RECT 1875.9000 1288.1800 1877.5000 1288.6600 ;
        RECT 1875.9000 1277.3000 1877.5000 1277.7800 ;
        RECT 1875.9000 1271.8600 1877.5000 1272.3400 ;
        RECT 1875.9000 1293.6200 1877.5000 1294.1000 ;
        RECT 1936.4400 1255.5400 1938.0400 1256.0200 ;
        RECT 1936.4400 1260.9800 1938.0400 1261.4600 ;
        RECT 1920.9000 1255.5400 1922.5000 1256.0200 ;
        RECT 1920.9000 1260.9800 1922.5000 1261.4600 ;
        RECT 1936.4400 1239.2200 1938.0400 1239.7000 ;
        RECT 1936.4400 1244.6600 1938.0400 1245.1400 ;
        RECT 1936.4400 1250.1000 1938.0400 1250.5800 ;
        RECT 1920.9000 1239.2200 1922.5000 1239.7000 ;
        RECT 1920.9000 1244.6600 1922.5000 1245.1400 ;
        RECT 1920.9000 1250.1000 1922.5000 1250.5800 ;
        RECT 1936.4400 1228.3400 1938.0400 1228.8200 ;
        RECT 1936.4400 1233.7800 1938.0400 1234.2600 ;
        RECT 1920.9000 1228.3400 1922.5000 1228.8200 ;
        RECT 1920.9000 1233.7800 1922.5000 1234.2600 ;
        RECT 1936.4400 1212.0200 1938.0400 1212.5000 ;
        RECT 1936.4400 1217.4600 1938.0400 1217.9400 ;
        RECT 1936.4400 1222.9000 1938.0400 1223.3800 ;
        RECT 1920.9000 1212.0200 1922.5000 1212.5000 ;
        RECT 1920.9000 1217.4600 1922.5000 1217.9400 ;
        RECT 1920.9000 1222.9000 1922.5000 1223.3800 ;
        RECT 1875.9000 1255.5400 1877.5000 1256.0200 ;
        RECT 1875.9000 1260.9800 1877.5000 1261.4600 ;
        RECT 1875.9000 1239.2200 1877.5000 1239.7000 ;
        RECT 1875.9000 1244.6600 1877.5000 1245.1400 ;
        RECT 1875.9000 1250.1000 1877.5000 1250.5800 ;
        RECT 1875.9000 1228.3400 1877.5000 1228.8200 ;
        RECT 1875.9000 1233.7800 1877.5000 1234.2600 ;
        RECT 1875.9000 1212.0200 1877.5000 1212.5000 ;
        RECT 1875.9000 1217.4600 1877.5000 1217.9400 ;
        RECT 1875.9000 1222.9000 1877.5000 1223.3800 ;
        RECT 1875.9000 1266.4200 1877.5000 1266.9000 ;
        RECT 1920.9000 1266.4200 1922.5000 1266.9000 ;
        RECT 1936.4400 1266.4200 1938.0400 1266.9000 ;
        RECT 1830.9000 1299.0600 1832.5000 1299.5400 ;
        RECT 1830.9000 1304.5000 1832.5000 1304.9800 ;
        RECT 1830.9000 1309.9400 1832.5000 1310.4200 ;
        RECT 1785.9000 1299.0600 1787.5000 1299.5400 ;
        RECT 1785.9000 1304.5000 1787.5000 1304.9800 ;
        RECT 1785.9000 1309.9400 1787.5000 1310.4200 ;
        RECT 1830.9000 1282.7400 1832.5000 1283.2200 ;
        RECT 1830.9000 1288.1800 1832.5000 1288.6600 ;
        RECT 1830.9000 1271.8600 1832.5000 1272.3400 ;
        RECT 1830.9000 1277.3000 1832.5000 1277.7800 ;
        RECT 1785.9000 1282.7400 1787.5000 1283.2200 ;
        RECT 1785.9000 1288.1800 1787.5000 1288.6600 ;
        RECT 1785.9000 1271.8600 1787.5000 1272.3400 ;
        RECT 1785.9000 1277.3000 1787.5000 1277.7800 ;
        RECT 1785.9000 1293.6200 1787.5000 1294.1000 ;
        RECT 1830.9000 1293.6200 1832.5000 1294.1000 ;
        RECT 1733.7400 1309.9400 1735.3400 1310.4200 ;
        RECT 1740.9000 1309.9400 1742.5000 1310.4200 ;
        RECT 1740.9000 1299.0600 1742.5000 1299.5400 ;
        RECT 1740.9000 1304.5000 1742.5000 1304.9800 ;
        RECT 1733.7400 1299.0600 1735.3400 1299.5400 ;
        RECT 1733.7400 1304.5000 1735.3400 1304.9800 ;
        RECT 1740.9000 1282.7400 1742.5000 1283.2200 ;
        RECT 1740.9000 1288.1800 1742.5000 1288.6600 ;
        RECT 1733.7400 1282.7400 1735.3400 1283.2200 ;
        RECT 1733.7400 1288.1800 1735.3400 1288.6600 ;
        RECT 1740.9000 1271.8600 1742.5000 1272.3400 ;
        RECT 1740.9000 1277.3000 1742.5000 1277.7800 ;
        RECT 1733.7400 1271.8600 1735.3400 1272.3400 ;
        RECT 1733.7400 1277.3000 1735.3400 1277.7800 ;
        RECT 1733.7400 1293.6200 1735.3400 1294.1000 ;
        RECT 1740.9000 1293.6200 1742.5000 1294.1000 ;
        RECT 1830.9000 1255.5400 1832.5000 1256.0200 ;
        RECT 1830.9000 1260.9800 1832.5000 1261.4600 ;
        RECT 1830.9000 1239.2200 1832.5000 1239.7000 ;
        RECT 1830.9000 1244.6600 1832.5000 1245.1400 ;
        RECT 1830.9000 1250.1000 1832.5000 1250.5800 ;
        RECT 1785.9000 1255.5400 1787.5000 1256.0200 ;
        RECT 1785.9000 1260.9800 1787.5000 1261.4600 ;
        RECT 1785.9000 1239.2200 1787.5000 1239.7000 ;
        RECT 1785.9000 1244.6600 1787.5000 1245.1400 ;
        RECT 1785.9000 1250.1000 1787.5000 1250.5800 ;
        RECT 1830.9000 1228.3400 1832.5000 1228.8200 ;
        RECT 1830.9000 1233.7800 1832.5000 1234.2600 ;
        RECT 1830.9000 1212.0200 1832.5000 1212.5000 ;
        RECT 1830.9000 1217.4600 1832.5000 1217.9400 ;
        RECT 1830.9000 1222.9000 1832.5000 1223.3800 ;
        RECT 1785.9000 1228.3400 1787.5000 1228.8200 ;
        RECT 1785.9000 1233.7800 1787.5000 1234.2600 ;
        RECT 1785.9000 1212.0200 1787.5000 1212.5000 ;
        RECT 1785.9000 1217.4600 1787.5000 1217.9400 ;
        RECT 1785.9000 1222.9000 1787.5000 1223.3800 ;
        RECT 1740.9000 1255.5400 1742.5000 1256.0200 ;
        RECT 1740.9000 1260.9800 1742.5000 1261.4600 ;
        RECT 1733.7400 1255.5400 1735.3400 1256.0200 ;
        RECT 1733.7400 1260.9800 1735.3400 1261.4600 ;
        RECT 1740.9000 1239.2200 1742.5000 1239.7000 ;
        RECT 1740.9000 1244.6600 1742.5000 1245.1400 ;
        RECT 1740.9000 1250.1000 1742.5000 1250.5800 ;
        RECT 1733.7400 1239.2200 1735.3400 1239.7000 ;
        RECT 1733.7400 1244.6600 1735.3400 1245.1400 ;
        RECT 1733.7400 1250.1000 1735.3400 1250.5800 ;
        RECT 1740.9000 1228.3400 1742.5000 1228.8200 ;
        RECT 1740.9000 1233.7800 1742.5000 1234.2600 ;
        RECT 1733.7400 1228.3400 1735.3400 1228.8200 ;
        RECT 1733.7400 1233.7800 1735.3400 1234.2600 ;
        RECT 1740.9000 1212.0200 1742.5000 1212.5000 ;
        RECT 1740.9000 1217.4600 1742.5000 1217.9400 ;
        RECT 1740.9000 1222.9000 1742.5000 1223.3800 ;
        RECT 1733.7400 1212.0200 1735.3400 1212.5000 ;
        RECT 1733.7400 1217.4600 1735.3400 1217.9400 ;
        RECT 1733.7400 1222.9000 1735.3400 1223.3800 ;
        RECT 1733.7400 1266.4200 1735.3400 1266.9000 ;
        RECT 1740.9000 1266.4200 1742.5000 1266.9000 ;
        RECT 1785.9000 1266.4200 1787.5000 1266.9000 ;
        RECT 1830.9000 1266.4200 1832.5000 1266.9000 ;
        RECT 1936.4400 1201.1400 1938.0400 1201.6200 ;
        RECT 1936.4400 1206.5800 1938.0400 1207.0600 ;
        RECT 1920.9000 1201.1400 1922.5000 1201.6200 ;
        RECT 1920.9000 1206.5800 1922.5000 1207.0600 ;
        RECT 1936.4400 1184.8200 1938.0400 1185.3000 ;
        RECT 1936.4400 1190.2600 1938.0400 1190.7400 ;
        RECT 1936.4400 1195.7000 1938.0400 1196.1800 ;
        RECT 1920.9000 1184.8200 1922.5000 1185.3000 ;
        RECT 1920.9000 1190.2600 1922.5000 1190.7400 ;
        RECT 1920.9000 1195.7000 1922.5000 1196.1800 ;
        RECT 1936.4400 1173.9400 1938.0400 1174.4200 ;
        RECT 1936.4400 1179.3800 1938.0400 1179.8600 ;
        RECT 1920.9000 1173.9400 1922.5000 1174.4200 ;
        RECT 1920.9000 1179.3800 1922.5000 1179.8600 ;
        RECT 1936.4400 1157.6200 1938.0400 1158.1000 ;
        RECT 1936.4400 1163.0600 1938.0400 1163.5400 ;
        RECT 1936.4400 1168.5000 1938.0400 1168.9800 ;
        RECT 1920.9000 1157.6200 1922.5000 1158.1000 ;
        RECT 1920.9000 1163.0600 1922.5000 1163.5400 ;
        RECT 1920.9000 1168.5000 1922.5000 1168.9800 ;
        RECT 1875.9000 1201.1400 1877.5000 1201.6200 ;
        RECT 1875.9000 1206.5800 1877.5000 1207.0600 ;
        RECT 1875.9000 1184.8200 1877.5000 1185.3000 ;
        RECT 1875.9000 1190.2600 1877.5000 1190.7400 ;
        RECT 1875.9000 1195.7000 1877.5000 1196.1800 ;
        RECT 1875.9000 1173.9400 1877.5000 1174.4200 ;
        RECT 1875.9000 1179.3800 1877.5000 1179.8600 ;
        RECT 1875.9000 1157.6200 1877.5000 1158.1000 ;
        RECT 1875.9000 1163.0600 1877.5000 1163.5400 ;
        RECT 1875.9000 1168.5000 1877.5000 1168.9800 ;
        RECT 1936.4400 1146.7400 1938.0400 1147.2200 ;
        RECT 1936.4400 1152.1800 1938.0400 1152.6600 ;
        RECT 1920.9000 1146.7400 1922.5000 1147.2200 ;
        RECT 1920.9000 1152.1800 1922.5000 1152.6600 ;
        RECT 1936.4400 1130.4200 1938.0400 1130.9000 ;
        RECT 1936.4400 1135.8600 1938.0400 1136.3400 ;
        RECT 1936.4400 1141.3000 1938.0400 1141.7800 ;
        RECT 1920.9000 1130.4200 1922.5000 1130.9000 ;
        RECT 1920.9000 1135.8600 1922.5000 1136.3400 ;
        RECT 1920.9000 1141.3000 1922.5000 1141.7800 ;
        RECT 1936.4400 1119.5400 1938.0400 1120.0200 ;
        RECT 1936.4400 1124.9800 1938.0400 1125.4600 ;
        RECT 1920.9000 1119.5400 1922.5000 1120.0200 ;
        RECT 1920.9000 1124.9800 1922.5000 1125.4600 ;
        RECT 1920.9000 1114.1000 1922.5000 1114.5800 ;
        RECT 1936.4400 1114.1000 1938.0400 1114.5800 ;
        RECT 1875.9000 1146.7400 1877.5000 1147.2200 ;
        RECT 1875.9000 1152.1800 1877.5000 1152.6600 ;
        RECT 1875.9000 1130.4200 1877.5000 1130.9000 ;
        RECT 1875.9000 1135.8600 1877.5000 1136.3400 ;
        RECT 1875.9000 1141.3000 1877.5000 1141.7800 ;
        RECT 1875.9000 1119.5400 1877.5000 1120.0200 ;
        RECT 1875.9000 1124.9800 1877.5000 1125.4600 ;
        RECT 1875.9000 1114.1000 1877.5000 1114.5800 ;
        RECT 1830.9000 1201.1400 1832.5000 1201.6200 ;
        RECT 1830.9000 1206.5800 1832.5000 1207.0600 ;
        RECT 1830.9000 1184.8200 1832.5000 1185.3000 ;
        RECT 1830.9000 1190.2600 1832.5000 1190.7400 ;
        RECT 1830.9000 1195.7000 1832.5000 1196.1800 ;
        RECT 1785.9000 1201.1400 1787.5000 1201.6200 ;
        RECT 1785.9000 1206.5800 1787.5000 1207.0600 ;
        RECT 1785.9000 1184.8200 1787.5000 1185.3000 ;
        RECT 1785.9000 1190.2600 1787.5000 1190.7400 ;
        RECT 1785.9000 1195.7000 1787.5000 1196.1800 ;
        RECT 1830.9000 1173.9400 1832.5000 1174.4200 ;
        RECT 1830.9000 1179.3800 1832.5000 1179.8600 ;
        RECT 1830.9000 1157.6200 1832.5000 1158.1000 ;
        RECT 1830.9000 1163.0600 1832.5000 1163.5400 ;
        RECT 1830.9000 1168.5000 1832.5000 1168.9800 ;
        RECT 1785.9000 1173.9400 1787.5000 1174.4200 ;
        RECT 1785.9000 1179.3800 1787.5000 1179.8600 ;
        RECT 1785.9000 1157.6200 1787.5000 1158.1000 ;
        RECT 1785.9000 1163.0600 1787.5000 1163.5400 ;
        RECT 1785.9000 1168.5000 1787.5000 1168.9800 ;
        RECT 1740.9000 1201.1400 1742.5000 1201.6200 ;
        RECT 1740.9000 1206.5800 1742.5000 1207.0600 ;
        RECT 1733.7400 1201.1400 1735.3400 1201.6200 ;
        RECT 1733.7400 1206.5800 1735.3400 1207.0600 ;
        RECT 1740.9000 1184.8200 1742.5000 1185.3000 ;
        RECT 1740.9000 1190.2600 1742.5000 1190.7400 ;
        RECT 1740.9000 1195.7000 1742.5000 1196.1800 ;
        RECT 1733.7400 1184.8200 1735.3400 1185.3000 ;
        RECT 1733.7400 1190.2600 1735.3400 1190.7400 ;
        RECT 1733.7400 1195.7000 1735.3400 1196.1800 ;
        RECT 1740.9000 1173.9400 1742.5000 1174.4200 ;
        RECT 1740.9000 1179.3800 1742.5000 1179.8600 ;
        RECT 1733.7400 1173.9400 1735.3400 1174.4200 ;
        RECT 1733.7400 1179.3800 1735.3400 1179.8600 ;
        RECT 1740.9000 1157.6200 1742.5000 1158.1000 ;
        RECT 1740.9000 1163.0600 1742.5000 1163.5400 ;
        RECT 1740.9000 1168.5000 1742.5000 1168.9800 ;
        RECT 1733.7400 1157.6200 1735.3400 1158.1000 ;
        RECT 1733.7400 1163.0600 1735.3400 1163.5400 ;
        RECT 1733.7400 1168.5000 1735.3400 1168.9800 ;
        RECT 1830.9000 1146.7400 1832.5000 1147.2200 ;
        RECT 1830.9000 1152.1800 1832.5000 1152.6600 ;
        RECT 1830.9000 1130.4200 1832.5000 1130.9000 ;
        RECT 1830.9000 1135.8600 1832.5000 1136.3400 ;
        RECT 1830.9000 1141.3000 1832.5000 1141.7800 ;
        RECT 1785.9000 1146.7400 1787.5000 1147.2200 ;
        RECT 1785.9000 1152.1800 1787.5000 1152.6600 ;
        RECT 1785.9000 1130.4200 1787.5000 1130.9000 ;
        RECT 1785.9000 1135.8600 1787.5000 1136.3400 ;
        RECT 1785.9000 1141.3000 1787.5000 1141.7800 ;
        RECT 1830.9000 1124.9800 1832.5000 1125.4600 ;
        RECT 1830.9000 1119.5400 1832.5000 1120.0200 ;
        RECT 1830.9000 1114.1000 1832.5000 1114.5800 ;
        RECT 1785.9000 1124.9800 1787.5000 1125.4600 ;
        RECT 1785.9000 1119.5400 1787.5000 1120.0200 ;
        RECT 1785.9000 1114.1000 1787.5000 1114.5800 ;
        RECT 1740.9000 1146.7400 1742.5000 1147.2200 ;
        RECT 1740.9000 1152.1800 1742.5000 1152.6600 ;
        RECT 1733.7400 1146.7400 1735.3400 1147.2200 ;
        RECT 1733.7400 1152.1800 1735.3400 1152.6600 ;
        RECT 1740.9000 1130.4200 1742.5000 1130.9000 ;
        RECT 1740.9000 1135.8600 1742.5000 1136.3400 ;
        RECT 1740.9000 1141.3000 1742.5000 1141.7800 ;
        RECT 1733.7400 1130.4200 1735.3400 1130.9000 ;
        RECT 1733.7400 1135.8600 1735.3400 1136.3400 ;
        RECT 1733.7400 1141.3000 1735.3400 1141.7800 ;
        RECT 1740.9000 1119.5400 1742.5000 1120.0200 ;
        RECT 1740.9000 1124.9800 1742.5000 1125.4600 ;
        RECT 1733.7400 1119.5400 1735.3400 1120.0200 ;
        RECT 1733.7400 1124.9800 1735.3400 1125.4600 ;
        RECT 1733.7400 1114.1000 1735.3400 1114.5800 ;
        RECT 1740.9000 1114.1000 1742.5000 1114.5800 ;
        RECT 1730.7800 1316.2900 1941.0000 1317.8900 ;
        RECT 1730.7800 1104.5900 1941.0000 1106.1900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1101.7600 1735.3400 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1319.8000 1735.3400 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1101.7600 1938.0400 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1319.8000 1938.0400 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1104.5900 1732.3800 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1104.5900 1941.0000 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1316.2900 1732.3800 1317.8900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1316.2900 1941.0000 1317.8900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 874.9500 1922.5000 1088.2500 ;
        RECT 1875.9000 874.9500 1877.5000 1088.2500 ;
        RECT 1830.9000 874.9500 1832.5000 1088.2500 ;
        RECT 1785.9000 874.9500 1787.5000 1088.2500 ;
        RECT 1740.9000 874.9500 1742.5000 1088.2500 ;
        RECT 1936.4400 872.1200 1938.0400 1091.7600 ;
        RECT 1733.7400 872.1200 1735.3400 1091.7600 ;
      LAYER met3 ;
        RECT 1920.9000 1080.3000 1922.5000 1080.7800 ;
        RECT 1936.4400 1080.3000 1938.0400 1080.7800 ;
        RECT 1936.4400 1069.4200 1938.0400 1069.9000 ;
        RECT 1936.4400 1074.8600 1938.0400 1075.3400 ;
        RECT 1920.9000 1069.4200 1922.5000 1069.9000 ;
        RECT 1920.9000 1074.8600 1922.5000 1075.3400 ;
        RECT 1936.4400 1053.1000 1938.0400 1053.5800 ;
        RECT 1936.4400 1058.5400 1938.0400 1059.0200 ;
        RECT 1920.9000 1053.1000 1922.5000 1053.5800 ;
        RECT 1920.9000 1058.5400 1922.5000 1059.0200 ;
        RECT 1936.4400 1042.2200 1938.0400 1042.7000 ;
        RECT 1936.4400 1047.6600 1938.0400 1048.1400 ;
        RECT 1920.9000 1042.2200 1922.5000 1042.7000 ;
        RECT 1920.9000 1047.6600 1922.5000 1048.1400 ;
        RECT 1920.9000 1063.9800 1922.5000 1064.4600 ;
        RECT 1936.4400 1063.9800 1938.0400 1064.4600 ;
        RECT 1875.9000 1069.4200 1877.5000 1069.9000 ;
        RECT 1875.9000 1074.8600 1877.5000 1075.3400 ;
        RECT 1875.9000 1080.3000 1877.5000 1080.7800 ;
        RECT 1875.9000 1053.1000 1877.5000 1053.5800 ;
        RECT 1875.9000 1058.5400 1877.5000 1059.0200 ;
        RECT 1875.9000 1047.6600 1877.5000 1048.1400 ;
        RECT 1875.9000 1042.2200 1877.5000 1042.7000 ;
        RECT 1875.9000 1063.9800 1877.5000 1064.4600 ;
        RECT 1936.4400 1025.9000 1938.0400 1026.3800 ;
        RECT 1936.4400 1031.3400 1938.0400 1031.8200 ;
        RECT 1920.9000 1025.9000 1922.5000 1026.3800 ;
        RECT 1920.9000 1031.3400 1922.5000 1031.8200 ;
        RECT 1936.4400 1009.5800 1938.0400 1010.0600 ;
        RECT 1936.4400 1015.0200 1938.0400 1015.5000 ;
        RECT 1936.4400 1020.4600 1938.0400 1020.9400 ;
        RECT 1920.9000 1009.5800 1922.5000 1010.0600 ;
        RECT 1920.9000 1015.0200 1922.5000 1015.5000 ;
        RECT 1920.9000 1020.4600 1922.5000 1020.9400 ;
        RECT 1936.4400 998.7000 1938.0400 999.1800 ;
        RECT 1936.4400 1004.1400 1938.0400 1004.6200 ;
        RECT 1920.9000 998.7000 1922.5000 999.1800 ;
        RECT 1920.9000 1004.1400 1922.5000 1004.6200 ;
        RECT 1936.4400 982.3800 1938.0400 982.8600 ;
        RECT 1936.4400 987.8200 1938.0400 988.3000 ;
        RECT 1936.4400 993.2600 1938.0400 993.7400 ;
        RECT 1920.9000 982.3800 1922.5000 982.8600 ;
        RECT 1920.9000 987.8200 1922.5000 988.3000 ;
        RECT 1920.9000 993.2600 1922.5000 993.7400 ;
        RECT 1875.9000 1025.9000 1877.5000 1026.3800 ;
        RECT 1875.9000 1031.3400 1877.5000 1031.8200 ;
        RECT 1875.9000 1009.5800 1877.5000 1010.0600 ;
        RECT 1875.9000 1015.0200 1877.5000 1015.5000 ;
        RECT 1875.9000 1020.4600 1877.5000 1020.9400 ;
        RECT 1875.9000 998.7000 1877.5000 999.1800 ;
        RECT 1875.9000 1004.1400 1877.5000 1004.6200 ;
        RECT 1875.9000 982.3800 1877.5000 982.8600 ;
        RECT 1875.9000 987.8200 1877.5000 988.3000 ;
        RECT 1875.9000 993.2600 1877.5000 993.7400 ;
        RECT 1875.9000 1036.7800 1877.5000 1037.2600 ;
        RECT 1920.9000 1036.7800 1922.5000 1037.2600 ;
        RECT 1936.4400 1036.7800 1938.0400 1037.2600 ;
        RECT 1830.9000 1069.4200 1832.5000 1069.9000 ;
        RECT 1830.9000 1074.8600 1832.5000 1075.3400 ;
        RECT 1830.9000 1080.3000 1832.5000 1080.7800 ;
        RECT 1785.9000 1069.4200 1787.5000 1069.9000 ;
        RECT 1785.9000 1074.8600 1787.5000 1075.3400 ;
        RECT 1785.9000 1080.3000 1787.5000 1080.7800 ;
        RECT 1830.9000 1053.1000 1832.5000 1053.5800 ;
        RECT 1830.9000 1058.5400 1832.5000 1059.0200 ;
        RECT 1830.9000 1042.2200 1832.5000 1042.7000 ;
        RECT 1830.9000 1047.6600 1832.5000 1048.1400 ;
        RECT 1785.9000 1053.1000 1787.5000 1053.5800 ;
        RECT 1785.9000 1058.5400 1787.5000 1059.0200 ;
        RECT 1785.9000 1042.2200 1787.5000 1042.7000 ;
        RECT 1785.9000 1047.6600 1787.5000 1048.1400 ;
        RECT 1785.9000 1063.9800 1787.5000 1064.4600 ;
        RECT 1830.9000 1063.9800 1832.5000 1064.4600 ;
        RECT 1733.7400 1080.3000 1735.3400 1080.7800 ;
        RECT 1740.9000 1080.3000 1742.5000 1080.7800 ;
        RECT 1740.9000 1069.4200 1742.5000 1069.9000 ;
        RECT 1740.9000 1074.8600 1742.5000 1075.3400 ;
        RECT 1733.7400 1069.4200 1735.3400 1069.9000 ;
        RECT 1733.7400 1074.8600 1735.3400 1075.3400 ;
        RECT 1740.9000 1053.1000 1742.5000 1053.5800 ;
        RECT 1740.9000 1058.5400 1742.5000 1059.0200 ;
        RECT 1733.7400 1053.1000 1735.3400 1053.5800 ;
        RECT 1733.7400 1058.5400 1735.3400 1059.0200 ;
        RECT 1740.9000 1042.2200 1742.5000 1042.7000 ;
        RECT 1740.9000 1047.6600 1742.5000 1048.1400 ;
        RECT 1733.7400 1042.2200 1735.3400 1042.7000 ;
        RECT 1733.7400 1047.6600 1735.3400 1048.1400 ;
        RECT 1733.7400 1063.9800 1735.3400 1064.4600 ;
        RECT 1740.9000 1063.9800 1742.5000 1064.4600 ;
        RECT 1830.9000 1025.9000 1832.5000 1026.3800 ;
        RECT 1830.9000 1031.3400 1832.5000 1031.8200 ;
        RECT 1830.9000 1009.5800 1832.5000 1010.0600 ;
        RECT 1830.9000 1015.0200 1832.5000 1015.5000 ;
        RECT 1830.9000 1020.4600 1832.5000 1020.9400 ;
        RECT 1785.9000 1025.9000 1787.5000 1026.3800 ;
        RECT 1785.9000 1031.3400 1787.5000 1031.8200 ;
        RECT 1785.9000 1009.5800 1787.5000 1010.0600 ;
        RECT 1785.9000 1015.0200 1787.5000 1015.5000 ;
        RECT 1785.9000 1020.4600 1787.5000 1020.9400 ;
        RECT 1830.9000 998.7000 1832.5000 999.1800 ;
        RECT 1830.9000 1004.1400 1832.5000 1004.6200 ;
        RECT 1830.9000 982.3800 1832.5000 982.8600 ;
        RECT 1830.9000 987.8200 1832.5000 988.3000 ;
        RECT 1830.9000 993.2600 1832.5000 993.7400 ;
        RECT 1785.9000 998.7000 1787.5000 999.1800 ;
        RECT 1785.9000 1004.1400 1787.5000 1004.6200 ;
        RECT 1785.9000 982.3800 1787.5000 982.8600 ;
        RECT 1785.9000 987.8200 1787.5000 988.3000 ;
        RECT 1785.9000 993.2600 1787.5000 993.7400 ;
        RECT 1740.9000 1025.9000 1742.5000 1026.3800 ;
        RECT 1740.9000 1031.3400 1742.5000 1031.8200 ;
        RECT 1733.7400 1025.9000 1735.3400 1026.3800 ;
        RECT 1733.7400 1031.3400 1735.3400 1031.8200 ;
        RECT 1740.9000 1009.5800 1742.5000 1010.0600 ;
        RECT 1740.9000 1015.0200 1742.5000 1015.5000 ;
        RECT 1740.9000 1020.4600 1742.5000 1020.9400 ;
        RECT 1733.7400 1009.5800 1735.3400 1010.0600 ;
        RECT 1733.7400 1015.0200 1735.3400 1015.5000 ;
        RECT 1733.7400 1020.4600 1735.3400 1020.9400 ;
        RECT 1740.9000 998.7000 1742.5000 999.1800 ;
        RECT 1740.9000 1004.1400 1742.5000 1004.6200 ;
        RECT 1733.7400 998.7000 1735.3400 999.1800 ;
        RECT 1733.7400 1004.1400 1735.3400 1004.6200 ;
        RECT 1740.9000 982.3800 1742.5000 982.8600 ;
        RECT 1740.9000 987.8200 1742.5000 988.3000 ;
        RECT 1740.9000 993.2600 1742.5000 993.7400 ;
        RECT 1733.7400 982.3800 1735.3400 982.8600 ;
        RECT 1733.7400 987.8200 1735.3400 988.3000 ;
        RECT 1733.7400 993.2600 1735.3400 993.7400 ;
        RECT 1733.7400 1036.7800 1735.3400 1037.2600 ;
        RECT 1740.9000 1036.7800 1742.5000 1037.2600 ;
        RECT 1785.9000 1036.7800 1787.5000 1037.2600 ;
        RECT 1830.9000 1036.7800 1832.5000 1037.2600 ;
        RECT 1936.4400 971.5000 1938.0400 971.9800 ;
        RECT 1936.4400 976.9400 1938.0400 977.4200 ;
        RECT 1920.9000 971.5000 1922.5000 971.9800 ;
        RECT 1920.9000 976.9400 1922.5000 977.4200 ;
        RECT 1936.4400 955.1800 1938.0400 955.6600 ;
        RECT 1936.4400 960.6200 1938.0400 961.1000 ;
        RECT 1936.4400 966.0600 1938.0400 966.5400 ;
        RECT 1920.9000 955.1800 1922.5000 955.6600 ;
        RECT 1920.9000 960.6200 1922.5000 961.1000 ;
        RECT 1920.9000 966.0600 1922.5000 966.5400 ;
        RECT 1936.4400 944.3000 1938.0400 944.7800 ;
        RECT 1936.4400 949.7400 1938.0400 950.2200 ;
        RECT 1920.9000 944.3000 1922.5000 944.7800 ;
        RECT 1920.9000 949.7400 1922.5000 950.2200 ;
        RECT 1936.4400 927.9800 1938.0400 928.4600 ;
        RECT 1936.4400 933.4200 1938.0400 933.9000 ;
        RECT 1936.4400 938.8600 1938.0400 939.3400 ;
        RECT 1920.9000 927.9800 1922.5000 928.4600 ;
        RECT 1920.9000 933.4200 1922.5000 933.9000 ;
        RECT 1920.9000 938.8600 1922.5000 939.3400 ;
        RECT 1875.9000 971.5000 1877.5000 971.9800 ;
        RECT 1875.9000 976.9400 1877.5000 977.4200 ;
        RECT 1875.9000 955.1800 1877.5000 955.6600 ;
        RECT 1875.9000 960.6200 1877.5000 961.1000 ;
        RECT 1875.9000 966.0600 1877.5000 966.5400 ;
        RECT 1875.9000 944.3000 1877.5000 944.7800 ;
        RECT 1875.9000 949.7400 1877.5000 950.2200 ;
        RECT 1875.9000 927.9800 1877.5000 928.4600 ;
        RECT 1875.9000 933.4200 1877.5000 933.9000 ;
        RECT 1875.9000 938.8600 1877.5000 939.3400 ;
        RECT 1936.4400 917.1000 1938.0400 917.5800 ;
        RECT 1936.4400 922.5400 1938.0400 923.0200 ;
        RECT 1920.9000 917.1000 1922.5000 917.5800 ;
        RECT 1920.9000 922.5400 1922.5000 923.0200 ;
        RECT 1936.4400 900.7800 1938.0400 901.2600 ;
        RECT 1936.4400 906.2200 1938.0400 906.7000 ;
        RECT 1936.4400 911.6600 1938.0400 912.1400 ;
        RECT 1920.9000 900.7800 1922.5000 901.2600 ;
        RECT 1920.9000 906.2200 1922.5000 906.7000 ;
        RECT 1920.9000 911.6600 1922.5000 912.1400 ;
        RECT 1936.4400 889.9000 1938.0400 890.3800 ;
        RECT 1936.4400 895.3400 1938.0400 895.8200 ;
        RECT 1920.9000 889.9000 1922.5000 890.3800 ;
        RECT 1920.9000 895.3400 1922.5000 895.8200 ;
        RECT 1920.9000 884.4600 1922.5000 884.9400 ;
        RECT 1936.4400 884.4600 1938.0400 884.9400 ;
        RECT 1875.9000 917.1000 1877.5000 917.5800 ;
        RECT 1875.9000 922.5400 1877.5000 923.0200 ;
        RECT 1875.9000 900.7800 1877.5000 901.2600 ;
        RECT 1875.9000 906.2200 1877.5000 906.7000 ;
        RECT 1875.9000 911.6600 1877.5000 912.1400 ;
        RECT 1875.9000 889.9000 1877.5000 890.3800 ;
        RECT 1875.9000 895.3400 1877.5000 895.8200 ;
        RECT 1875.9000 884.4600 1877.5000 884.9400 ;
        RECT 1830.9000 971.5000 1832.5000 971.9800 ;
        RECT 1830.9000 976.9400 1832.5000 977.4200 ;
        RECT 1830.9000 955.1800 1832.5000 955.6600 ;
        RECT 1830.9000 960.6200 1832.5000 961.1000 ;
        RECT 1830.9000 966.0600 1832.5000 966.5400 ;
        RECT 1785.9000 971.5000 1787.5000 971.9800 ;
        RECT 1785.9000 976.9400 1787.5000 977.4200 ;
        RECT 1785.9000 955.1800 1787.5000 955.6600 ;
        RECT 1785.9000 960.6200 1787.5000 961.1000 ;
        RECT 1785.9000 966.0600 1787.5000 966.5400 ;
        RECT 1830.9000 944.3000 1832.5000 944.7800 ;
        RECT 1830.9000 949.7400 1832.5000 950.2200 ;
        RECT 1830.9000 927.9800 1832.5000 928.4600 ;
        RECT 1830.9000 933.4200 1832.5000 933.9000 ;
        RECT 1830.9000 938.8600 1832.5000 939.3400 ;
        RECT 1785.9000 944.3000 1787.5000 944.7800 ;
        RECT 1785.9000 949.7400 1787.5000 950.2200 ;
        RECT 1785.9000 927.9800 1787.5000 928.4600 ;
        RECT 1785.9000 933.4200 1787.5000 933.9000 ;
        RECT 1785.9000 938.8600 1787.5000 939.3400 ;
        RECT 1740.9000 971.5000 1742.5000 971.9800 ;
        RECT 1740.9000 976.9400 1742.5000 977.4200 ;
        RECT 1733.7400 971.5000 1735.3400 971.9800 ;
        RECT 1733.7400 976.9400 1735.3400 977.4200 ;
        RECT 1740.9000 955.1800 1742.5000 955.6600 ;
        RECT 1740.9000 960.6200 1742.5000 961.1000 ;
        RECT 1740.9000 966.0600 1742.5000 966.5400 ;
        RECT 1733.7400 955.1800 1735.3400 955.6600 ;
        RECT 1733.7400 960.6200 1735.3400 961.1000 ;
        RECT 1733.7400 966.0600 1735.3400 966.5400 ;
        RECT 1740.9000 944.3000 1742.5000 944.7800 ;
        RECT 1740.9000 949.7400 1742.5000 950.2200 ;
        RECT 1733.7400 944.3000 1735.3400 944.7800 ;
        RECT 1733.7400 949.7400 1735.3400 950.2200 ;
        RECT 1740.9000 927.9800 1742.5000 928.4600 ;
        RECT 1740.9000 933.4200 1742.5000 933.9000 ;
        RECT 1740.9000 938.8600 1742.5000 939.3400 ;
        RECT 1733.7400 927.9800 1735.3400 928.4600 ;
        RECT 1733.7400 933.4200 1735.3400 933.9000 ;
        RECT 1733.7400 938.8600 1735.3400 939.3400 ;
        RECT 1830.9000 917.1000 1832.5000 917.5800 ;
        RECT 1830.9000 922.5400 1832.5000 923.0200 ;
        RECT 1830.9000 900.7800 1832.5000 901.2600 ;
        RECT 1830.9000 906.2200 1832.5000 906.7000 ;
        RECT 1830.9000 911.6600 1832.5000 912.1400 ;
        RECT 1785.9000 917.1000 1787.5000 917.5800 ;
        RECT 1785.9000 922.5400 1787.5000 923.0200 ;
        RECT 1785.9000 900.7800 1787.5000 901.2600 ;
        RECT 1785.9000 906.2200 1787.5000 906.7000 ;
        RECT 1785.9000 911.6600 1787.5000 912.1400 ;
        RECT 1830.9000 895.3400 1832.5000 895.8200 ;
        RECT 1830.9000 889.9000 1832.5000 890.3800 ;
        RECT 1830.9000 884.4600 1832.5000 884.9400 ;
        RECT 1785.9000 895.3400 1787.5000 895.8200 ;
        RECT 1785.9000 889.9000 1787.5000 890.3800 ;
        RECT 1785.9000 884.4600 1787.5000 884.9400 ;
        RECT 1740.9000 917.1000 1742.5000 917.5800 ;
        RECT 1740.9000 922.5400 1742.5000 923.0200 ;
        RECT 1733.7400 917.1000 1735.3400 917.5800 ;
        RECT 1733.7400 922.5400 1735.3400 923.0200 ;
        RECT 1740.9000 900.7800 1742.5000 901.2600 ;
        RECT 1740.9000 906.2200 1742.5000 906.7000 ;
        RECT 1740.9000 911.6600 1742.5000 912.1400 ;
        RECT 1733.7400 900.7800 1735.3400 901.2600 ;
        RECT 1733.7400 906.2200 1735.3400 906.7000 ;
        RECT 1733.7400 911.6600 1735.3400 912.1400 ;
        RECT 1740.9000 889.9000 1742.5000 890.3800 ;
        RECT 1740.9000 895.3400 1742.5000 895.8200 ;
        RECT 1733.7400 889.9000 1735.3400 890.3800 ;
        RECT 1733.7400 895.3400 1735.3400 895.8200 ;
        RECT 1733.7400 884.4600 1735.3400 884.9400 ;
        RECT 1740.9000 884.4600 1742.5000 884.9400 ;
        RECT 1730.7800 1086.6500 1941.0000 1088.2500 ;
        RECT 1730.7800 874.9500 1941.0000 876.5500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 872.1200 1735.3400 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 1090.1600 1735.3400 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 872.1200 1938.0400 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 1090.1600 1938.0400 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 874.9500 1732.3800 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 874.9500 1941.0000 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1086.6500 1732.3800 1088.2500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1086.6500 1941.0000 1088.2500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 645.3100 1922.5000 858.6100 ;
        RECT 1875.9000 645.3100 1877.5000 858.6100 ;
        RECT 1830.9000 645.3100 1832.5000 858.6100 ;
        RECT 1785.9000 645.3100 1787.5000 858.6100 ;
        RECT 1740.9000 645.3100 1742.5000 858.6100 ;
        RECT 1936.4400 642.4800 1938.0400 862.1200 ;
        RECT 1733.7400 642.4800 1735.3400 862.1200 ;
      LAYER met3 ;
        RECT 1920.9000 850.6600 1922.5000 851.1400 ;
        RECT 1936.4400 850.6600 1938.0400 851.1400 ;
        RECT 1936.4400 839.7800 1938.0400 840.2600 ;
        RECT 1936.4400 845.2200 1938.0400 845.7000 ;
        RECT 1920.9000 839.7800 1922.5000 840.2600 ;
        RECT 1920.9000 845.2200 1922.5000 845.7000 ;
        RECT 1936.4400 823.4600 1938.0400 823.9400 ;
        RECT 1936.4400 828.9000 1938.0400 829.3800 ;
        RECT 1920.9000 823.4600 1922.5000 823.9400 ;
        RECT 1920.9000 828.9000 1922.5000 829.3800 ;
        RECT 1936.4400 812.5800 1938.0400 813.0600 ;
        RECT 1936.4400 818.0200 1938.0400 818.5000 ;
        RECT 1920.9000 812.5800 1922.5000 813.0600 ;
        RECT 1920.9000 818.0200 1922.5000 818.5000 ;
        RECT 1920.9000 834.3400 1922.5000 834.8200 ;
        RECT 1936.4400 834.3400 1938.0400 834.8200 ;
        RECT 1875.9000 839.7800 1877.5000 840.2600 ;
        RECT 1875.9000 845.2200 1877.5000 845.7000 ;
        RECT 1875.9000 850.6600 1877.5000 851.1400 ;
        RECT 1875.9000 823.4600 1877.5000 823.9400 ;
        RECT 1875.9000 828.9000 1877.5000 829.3800 ;
        RECT 1875.9000 818.0200 1877.5000 818.5000 ;
        RECT 1875.9000 812.5800 1877.5000 813.0600 ;
        RECT 1875.9000 834.3400 1877.5000 834.8200 ;
        RECT 1936.4400 796.2600 1938.0400 796.7400 ;
        RECT 1936.4400 801.7000 1938.0400 802.1800 ;
        RECT 1920.9000 796.2600 1922.5000 796.7400 ;
        RECT 1920.9000 801.7000 1922.5000 802.1800 ;
        RECT 1936.4400 779.9400 1938.0400 780.4200 ;
        RECT 1936.4400 785.3800 1938.0400 785.8600 ;
        RECT 1936.4400 790.8200 1938.0400 791.3000 ;
        RECT 1920.9000 779.9400 1922.5000 780.4200 ;
        RECT 1920.9000 785.3800 1922.5000 785.8600 ;
        RECT 1920.9000 790.8200 1922.5000 791.3000 ;
        RECT 1936.4400 769.0600 1938.0400 769.5400 ;
        RECT 1936.4400 774.5000 1938.0400 774.9800 ;
        RECT 1920.9000 769.0600 1922.5000 769.5400 ;
        RECT 1920.9000 774.5000 1922.5000 774.9800 ;
        RECT 1936.4400 752.7400 1938.0400 753.2200 ;
        RECT 1936.4400 758.1800 1938.0400 758.6600 ;
        RECT 1936.4400 763.6200 1938.0400 764.1000 ;
        RECT 1920.9000 752.7400 1922.5000 753.2200 ;
        RECT 1920.9000 758.1800 1922.5000 758.6600 ;
        RECT 1920.9000 763.6200 1922.5000 764.1000 ;
        RECT 1875.9000 796.2600 1877.5000 796.7400 ;
        RECT 1875.9000 801.7000 1877.5000 802.1800 ;
        RECT 1875.9000 779.9400 1877.5000 780.4200 ;
        RECT 1875.9000 785.3800 1877.5000 785.8600 ;
        RECT 1875.9000 790.8200 1877.5000 791.3000 ;
        RECT 1875.9000 769.0600 1877.5000 769.5400 ;
        RECT 1875.9000 774.5000 1877.5000 774.9800 ;
        RECT 1875.9000 752.7400 1877.5000 753.2200 ;
        RECT 1875.9000 758.1800 1877.5000 758.6600 ;
        RECT 1875.9000 763.6200 1877.5000 764.1000 ;
        RECT 1875.9000 807.1400 1877.5000 807.6200 ;
        RECT 1920.9000 807.1400 1922.5000 807.6200 ;
        RECT 1936.4400 807.1400 1938.0400 807.6200 ;
        RECT 1830.9000 839.7800 1832.5000 840.2600 ;
        RECT 1830.9000 845.2200 1832.5000 845.7000 ;
        RECT 1830.9000 850.6600 1832.5000 851.1400 ;
        RECT 1785.9000 839.7800 1787.5000 840.2600 ;
        RECT 1785.9000 845.2200 1787.5000 845.7000 ;
        RECT 1785.9000 850.6600 1787.5000 851.1400 ;
        RECT 1830.9000 823.4600 1832.5000 823.9400 ;
        RECT 1830.9000 828.9000 1832.5000 829.3800 ;
        RECT 1830.9000 812.5800 1832.5000 813.0600 ;
        RECT 1830.9000 818.0200 1832.5000 818.5000 ;
        RECT 1785.9000 823.4600 1787.5000 823.9400 ;
        RECT 1785.9000 828.9000 1787.5000 829.3800 ;
        RECT 1785.9000 812.5800 1787.5000 813.0600 ;
        RECT 1785.9000 818.0200 1787.5000 818.5000 ;
        RECT 1785.9000 834.3400 1787.5000 834.8200 ;
        RECT 1830.9000 834.3400 1832.5000 834.8200 ;
        RECT 1733.7400 850.6600 1735.3400 851.1400 ;
        RECT 1740.9000 850.6600 1742.5000 851.1400 ;
        RECT 1740.9000 839.7800 1742.5000 840.2600 ;
        RECT 1740.9000 845.2200 1742.5000 845.7000 ;
        RECT 1733.7400 839.7800 1735.3400 840.2600 ;
        RECT 1733.7400 845.2200 1735.3400 845.7000 ;
        RECT 1740.9000 823.4600 1742.5000 823.9400 ;
        RECT 1740.9000 828.9000 1742.5000 829.3800 ;
        RECT 1733.7400 823.4600 1735.3400 823.9400 ;
        RECT 1733.7400 828.9000 1735.3400 829.3800 ;
        RECT 1740.9000 812.5800 1742.5000 813.0600 ;
        RECT 1740.9000 818.0200 1742.5000 818.5000 ;
        RECT 1733.7400 812.5800 1735.3400 813.0600 ;
        RECT 1733.7400 818.0200 1735.3400 818.5000 ;
        RECT 1733.7400 834.3400 1735.3400 834.8200 ;
        RECT 1740.9000 834.3400 1742.5000 834.8200 ;
        RECT 1830.9000 796.2600 1832.5000 796.7400 ;
        RECT 1830.9000 801.7000 1832.5000 802.1800 ;
        RECT 1830.9000 779.9400 1832.5000 780.4200 ;
        RECT 1830.9000 785.3800 1832.5000 785.8600 ;
        RECT 1830.9000 790.8200 1832.5000 791.3000 ;
        RECT 1785.9000 796.2600 1787.5000 796.7400 ;
        RECT 1785.9000 801.7000 1787.5000 802.1800 ;
        RECT 1785.9000 779.9400 1787.5000 780.4200 ;
        RECT 1785.9000 785.3800 1787.5000 785.8600 ;
        RECT 1785.9000 790.8200 1787.5000 791.3000 ;
        RECT 1830.9000 769.0600 1832.5000 769.5400 ;
        RECT 1830.9000 774.5000 1832.5000 774.9800 ;
        RECT 1830.9000 752.7400 1832.5000 753.2200 ;
        RECT 1830.9000 758.1800 1832.5000 758.6600 ;
        RECT 1830.9000 763.6200 1832.5000 764.1000 ;
        RECT 1785.9000 769.0600 1787.5000 769.5400 ;
        RECT 1785.9000 774.5000 1787.5000 774.9800 ;
        RECT 1785.9000 752.7400 1787.5000 753.2200 ;
        RECT 1785.9000 758.1800 1787.5000 758.6600 ;
        RECT 1785.9000 763.6200 1787.5000 764.1000 ;
        RECT 1740.9000 796.2600 1742.5000 796.7400 ;
        RECT 1740.9000 801.7000 1742.5000 802.1800 ;
        RECT 1733.7400 796.2600 1735.3400 796.7400 ;
        RECT 1733.7400 801.7000 1735.3400 802.1800 ;
        RECT 1740.9000 779.9400 1742.5000 780.4200 ;
        RECT 1740.9000 785.3800 1742.5000 785.8600 ;
        RECT 1740.9000 790.8200 1742.5000 791.3000 ;
        RECT 1733.7400 779.9400 1735.3400 780.4200 ;
        RECT 1733.7400 785.3800 1735.3400 785.8600 ;
        RECT 1733.7400 790.8200 1735.3400 791.3000 ;
        RECT 1740.9000 769.0600 1742.5000 769.5400 ;
        RECT 1740.9000 774.5000 1742.5000 774.9800 ;
        RECT 1733.7400 769.0600 1735.3400 769.5400 ;
        RECT 1733.7400 774.5000 1735.3400 774.9800 ;
        RECT 1740.9000 752.7400 1742.5000 753.2200 ;
        RECT 1740.9000 758.1800 1742.5000 758.6600 ;
        RECT 1740.9000 763.6200 1742.5000 764.1000 ;
        RECT 1733.7400 752.7400 1735.3400 753.2200 ;
        RECT 1733.7400 758.1800 1735.3400 758.6600 ;
        RECT 1733.7400 763.6200 1735.3400 764.1000 ;
        RECT 1733.7400 807.1400 1735.3400 807.6200 ;
        RECT 1740.9000 807.1400 1742.5000 807.6200 ;
        RECT 1785.9000 807.1400 1787.5000 807.6200 ;
        RECT 1830.9000 807.1400 1832.5000 807.6200 ;
        RECT 1936.4400 741.8600 1938.0400 742.3400 ;
        RECT 1936.4400 747.3000 1938.0400 747.7800 ;
        RECT 1920.9000 741.8600 1922.5000 742.3400 ;
        RECT 1920.9000 747.3000 1922.5000 747.7800 ;
        RECT 1936.4400 725.5400 1938.0400 726.0200 ;
        RECT 1936.4400 730.9800 1938.0400 731.4600 ;
        RECT 1936.4400 736.4200 1938.0400 736.9000 ;
        RECT 1920.9000 725.5400 1922.5000 726.0200 ;
        RECT 1920.9000 730.9800 1922.5000 731.4600 ;
        RECT 1920.9000 736.4200 1922.5000 736.9000 ;
        RECT 1936.4400 714.6600 1938.0400 715.1400 ;
        RECT 1936.4400 720.1000 1938.0400 720.5800 ;
        RECT 1920.9000 714.6600 1922.5000 715.1400 ;
        RECT 1920.9000 720.1000 1922.5000 720.5800 ;
        RECT 1936.4400 698.3400 1938.0400 698.8200 ;
        RECT 1936.4400 703.7800 1938.0400 704.2600 ;
        RECT 1936.4400 709.2200 1938.0400 709.7000 ;
        RECT 1920.9000 698.3400 1922.5000 698.8200 ;
        RECT 1920.9000 703.7800 1922.5000 704.2600 ;
        RECT 1920.9000 709.2200 1922.5000 709.7000 ;
        RECT 1875.9000 741.8600 1877.5000 742.3400 ;
        RECT 1875.9000 747.3000 1877.5000 747.7800 ;
        RECT 1875.9000 725.5400 1877.5000 726.0200 ;
        RECT 1875.9000 730.9800 1877.5000 731.4600 ;
        RECT 1875.9000 736.4200 1877.5000 736.9000 ;
        RECT 1875.9000 714.6600 1877.5000 715.1400 ;
        RECT 1875.9000 720.1000 1877.5000 720.5800 ;
        RECT 1875.9000 698.3400 1877.5000 698.8200 ;
        RECT 1875.9000 703.7800 1877.5000 704.2600 ;
        RECT 1875.9000 709.2200 1877.5000 709.7000 ;
        RECT 1936.4400 687.4600 1938.0400 687.9400 ;
        RECT 1936.4400 692.9000 1938.0400 693.3800 ;
        RECT 1920.9000 687.4600 1922.5000 687.9400 ;
        RECT 1920.9000 692.9000 1922.5000 693.3800 ;
        RECT 1936.4400 671.1400 1938.0400 671.6200 ;
        RECT 1936.4400 676.5800 1938.0400 677.0600 ;
        RECT 1936.4400 682.0200 1938.0400 682.5000 ;
        RECT 1920.9000 671.1400 1922.5000 671.6200 ;
        RECT 1920.9000 676.5800 1922.5000 677.0600 ;
        RECT 1920.9000 682.0200 1922.5000 682.5000 ;
        RECT 1936.4400 660.2600 1938.0400 660.7400 ;
        RECT 1936.4400 665.7000 1938.0400 666.1800 ;
        RECT 1920.9000 660.2600 1922.5000 660.7400 ;
        RECT 1920.9000 665.7000 1922.5000 666.1800 ;
        RECT 1920.9000 654.8200 1922.5000 655.3000 ;
        RECT 1936.4400 654.8200 1938.0400 655.3000 ;
        RECT 1875.9000 687.4600 1877.5000 687.9400 ;
        RECT 1875.9000 692.9000 1877.5000 693.3800 ;
        RECT 1875.9000 671.1400 1877.5000 671.6200 ;
        RECT 1875.9000 676.5800 1877.5000 677.0600 ;
        RECT 1875.9000 682.0200 1877.5000 682.5000 ;
        RECT 1875.9000 660.2600 1877.5000 660.7400 ;
        RECT 1875.9000 665.7000 1877.5000 666.1800 ;
        RECT 1875.9000 654.8200 1877.5000 655.3000 ;
        RECT 1830.9000 741.8600 1832.5000 742.3400 ;
        RECT 1830.9000 747.3000 1832.5000 747.7800 ;
        RECT 1830.9000 725.5400 1832.5000 726.0200 ;
        RECT 1830.9000 730.9800 1832.5000 731.4600 ;
        RECT 1830.9000 736.4200 1832.5000 736.9000 ;
        RECT 1785.9000 741.8600 1787.5000 742.3400 ;
        RECT 1785.9000 747.3000 1787.5000 747.7800 ;
        RECT 1785.9000 725.5400 1787.5000 726.0200 ;
        RECT 1785.9000 730.9800 1787.5000 731.4600 ;
        RECT 1785.9000 736.4200 1787.5000 736.9000 ;
        RECT 1830.9000 714.6600 1832.5000 715.1400 ;
        RECT 1830.9000 720.1000 1832.5000 720.5800 ;
        RECT 1830.9000 698.3400 1832.5000 698.8200 ;
        RECT 1830.9000 703.7800 1832.5000 704.2600 ;
        RECT 1830.9000 709.2200 1832.5000 709.7000 ;
        RECT 1785.9000 714.6600 1787.5000 715.1400 ;
        RECT 1785.9000 720.1000 1787.5000 720.5800 ;
        RECT 1785.9000 698.3400 1787.5000 698.8200 ;
        RECT 1785.9000 703.7800 1787.5000 704.2600 ;
        RECT 1785.9000 709.2200 1787.5000 709.7000 ;
        RECT 1740.9000 741.8600 1742.5000 742.3400 ;
        RECT 1740.9000 747.3000 1742.5000 747.7800 ;
        RECT 1733.7400 741.8600 1735.3400 742.3400 ;
        RECT 1733.7400 747.3000 1735.3400 747.7800 ;
        RECT 1740.9000 725.5400 1742.5000 726.0200 ;
        RECT 1740.9000 730.9800 1742.5000 731.4600 ;
        RECT 1740.9000 736.4200 1742.5000 736.9000 ;
        RECT 1733.7400 725.5400 1735.3400 726.0200 ;
        RECT 1733.7400 730.9800 1735.3400 731.4600 ;
        RECT 1733.7400 736.4200 1735.3400 736.9000 ;
        RECT 1740.9000 714.6600 1742.5000 715.1400 ;
        RECT 1740.9000 720.1000 1742.5000 720.5800 ;
        RECT 1733.7400 714.6600 1735.3400 715.1400 ;
        RECT 1733.7400 720.1000 1735.3400 720.5800 ;
        RECT 1740.9000 698.3400 1742.5000 698.8200 ;
        RECT 1740.9000 703.7800 1742.5000 704.2600 ;
        RECT 1740.9000 709.2200 1742.5000 709.7000 ;
        RECT 1733.7400 698.3400 1735.3400 698.8200 ;
        RECT 1733.7400 703.7800 1735.3400 704.2600 ;
        RECT 1733.7400 709.2200 1735.3400 709.7000 ;
        RECT 1830.9000 687.4600 1832.5000 687.9400 ;
        RECT 1830.9000 692.9000 1832.5000 693.3800 ;
        RECT 1830.9000 671.1400 1832.5000 671.6200 ;
        RECT 1830.9000 676.5800 1832.5000 677.0600 ;
        RECT 1830.9000 682.0200 1832.5000 682.5000 ;
        RECT 1785.9000 687.4600 1787.5000 687.9400 ;
        RECT 1785.9000 692.9000 1787.5000 693.3800 ;
        RECT 1785.9000 671.1400 1787.5000 671.6200 ;
        RECT 1785.9000 676.5800 1787.5000 677.0600 ;
        RECT 1785.9000 682.0200 1787.5000 682.5000 ;
        RECT 1830.9000 665.7000 1832.5000 666.1800 ;
        RECT 1830.9000 660.2600 1832.5000 660.7400 ;
        RECT 1830.9000 654.8200 1832.5000 655.3000 ;
        RECT 1785.9000 665.7000 1787.5000 666.1800 ;
        RECT 1785.9000 660.2600 1787.5000 660.7400 ;
        RECT 1785.9000 654.8200 1787.5000 655.3000 ;
        RECT 1740.9000 687.4600 1742.5000 687.9400 ;
        RECT 1740.9000 692.9000 1742.5000 693.3800 ;
        RECT 1733.7400 687.4600 1735.3400 687.9400 ;
        RECT 1733.7400 692.9000 1735.3400 693.3800 ;
        RECT 1740.9000 671.1400 1742.5000 671.6200 ;
        RECT 1740.9000 676.5800 1742.5000 677.0600 ;
        RECT 1740.9000 682.0200 1742.5000 682.5000 ;
        RECT 1733.7400 671.1400 1735.3400 671.6200 ;
        RECT 1733.7400 676.5800 1735.3400 677.0600 ;
        RECT 1733.7400 682.0200 1735.3400 682.5000 ;
        RECT 1740.9000 660.2600 1742.5000 660.7400 ;
        RECT 1740.9000 665.7000 1742.5000 666.1800 ;
        RECT 1733.7400 660.2600 1735.3400 660.7400 ;
        RECT 1733.7400 665.7000 1735.3400 666.1800 ;
        RECT 1733.7400 654.8200 1735.3400 655.3000 ;
        RECT 1740.9000 654.8200 1742.5000 655.3000 ;
        RECT 1730.7800 857.0100 1941.0000 858.6100 ;
        RECT 1730.7800 645.3100 1941.0000 646.9100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 642.4800 1735.3400 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 860.5200 1735.3400 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 642.4800 1938.0400 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 860.5200 1938.0400 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 645.3100 1732.3800 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 645.3100 1941.0000 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 857.0100 1732.3800 858.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 857.0100 1941.0000 858.6100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1920.9000 415.6700 1922.5000 628.9700 ;
        RECT 1875.9000 415.6700 1877.5000 628.9700 ;
        RECT 1830.9000 415.6700 1832.5000 628.9700 ;
        RECT 1785.9000 415.6700 1787.5000 628.9700 ;
        RECT 1740.9000 415.6700 1742.5000 628.9700 ;
        RECT 1936.4400 412.8400 1938.0400 632.4800 ;
        RECT 1733.7400 412.8400 1735.3400 632.4800 ;
      LAYER met3 ;
        RECT 1920.9000 621.0200 1922.5000 621.5000 ;
        RECT 1936.4400 621.0200 1938.0400 621.5000 ;
        RECT 1936.4400 610.1400 1938.0400 610.6200 ;
        RECT 1936.4400 615.5800 1938.0400 616.0600 ;
        RECT 1920.9000 610.1400 1922.5000 610.6200 ;
        RECT 1920.9000 615.5800 1922.5000 616.0600 ;
        RECT 1936.4400 593.8200 1938.0400 594.3000 ;
        RECT 1936.4400 599.2600 1938.0400 599.7400 ;
        RECT 1920.9000 593.8200 1922.5000 594.3000 ;
        RECT 1920.9000 599.2600 1922.5000 599.7400 ;
        RECT 1936.4400 582.9400 1938.0400 583.4200 ;
        RECT 1936.4400 588.3800 1938.0400 588.8600 ;
        RECT 1920.9000 582.9400 1922.5000 583.4200 ;
        RECT 1920.9000 588.3800 1922.5000 588.8600 ;
        RECT 1920.9000 604.7000 1922.5000 605.1800 ;
        RECT 1936.4400 604.7000 1938.0400 605.1800 ;
        RECT 1875.9000 610.1400 1877.5000 610.6200 ;
        RECT 1875.9000 615.5800 1877.5000 616.0600 ;
        RECT 1875.9000 621.0200 1877.5000 621.5000 ;
        RECT 1875.9000 593.8200 1877.5000 594.3000 ;
        RECT 1875.9000 599.2600 1877.5000 599.7400 ;
        RECT 1875.9000 588.3800 1877.5000 588.8600 ;
        RECT 1875.9000 582.9400 1877.5000 583.4200 ;
        RECT 1875.9000 604.7000 1877.5000 605.1800 ;
        RECT 1936.4400 566.6200 1938.0400 567.1000 ;
        RECT 1936.4400 572.0600 1938.0400 572.5400 ;
        RECT 1920.9000 566.6200 1922.5000 567.1000 ;
        RECT 1920.9000 572.0600 1922.5000 572.5400 ;
        RECT 1936.4400 550.3000 1938.0400 550.7800 ;
        RECT 1936.4400 555.7400 1938.0400 556.2200 ;
        RECT 1936.4400 561.1800 1938.0400 561.6600 ;
        RECT 1920.9000 550.3000 1922.5000 550.7800 ;
        RECT 1920.9000 555.7400 1922.5000 556.2200 ;
        RECT 1920.9000 561.1800 1922.5000 561.6600 ;
        RECT 1936.4400 539.4200 1938.0400 539.9000 ;
        RECT 1936.4400 544.8600 1938.0400 545.3400 ;
        RECT 1920.9000 539.4200 1922.5000 539.9000 ;
        RECT 1920.9000 544.8600 1922.5000 545.3400 ;
        RECT 1936.4400 523.1000 1938.0400 523.5800 ;
        RECT 1936.4400 528.5400 1938.0400 529.0200 ;
        RECT 1936.4400 533.9800 1938.0400 534.4600 ;
        RECT 1920.9000 523.1000 1922.5000 523.5800 ;
        RECT 1920.9000 528.5400 1922.5000 529.0200 ;
        RECT 1920.9000 533.9800 1922.5000 534.4600 ;
        RECT 1875.9000 566.6200 1877.5000 567.1000 ;
        RECT 1875.9000 572.0600 1877.5000 572.5400 ;
        RECT 1875.9000 550.3000 1877.5000 550.7800 ;
        RECT 1875.9000 555.7400 1877.5000 556.2200 ;
        RECT 1875.9000 561.1800 1877.5000 561.6600 ;
        RECT 1875.9000 539.4200 1877.5000 539.9000 ;
        RECT 1875.9000 544.8600 1877.5000 545.3400 ;
        RECT 1875.9000 523.1000 1877.5000 523.5800 ;
        RECT 1875.9000 528.5400 1877.5000 529.0200 ;
        RECT 1875.9000 533.9800 1877.5000 534.4600 ;
        RECT 1875.9000 577.5000 1877.5000 577.9800 ;
        RECT 1920.9000 577.5000 1922.5000 577.9800 ;
        RECT 1936.4400 577.5000 1938.0400 577.9800 ;
        RECT 1830.9000 610.1400 1832.5000 610.6200 ;
        RECT 1830.9000 615.5800 1832.5000 616.0600 ;
        RECT 1830.9000 621.0200 1832.5000 621.5000 ;
        RECT 1785.9000 610.1400 1787.5000 610.6200 ;
        RECT 1785.9000 615.5800 1787.5000 616.0600 ;
        RECT 1785.9000 621.0200 1787.5000 621.5000 ;
        RECT 1830.9000 593.8200 1832.5000 594.3000 ;
        RECT 1830.9000 599.2600 1832.5000 599.7400 ;
        RECT 1830.9000 582.9400 1832.5000 583.4200 ;
        RECT 1830.9000 588.3800 1832.5000 588.8600 ;
        RECT 1785.9000 593.8200 1787.5000 594.3000 ;
        RECT 1785.9000 599.2600 1787.5000 599.7400 ;
        RECT 1785.9000 582.9400 1787.5000 583.4200 ;
        RECT 1785.9000 588.3800 1787.5000 588.8600 ;
        RECT 1785.9000 604.7000 1787.5000 605.1800 ;
        RECT 1830.9000 604.7000 1832.5000 605.1800 ;
        RECT 1733.7400 621.0200 1735.3400 621.5000 ;
        RECT 1740.9000 621.0200 1742.5000 621.5000 ;
        RECT 1740.9000 610.1400 1742.5000 610.6200 ;
        RECT 1740.9000 615.5800 1742.5000 616.0600 ;
        RECT 1733.7400 610.1400 1735.3400 610.6200 ;
        RECT 1733.7400 615.5800 1735.3400 616.0600 ;
        RECT 1740.9000 593.8200 1742.5000 594.3000 ;
        RECT 1740.9000 599.2600 1742.5000 599.7400 ;
        RECT 1733.7400 593.8200 1735.3400 594.3000 ;
        RECT 1733.7400 599.2600 1735.3400 599.7400 ;
        RECT 1740.9000 582.9400 1742.5000 583.4200 ;
        RECT 1740.9000 588.3800 1742.5000 588.8600 ;
        RECT 1733.7400 582.9400 1735.3400 583.4200 ;
        RECT 1733.7400 588.3800 1735.3400 588.8600 ;
        RECT 1733.7400 604.7000 1735.3400 605.1800 ;
        RECT 1740.9000 604.7000 1742.5000 605.1800 ;
        RECT 1830.9000 566.6200 1832.5000 567.1000 ;
        RECT 1830.9000 572.0600 1832.5000 572.5400 ;
        RECT 1830.9000 550.3000 1832.5000 550.7800 ;
        RECT 1830.9000 555.7400 1832.5000 556.2200 ;
        RECT 1830.9000 561.1800 1832.5000 561.6600 ;
        RECT 1785.9000 566.6200 1787.5000 567.1000 ;
        RECT 1785.9000 572.0600 1787.5000 572.5400 ;
        RECT 1785.9000 550.3000 1787.5000 550.7800 ;
        RECT 1785.9000 555.7400 1787.5000 556.2200 ;
        RECT 1785.9000 561.1800 1787.5000 561.6600 ;
        RECT 1830.9000 539.4200 1832.5000 539.9000 ;
        RECT 1830.9000 544.8600 1832.5000 545.3400 ;
        RECT 1830.9000 523.1000 1832.5000 523.5800 ;
        RECT 1830.9000 528.5400 1832.5000 529.0200 ;
        RECT 1830.9000 533.9800 1832.5000 534.4600 ;
        RECT 1785.9000 539.4200 1787.5000 539.9000 ;
        RECT 1785.9000 544.8600 1787.5000 545.3400 ;
        RECT 1785.9000 523.1000 1787.5000 523.5800 ;
        RECT 1785.9000 528.5400 1787.5000 529.0200 ;
        RECT 1785.9000 533.9800 1787.5000 534.4600 ;
        RECT 1740.9000 566.6200 1742.5000 567.1000 ;
        RECT 1740.9000 572.0600 1742.5000 572.5400 ;
        RECT 1733.7400 566.6200 1735.3400 567.1000 ;
        RECT 1733.7400 572.0600 1735.3400 572.5400 ;
        RECT 1740.9000 550.3000 1742.5000 550.7800 ;
        RECT 1740.9000 555.7400 1742.5000 556.2200 ;
        RECT 1740.9000 561.1800 1742.5000 561.6600 ;
        RECT 1733.7400 550.3000 1735.3400 550.7800 ;
        RECT 1733.7400 555.7400 1735.3400 556.2200 ;
        RECT 1733.7400 561.1800 1735.3400 561.6600 ;
        RECT 1740.9000 539.4200 1742.5000 539.9000 ;
        RECT 1740.9000 544.8600 1742.5000 545.3400 ;
        RECT 1733.7400 539.4200 1735.3400 539.9000 ;
        RECT 1733.7400 544.8600 1735.3400 545.3400 ;
        RECT 1740.9000 523.1000 1742.5000 523.5800 ;
        RECT 1740.9000 528.5400 1742.5000 529.0200 ;
        RECT 1740.9000 533.9800 1742.5000 534.4600 ;
        RECT 1733.7400 523.1000 1735.3400 523.5800 ;
        RECT 1733.7400 528.5400 1735.3400 529.0200 ;
        RECT 1733.7400 533.9800 1735.3400 534.4600 ;
        RECT 1733.7400 577.5000 1735.3400 577.9800 ;
        RECT 1740.9000 577.5000 1742.5000 577.9800 ;
        RECT 1785.9000 577.5000 1787.5000 577.9800 ;
        RECT 1830.9000 577.5000 1832.5000 577.9800 ;
        RECT 1936.4400 512.2200 1938.0400 512.7000 ;
        RECT 1936.4400 517.6600 1938.0400 518.1400 ;
        RECT 1920.9000 512.2200 1922.5000 512.7000 ;
        RECT 1920.9000 517.6600 1922.5000 518.1400 ;
        RECT 1936.4400 495.9000 1938.0400 496.3800 ;
        RECT 1936.4400 501.3400 1938.0400 501.8200 ;
        RECT 1936.4400 506.7800 1938.0400 507.2600 ;
        RECT 1920.9000 495.9000 1922.5000 496.3800 ;
        RECT 1920.9000 501.3400 1922.5000 501.8200 ;
        RECT 1920.9000 506.7800 1922.5000 507.2600 ;
        RECT 1936.4400 485.0200 1938.0400 485.5000 ;
        RECT 1936.4400 490.4600 1938.0400 490.9400 ;
        RECT 1920.9000 485.0200 1922.5000 485.5000 ;
        RECT 1920.9000 490.4600 1922.5000 490.9400 ;
        RECT 1936.4400 468.7000 1938.0400 469.1800 ;
        RECT 1936.4400 474.1400 1938.0400 474.6200 ;
        RECT 1936.4400 479.5800 1938.0400 480.0600 ;
        RECT 1920.9000 468.7000 1922.5000 469.1800 ;
        RECT 1920.9000 474.1400 1922.5000 474.6200 ;
        RECT 1920.9000 479.5800 1922.5000 480.0600 ;
        RECT 1875.9000 512.2200 1877.5000 512.7000 ;
        RECT 1875.9000 517.6600 1877.5000 518.1400 ;
        RECT 1875.9000 495.9000 1877.5000 496.3800 ;
        RECT 1875.9000 501.3400 1877.5000 501.8200 ;
        RECT 1875.9000 506.7800 1877.5000 507.2600 ;
        RECT 1875.9000 485.0200 1877.5000 485.5000 ;
        RECT 1875.9000 490.4600 1877.5000 490.9400 ;
        RECT 1875.9000 468.7000 1877.5000 469.1800 ;
        RECT 1875.9000 474.1400 1877.5000 474.6200 ;
        RECT 1875.9000 479.5800 1877.5000 480.0600 ;
        RECT 1936.4400 457.8200 1938.0400 458.3000 ;
        RECT 1936.4400 463.2600 1938.0400 463.7400 ;
        RECT 1920.9000 457.8200 1922.5000 458.3000 ;
        RECT 1920.9000 463.2600 1922.5000 463.7400 ;
        RECT 1936.4400 441.5000 1938.0400 441.9800 ;
        RECT 1936.4400 446.9400 1938.0400 447.4200 ;
        RECT 1936.4400 452.3800 1938.0400 452.8600 ;
        RECT 1920.9000 441.5000 1922.5000 441.9800 ;
        RECT 1920.9000 446.9400 1922.5000 447.4200 ;
        RECT 1920.9000 452.3800 1922.5000 452.8600 ;
        RECT 1936.4400 430.6200 1938.0400 431.1000 ;
        RECT 1936.4400 436.0600 1938.0400 436.5400 ;
        RECT 1920.9000 430.6200 1922.5000 431.1000 ;
        RECT 1920.9000 436.0600 1922.5000 436.5400 ;
        RECT 1920.9000 425.1800 1922.5000 425.6600 ;
        RECT 1936.4400 425.1800 1938.0400 425.6600 ;
        RECT 1875.9000 457.8200 1877.5000 458.3000 ;
        RECT 1875.9000 463.2600 1877.5000 463.7400 ;
        RECT 1875.9000 441.5000 1877.5000 441.9800 ;
        RECT 1875.9000 446.9400 1877.5000 447.4200 ;
        RECT 1875.9000 452.3800 1877.5000 452.8600 ;
        RECT 1875.9000 430.6200 1877.5000 431.1000 ;
        RECT 1875.9000 436.0600 1877.5000 436.5400 ;
        RECT 1875.9000 425.1800 1877.5000 425.6600 ;
        RECT 1830.9000 512.2200 1832.5000 512.7000 ;
        RECT 1830.9000 517.6600 1832.5000 518.1400 ;
        RECT 1830.9000 495.9000 1832.5000 496.3800 ;
        RECT 1830.9000 501.3400 1832.5000 501.8200 ;
        RECT 1830.9000 506.7800 1832.5000 507.2600 ;
        RECT 1785.9000 512.2200 1787.5000 512.7000 ;
        RECT 1785.9000 517.6600 1787.5000 518.1400 ;
        RECT 1785.9000 495.9000 1787.5000 496.3800 ;
        RECT 1785.9000 501.3400 1787.5000 501.8200 ;
        RECT 1785.9000 506.7800 1787.5000 507.2600 ;
        RECT 1830.9000 485.0200 1832.5000 485.5000 ;
        RECT 1830.9000 490.4600 1832.5000 490.9400 ;
        RECT 1830.9000 468.7000 1832.5000 469.1800 ;
        RECT 1830.9000 474.1400 1832.5000 474.6200 ;
        RECT 1830.9000 479.5800 1832.5000 480.0600 ;
        RECT 1785.9000 485.0200 1787.5000 485.5000 ;
        RECT 1785.9000 490.4600 1787.5000 490.9400 ;
        RECT 1785.9000 468.7000 1787.5000 469.1800 ;
        RECT 1785.9000 474.1400 1787.5000 474.6200 ;
        RECT 1785.9000 479.5800 1787.5000 480.0600 ;
        RECT 1740.9000 512.2200 1742.5000 512.7000 ;
        RECT 1740.9000 517.6600 1742.5000 518.1400 ;
        RECT 1733.7400 512.2200 1735.3400 512.7000 ;
        RECT 1733.7400 517.6600 1735.3400 518.1400 ;
        RECT 1740.9000 495.9000 1742.5000 496.3800 ;
        RECT 1740.9000 501.3400 1742.5000 501.8200 ;
        RECT 1740.9000 506.7800 1742.5000 507.2600 ;
        RECT 1733.7400 495.9000 1735.3400 496.3800 ;
        RECT 1733.7400 501.3400 1735.3400 501.8200 ;
        RECT 1733.7400 506.7800 1735.3400 507.2600 ;
        RECT 1740.9000 485.0200 1742.5000 485.5000 ;
        RECT 1740.9000 490.4600 1742.5000 490.9400 ;
        RECT 1733.7400 485.0200 1735.3400 485.5000 ;
        RECT 1733.7400 490.4600 1735.3400 490.9400 ;
        RECT 1740.9000 468.7000 1742.5000 469.1800 ;
        RECT 1740.9000 474.1400 1742.5000 474.6200 ;
        RECT 1740.9000 479.5800 1742.5000 480.0600 ;
        RECT 1733.7400 468.7000 1735.3400 469.1800 ;
        RECT 1733.7400 474.1400 1735.3400 474.6200 ;
        RECT 1733.7400 479.5800 1735.3400 480.0600 ;
        RECT 1830.9000 457.8200 1832.5000 458.3000 ;
        RECT 1830.9000 463.2600 1832.5000 463.7400 ;
        RECT 1830.9000 441.5000 1832.5000 441.9800 ;
        RECT 1830.9000 446.9400 1832.5000 447.4200 ;
        RECT 1830.9000 452.3800 1832.5000 452.8600 ;
        RECT 1785.9000 457.8200 1787.5000 458.3000 ;
        RECT 1785.9000 463.2600 1787.5000 463.7400 ;
        RECT 1785.9000 441.5000 1787.5000 441.9800 ;
        RECT 1785.9000 446.9400 1787.5000 447.4200 ;
        RECT 1785.9000 452.3800 1787.5000 452.8600 ;
        RECT 1830.9000 436.0600 1832.5000 436.5400 ;
        RECT 1830.9000 430.6200 1832.5000 431.1000 ;
        RECT 1830.9000 425.1800 1832.5000 425.6600 ;
        RECT 1785.9000 436.0600 1787.5000 436.5400 ;
        RECT 1785.9000 430.6200 1787.5000 431.1000 ;
        RECT 1785.9000 425.1800 1787.5000 425.6600 ;
        RECT 1740.9000 457.8200 1742.5000 458.3000 ;
        RECT 1740.9000 463.2600 1742.5000 463.7400 ;
        RECT 1733.7400 457.8200 1735.3400 458.3000 ;
        RECT 1733.7400 463.2600 1735.3400 463.7400 ;
        RECT 1740.9000 441.5000 1742.5000 441.9800 ;
        RECT 1740.9000 446.9400 1742.5000 447.4200 ;
        RECT 1740.9000 452.3800 1742.5000 452.8600 ;
        RECT 1733.7400 441.5000 1735.3400 441.9800 ;
        RECT 1733.7400 446.9400 1735.3400 447.4200 ;
        RECT 1733.7400 452.3800 1735.3400 452.8600 ;
        RECT 1740.9000 430.6200 1742.5000 431.1000 ;
        RECT 1740.9000 436.0600 1742.5000 436.5400 ;
        RECT 1733.7400 430.6200 1735.3400 431.1000 ;
        RECT 1733.7400 436.0600 1735.3400 436.5400 ;
        RECT 1733.7400 425.1800 1735.3400 425.6600 ;
        RECT 1740.9000 425.1800 1742.5000 425.6600 ;
        RECT 1730.7800 627.3700 1941.0000 628.9700 ;
        RECT 1730.7800 415.6700 1941.0000 417.2700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 412.8400 1735.3400 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.7400 630.8800 1735.3400 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 412.8400 1938.0400 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1936.4400 630.8800 1938.0400 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 415.6700 1732.3800 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 415.6700 1941.0000 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 627.3700 1732.3800 628.9700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 627.3700 1941.0000 628.9700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1954.0600 2479.6000 1955.6600 2509.8600 ;
        RECT 2156.5600 2479.6000 2158.1600 2509.8600 ;
      LAYER met3 ;
        RECT 2156.5600 2500.1000 2158.1600 2500.5800 ;
        RECT 1954.0600 2500.1000 1955.6600 2500.5800 ;
        RECT 2156.5600 2489.2200 2158.1600 2489.7000 ;
        RECT 1954.0600 2489.2200 1955.6600 2489.7000 ;
        RECT 2156.5600 2494.6600 2158.1600 2495.1400 ;
        RECT 1954.0600 2494.6600 1955.6600 2495.1400 ;
        RECT 1951.0000 2505.5000 2161.2200 2507.1000 ;
        RECT 1951.0000 2481.1700 2161.2200 2482.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.0600 2479.6000 1955.6600 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.0600 2508.2600 1955.6600 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.5600 2479.6000 2158.1600 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.5600 2508.2600 2158.1600 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2481.1700 1952.6000 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2481.1700 2161.2200 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2505.5000 1952.6000 2507.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2505.5000 2161.2200 2507.1000 ;
    END
# end of P/G pin shape extracted from block 'N_term_DSP'


# P/G pin shape extracted from block 'S_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1954.0600 142.9400 1955.6600 173.2000 ;
        RECT 2156.5600 142.9400 2158.1600 173.2000 ;
      LAYER met3 ;
        RECT 2156.5600 163.4400 2158.1600 163.9200 ;
        RECT 1954.0600 163.4400 1955.6600 163.9200 ;
        RECT 2156.5600 152.5600 2158.1600 153.0400 ;
        RECT 1954.0600 152.5600 1955.6600 153.0400 ;
        RECT 2156.5600 158.0000 2158.1600 158.4800 ;
        RECT 1954.0600 158.0000 1955.6600 158.4800 ;
        RECT 1951.0000 168.8400 2161.2200 170.4400 ;
        RECT 1951.0000 144.5100 2161.2200 146.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.0600 142.9400 1955.6600 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1954.0600 171.6000 1955.6600 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.5600 142.9400 2158.1600 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.5600 171.6000 2158.1600 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 144.5100 1952.6000 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 144.5100 2161.2200 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 168.8400 1952.6000 170.4400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 168.8400 2161.2200 170.4400 ;
    END
# end of P/G pin shape extracted from block 'S_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1953.9600 2020.3200 1955.5600 2470.1400 ;
        RECT 2156.6600 2020.3200 2158.2600 2470.1400 ;
        RECT 1961.1200 2023.1500 1962.7200 2467.1400 ;
        RECT 2006.1200 2023.1500 2007.7200 2467.1400 ;
        RECT 2051.1200 2023.1500 2052.7200 2467.1400 ;
        RECT 2096.1200 2023.1500 2097.7200 2467.1400 ;
        RECT 2141.1200 2023.1500 2142.7200 2467.1400 ;
      LAYER met3 ;
        RECT 2156.6600 2456.9800 2158.2600 2457.4600 ;
        RECT 2156.6600 2451.5400 2158.2600 2452.0200 ;
        RECT 2156.6600 2446.1000 2158.2600 2446.5800 ;
        RECT 2156.6600 2440.6600 2158.2600 2441.1400 ;
        RECT 2156.6600 2435.2200 2158.2600 2435.7000 ;
        RECT 2156.6600 2429.7800 2158.2600 2430.2600 ;
        RECT 2156.6600 2424.3400 2158.2600 2424.8200 ;
        RECT 2156.6600 2418.9000 2158.2600 2419.3800 ;
        RECT 2156.6600 2408.0200 2158.2600 2408.5000 ;
        RECT 2156.6600 2402.5800 2158.2600 2403.0600 ;
        RECT 2156.6600 2397.1400 2158.2600 2397.6200 ;
        RECT 2156.6600 2391.7000 2158.2600 2392.1800 ;
        RECT 2156.6600 2386.2600 2158.2600 2386.7400 ;
        RECT 2156.6600 2380.8200 2158.2600 2381.3000 ;
        RECT 2156.6600 2375.3800 2158.2600 2375.8600 ;
        RECT 2156.6600 2369.9400 2158.2600 2370.4200 ;
        RECT 2156.6600 2364.5000 2158.2600 2364.9800 ;
        RECT 2156.6600 2359.0600 2158.2600 2359.5400 ;
        RECT 2156.6600 2413.4600 2158.2600 2413.9400 ;
        RECT 2156.6600 2353.6200 2158.2600 2354.1000 ;
        RECT 2156.6600 2348.1800 2158.2600 2348.6600 ;
        RECT 2156.6600 2342.7400 2158.2600 2343.2200 ;
        RECT 2156.6600 2337.3000 2158.2600 2337.7800 ;
        RECT 2156.6600 2331.8600 2158.2600 2332.3400 ;
        RECT 2156.6600 2326.4200 2158.2600 2326.9000 ;
        RECT 2156.6600 2320.9800 2158.2600 2321.4600 ;
        RECT 2156.6600 2315.5400 2158.2600 2316.0200 ;
        RECT 2156.6600 2310.1000 2158.2600 2310.5800 ;
        RECT 2156.6600 2304.6600 2158.2600 2305.1400 ;
        RECT 2156.6600 2299.2200 2158.2600 2299.7000 ;
        RECT 2156.6600 2293.7800 2158.2600 2294.2600 ;
        RECT 2156.6600 2288.3400 2158.2600 2288.8200 ;
        RECT 2156.6600 2282.9000 2158.2600 2283.3800 ;
        RECT 2156.6600 2277.4600 2158.2600 2277.9400 ;
        RECT 2156.6600 2272.0200 2158.2600 2272.5000 ;
        RECT 2156.6600 2266.5800 2158.2600 2267.0600 ;
        RECT 2156.6600 2261.1400 2158.2600 2261.6200 ;
        RECT 2156.6600 2255.7000 2158.2600 2256.1800 ;
        RECT 2156.6600 2250.2600 2158.2600 2250.7400 ;
        RECT 1953.9600 2456.9800 1955.5600 2457.4600 ;
        RECT 1953.9600 2451.5400 1955.5600 2452.0200 ;
        RECT 1953.9600 2446.1000 1955.5600 2446.5800 ;
        RECT 1953.9600 2440.6600 1955.5600 2441.1400 ;
        RECT 1953.9600 2435.2200 1955.5600 2435.7000 ;
        RECT 1953.9600 2429.7800 1955.5600 2430.2600 ;
        RECT 1953.9600 2424.3400 1955.5600 2424.8200 ;
        RECT 1953.9600 2418.9000 1955.5600 2419.3800 ;
        RECT 1953.9600 2408.0200 1955.5600 2408.5000 ;
        RECT 1953.9600 2402.5800 1955.5600 2403.0600 ;
        RECT 1953.9600 2397.1400 1955.5600 2397.6200 ;
        RECT 1953.9600 2391.7000 1955.5600 2392.1800 ;
        RECT 1953.9600 2386.2600 1955.5600 2386.7400 ;
        RECT 1953.9600 2380.8200 1955.5600 2381.3000 ;
        RECT 1953.9600 2375.3800 1955.5600 2375.8600 ;
        RECT 1953.9600 2369.9400 1955.5600 2370.4200 ;
        RECT 1953.9600 2364.5000 1955.5600 2364.9800 ;
        RECT 1953.9600 2359.0600 1955.5600 2359.5400 ;
        RECT 1953.9600 2413.4600 1955.5600 2413.9400 ;
        RECT 1953.9600 2353.6200 1955.5600 2354.1000 ;
        RECT 1953.9600 2348.1800 1955.5600 2348.6600 ;
        RECT 1953.9600 2342.7400 1955.5600 2343.2200 ;
        RECT 1953.9600 2337.3000 1955.5600 2337.7800 ;
        RECT 1953.9600 2331.8600 1955.5600 2332.3400 ;
        RECT 1953.9600 2326.4200 1955.5600 2326.9000 ;
        RECT 1953.9600 2320.9800 1955.5600 2321.4600 ;
        RECT 1953.9600 2315.5400 1955.5600 2316.0200 ;
        RECT 1953.9600 2310.1000 1955.5600 2310.5800 ;
        RECT 1953.9600 2304.6600 1955.5600 2305.1400 ;
        RECT 1953.9600 2299.2200 1955.5600 2299.7000 ;
        RECT 1953.9600 2293.7800 1955.5600 2294.2600 ;
        RECT 1953.9600 2288.3400 1955.5600 2288.8200 ;
        RECT 1953.9600 2282.9000 1955.5600 2283.3800 ;
        RECT 1953.9600 2277.4600 1955.5600 2277.9400 ;
        RECT 1953.9600 2272.0200 1955.5600 2272.5000 ;
        RECT 1953.9600 2266.5800 1955.5600 2267.0600 ;
        RECT 1953.9600 2261.1400 1955.5600 2261.6200 ;
        RECT 1953.9600 2255.7000 1955.5600 2256.1800 ;
        RECT 1953.9600 2250.2600 1955.5600 2250.7400 ;
        RECT 2156.6600 2239.3800 2158.2600 2239.8600 ;
        RECT 2156.6600 2233.9400 2158.2600 2234.4200 ;
        RECT 2156.6600 2228.5000 2158.2600 2228.9800 ;
        RECT 2156.6600 2223.0600 2158.2600 2223.5400 ;
        RECT 2156.6600 2217.6200 2158.2600 2218.1000 ;
        RECT 2156.6600 2212.1800 2158.2600 2212.6600 ;
        RECT 2156.6600 2206.7400 2158.2600 2207.2200 ;
        RECT 2156.6600 2201.3000 2158.2600 2201.7800 ;
        RECT 2156.6600 2195.8600 2158.2600 2196.3400 ;
        RECT 2156.6600 2190.4200 2158.2600 2190.9000 ;
        RECT 2156.6600 2184.9800 2158.2600 2185.4600 ;
        RECT 2156.6600 2179.5400 2158.2600 2180.0200 ;
        RECT 2156.6600 2174.1000 2158.2600 2174.5800 ;
        RECT 2156.6600 2168.6600 2158.2600 2169.1400 ;
        RECT 2156.6600 2163.2200 2158.2600 2163.7000 ;
        RECT 2156.6600 2157.7800 2158.2600 2158.2600 ;
        RECT 2156.6600 2152.3400 2158.2600 2152.8200 ;
        RECT 2156.6600 2146.9000 2158.2600 2147.3800 ;
        RECT 2156.6600 2141.4600 2158.2600 2141.9400 ;
        RECT 2156.6600 2136.0200 2158.2600 2136.5000 ;
        RECT 2156.6600 2130.5800 2158.2600 2131.0600 ;
        RECT 2156.6600 2125.1400 2158.2600 2125.6200 ;
        RECT 2156.6600 2119.7000 2158.2600 2120.1800 ;
        RECT 2156.6600 2114.2600 2158.2600 2114.7400 ;
        RECT 2156.6600 2108.8200 2158.2600 2109.3000 ;
        RECT 2156.6600 2103.3800 2158.2600 2103.8600 ;
        RECT 2156.6600 2097.9400 2158.2600 2098.4200 ;
        RECT 2156.6600 2092.5000 2158.2600 2092.9800 ;
        RECT 2156.6600 2087.0600 2158.2600 2087.5400 ;
        RECT 2156.6600 2081.6200 2158.2600 2082.1000 ;
        RECT 2156.6600 2070.7400 2158.2600 2071.2200 ;
        RECT 2156.6600 2065.3000 2158.2600 2065.7800 ;
        RECT 2156.6600 2059.8600 2158.2600 2060.3400 ;
        RECT 2156.6600 2054.4200 2158.2600 2054.9000 ;
        RECT 2156.6600 2048.9800 2158.2600 2049.4600 ;
        RECT 2156.6600 2043.5400 2158.2600 2044.0200 ;
        RECT 2156.6600 2038.1000 2158.2600 2038.5800 ;
        RECT 2156.6600 2032.6600 2158.2600 2033.1400 ;
        RECT 2156.6600 2076.1800 2158.2600 2076.6600 ;
        RECT 1953.9600 2239.3800 1955.5600 2239.8600 ;
        RECT 1953.9600 2233.9400 1955.5600 2234.4200 ;
        RECT 1953.9600 2228.5000 1955.5600 2228.9800 ;
        RECT 1953.9600 2223.0600 1955.5600 2223.5400 ;
        RECT 1953.9600 2217.6200 1955.5600 2218.1000 ;
        RECT 1953.9600 2212.1800 1955.5600 2212.6600 ;
        RECT 1953.9600 2206.7400 1955.5600 2207.2200 ;
        RECT 1953.9600 2201.3000 1955.5600 2201.7800 ;
        RECT 1953.9600 2195.8600 1955.5600 2196.3400 ;
        RECT 1953.9600 2190.4200 1955.5600 2190.9000 ;
        RECT 1953.9600 2184.9800 1955.5600 2185.4600 ;
        RECT 1953.9600 2179.5400 1955.5600 2180.0200 ;
        RECT 1953.9600 2174.1000 1955.5600 2174.5800 ;
        RECT 1953.9600 2168.6600 1955.5600 2169.1400 ;
        RECT 1953.9600 2163.2200 1955.5600 2163.7000 ;
        RECT 1953.9600 2157.7800 1955.5600 2158.2600 ;
        RECT 1953.9600 2152.3400 1955.5600 2152.8200 ;
        RECT 1953.9600 2146.9000 1955.5600 2147.3800 ;
        RECT 1953.9600 2141.4600 1955.5600 2141.9400 ;
        RECT 1953.9600 2136.0200 1955.5600 2136.5000 ;
        RECT 1953.9600 2130.5800 1955.5600 2131.0600 ;
        RECT 1953.9600 2125.1400 1955.5600 2125.6200 ;
        RECT 1953.9600 2119.7000 1955.5600 2120.1800 ;
        RECT 1953.9600 2114.2600 1955.5600 2114.7400 ;
        RECT 1953.9600 2108.8200 1955.5600 2109.3000 ;
        RECT 1953.9600 2103.3800 1955.5600 2103.8600 ;
        RECT 1953.9600 2097.9400 1955.5600 2098.4200 ;
        RECT 1953.9600 2092.5000 1955.5600 2092.9800 ;
        RECT 1953.9600 2087.0600 1955.5600 2087.5400 ;
        RECT 1953.9600 2081.6200 1955.5600 2082.1000 ;
        RECT 1953.9600 2070.7400 1955.5600 2071.2200 ;
        RECT 1953.9600 2065.3000 1955.5600 2065.7800 ;
        RECT 1953.9600 2059.8600 1955.5600 2060.3400 ;
        RECT 1953.9600 2054.4200 1955.5600 2054.9000 ;
        RECT 1953.9600 2048.9800 1955.5600 2049.4600 ;
        RECT 1953.9600 2043.5400 1955.5600 2044.0200 ;
        RECT 1953.9600 2038.1000 1955.5600 2038.5800 ;
        RECT 1953.9600 2032.6600 1955.5600 2033.1400 ;
        RECT 1953.9600 2076.1800 1955.5600 2076.6600 ;
        RECT 2156.6600 2244.8200 2158.2600 2245.3000 ;
        RECT 1953.9600 2244.8200 1955.5600 2245.3000 ;
        RECT 1951.0000 2465.5400 2161.2200 2467.1400 ;
        RECT 1951.0000 2023.1500 2161.2200 2024.7500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 2020.3200 1955.5600 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 2468.5400 1955.5600 2470.1400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 2020.3200 2158.2600 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 2468.5400 2158.2600 2470.1400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2023.1500 1952.6000 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2023.1500 2161.2200 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2465.5400 1952.6000 2467.1400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2465.5400 2161.2200 2467.1400 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1953.9600 1561.0400 1955.5600 2010.8600 ;
        RECT 2156.6600 1561.0400 2158.2600 2010.8600 ;
        RECT 1961.1200 1563.8700 1962.7200 2007.8600 ;
        RECT 2006.1200 1563.8700 2007.7200 2007.8600 ;
        RECT 2051.1200 1563.8700 2052.7200 2007.8600 ;
        RECT 2096.1200 1563.8700 2097.7200 2007.8600 ;
        RECT 2141.1200 1563.8700 2142.7200 2007.8600 ;
      LAYER met3 ;
        RECT 2156.6600 1997.7000 2158.2600 1998.1800 ;
        RECT 2156.6600 1992.2600 2158.2600 1992.7400 ;
        RECT 2156.6600 1986.8200 2158.2600 1987.3000 ;
        RECT 2156.6600 1981.3800 2158.2600 1981.8600 ;
        RECT 2156.6600 1975.9400 2158.2600 1976.4200 ;
        RECT 2156.6600 1970.5000 2158.2600 1970.9800 ;
        RECT 2156.6600 1965.0600 2158.2600 1965.5400 ;
        RECT 2156.6600 1959.6200 2158.2600 1960.1000 ;
        RECT 2156.6600 1948.7400 2158.2600 1949.2200 ;
        RECT 2156.6600 1943.3000 2158.2600 1943.7800 ;
        RECT 2156.6600 1937.8600 2158.2600 1938.3400 ;
        RECT 2156.6600 1932.4200 2158.2600 1932.9000 ;
        RECT 2156.6600 1926.9800 2158.2600 1927.4600 ;
        RECT 2156.6600 1921.5400 2158.2600 1922.0200 ;
        RECT 2156.6600 1916.1000 2158.2600 1916.5800 ;
        RECT 2156.6600 1910.6600 2158.2600 1911.1400 ;
        RECT 2156.6600 1905.2200 2158.2600 1905.7000 ;
        RECT 2156.6600 1899.7800 2158.2600 1900.2600 ;
        RECT 2156.6600 1954.1800 2158.2600 1954.6600 ;
        RECT 2156.6600 1894.3400 2158.2600 1894.8200 ;
        RECT 2156.6600 1888.9000 2158.2600 1889.3800 ;
        RECT 2156.6600 1883.4600 2158.2600 1883.9400 ;
        RECT 2156.6600 1878.0200 2158.2600 1878.5000 ;
        RECT 2156.6600 1872.5800 2158.2600 1873.0600 ;
        RECT 2156.6600 1867.1400 2158.2600 1867.6200 ;
        RECT 2156.6600 1861.7000 2158.2600 1862.1800 ;
        RECT 2156.6600 1856.2600 2158.2600 1856.7400 ;
        RECT 2156.6600 1850.8200 2158.2600 1851.3000 ;
        RECT 2156.6600 1845.3800 2158.2600 1845.8600 ;
        RECT 2156.6600 1839.9400 2158.2600 1840.4200 ;
        RECT 2156.6600 1834.5000 2158.2600 1834.9800 ;
        RECT 2156.6600 1829.0600 2158.2600 1829.5400 ;
        RECT 2156.6600 1823.6200 2158.2600 1824.1000 ;
        RECT 2156.6600 1818.1800 2158.2600 1818.6600 ;
        RECT 2156.6600 1812.7400 2158.2600 1813.2200 ;
        RECT 2156.6600 1807.3000 2158.2600 1807.7800 ;
        RECT 2156.6600 1801.8600 2158.2600 1802.3400 ;
        RECT 2156.6600 1796.4200 2158.2600 1796.9000 ;
        RECT 2156.6600 1790.9800 2158.2600 1791.4600 ;
        RECT 1953.9600 1997.7000 1955.5600 1998.1800 ;
        RECT 1953.9600 1992.2600 1955.5600 1992.7400 ;
        RECT 1953.9600 1986.8200 1955.5600 1987.3000 ;
        RECT 1953.9600 1981.3800 1955.5600 1981.8600 ;
        RECT 1953.9600 1975.9400 1955.5600 1976.4200 ;
        RECT 1953.9600 1970.5000 1955.5600 1970.9800 ;
        RECT 1953.9600 1965.0600 1955.5600 1965.5400 ;
        RECT 1953.9600 1959.6200 1955.5600 1960.1000 ;
        RECT 1953.9600 1948.7400 1955.5600 1949.2200 ;
        RECT 1953.9600 1943.3000 1955.5600 1943.7800 ;
        RECT 1953.9600 1937.8600 1955.5600 1938.3400 ;
        RECT 1953.9600 1932.4200 1955.5600 1932.9000 ;
        RECT 1953.9600 1926.9800 1955.5600 1927.4600 ;
        RECT 1953.9600 1921.5400 1955.5600 1922.0200 ;
        RECT 1953.9600 1916.1000 1955.5600 1916.5800 ;
        RECT 1953.9600 1910.6600 1955.5600 1911.1400 ;
        RECT 1953.9600 1905.2200 1955.5600 1905.7000 ;
        RECT 1953.9600 1899.7800 1955.5600 1900.2600 ;
        RECT 1953.9600 1954.1800 1955.5600 1954.6600 ;
        RECT 1953.9600 1894.3400 1955.5600 1894.8200 ;
        RECT 1953.9600 1888.9000 1955.5600 1889.3800 ;
        RECT 1953.9600 1883.4600 1955.5600 1883.9400 ;
        RECT 1953.9600 1878.0200 1955.5600 1878.5000 ;
        RECT 1953.9600 1872.5800 1955.5600 1873.0600 ;
        RECT 1953.9600 1867.1400 1955.5600 1867.6200 ;
        RECT 1953.9600 1861.7000 1955.5600 1862.1800 ;
        RECT 1953.9600 1856.2600 1955.5600 1856.7400 ;
        RECT 1953.9600 1850.8200 1955.5600 1851.3000 ;
        RECT 1953.9600 1845.3800 1955.5600 1845.8600 ;
        RECT 1953.9600 1839.9400 1955.5600 1840.4200 ;
        RECT 1953.9600 1834.5000 1955.5600 1834.9800 ;
        RECT 1953.9600 1829.0600 1955.5600 1829.5400 ;
        RECT 1953.9600 1823.6200 1955.5600 1824.1000 ;
        RECT 1953.9600 1818.1800 1955.5600 1818.6600 ;
        RECT 1953.9600 1812.7400 1955.5600 1813.2200 ;
        RECT 1953.9600 1807.3000 1955.5600 1807.7800 ;
        RECT 1953.9600 1801.8600 1955.5600 1802.3400 ;
        RECT 1953.9600 1796.4200 1955.5600 1796.9000 ;
        RECT 1953.9600 1790.9800 1955.5600 1791.4600 ;
        RECT 2156.6600 1780.1000 2158.2600 1780.5800 ;
        RECT 2156.6600 1774.6600 2158.2600 1775.1400 ;
        RECT 2156.6600 1769.2200 2158.2600 1769.7000 ;
        RECT 2156.6600 1763.7800 2158.2600 1764.2600 ;
        RECT 2156.6600 1758.3400 2158.2600 1758.8200 ;
        RECT 2156.6600 1752.9000 2158.2600 1753.3800 ;
        RECT 2156.6600 1747.4600 2158.2600 1747.9400 ;
        RECT 2156.6600 1742.0200 2158.2600 1742.5000 ;
        RECT 2156.6600 1736.5800 2158.2600 1737.0600 ;
        RECT 2156.6600 1731.1400 2158.2600 1731.6200 ;
        RECT 2156.6600 1725.7000 2158.2600 1726.1800 ;
        RECT 2156.6600 1720.2600 2158.2600 1720.7400 ;
        RECT 2156.6600 1714.8200 2158.2600 1715.3000 ;
        RECT 2156.6600 1709.3800 2158.2600 1709.8600 ;
        RECT 2156.6600 1703.9400 2158.2600 1704.4200 ;
        RECT 2156.6600 1698.5000 2158.2600 1698.9800 ;
        RECT 2156.6600 1693.0600 2158.2600 1693.5400 ;
        RECT 2156.6600 1687.6200 2158.2600 1688.1000 ;
        RECT 2156.6600 1682.1800 2158.2600 1682.6600 ;
        RECT 2156.6600 1676.7400 2158.2600 1677.2200 ;
        RECT 2156.6600 1671.3000 2158.2600 1671.7800 ;
        RECT 2156.6600 1665.8600 2158.2600 1666.3400 ;
        RECT 2156.6600 1660.4200 2158.2600 1660.9000 ;
        RECT 2156.6600 1654.9800 2158.2600 1655.4600 ;
        RECT 2156.6600 1649.5400 2158.2600 1650.0200 ;
        RECT 2156.6600 1644.1000 2158.2600 1644.5800 ;
        RECT 2156.6600 1638.6600 2158.2600 1639.1400 ;
        RECT 2156.6600 1633.2200 2158.2600 1633.7000 ;
        RECT 2156.6600 1627.7800 2158.2600 1628.2600 ;
        RECT 2156.6600 1622.3400 2158.2600 1622.8200 ;
        RECT 2156.6600 1611.4600 2158.2600 1611.9400 ;
        RECT 2156.6600 1606.0200 2158.2600 1606.5000 ;
        RECT 2156.6600 1600.5800 2158.2600 1601.0600 ;
        RECT 2156.6600 1595.1400 2158.2600 1595.6200 ;
        RECT 2156.6600 1589.7000 2158.2600 1590.1800 ;
        RECT 2156.6600 1584.2600 2158.2600 1584.7400 ;
        RECT 2156.6600 1578.8200 2158.2600 1579.3000 ;
        RECT 2156.6600 1573.3800 2158.2600 1573.8600 ;
        RECT 2156.6600 1616.9000 2158.2600 1617.3800 ;
        RECT 1953.9600 1780.1000 1955.5600 1780.5800 ;
        RECT 1953.9600 1774.6600 1955.5600 1775.1400 ;
        RECT 1953.9600 1769.2200 1955.5600 1769.7000 ;
        RECT 1953.9600 1763.7800 1955.5600 1764.2600 ;
        RECT 1953.9600 1758.3400 1955.5600 1758.8200 ;
        RECT 1953.9600 1752.9000 1955.5600 1753.3800 ;
        RECT 1953.9600 1747.4600 1955.5600 1747.9400 ;
        RECT 1953.9600 1742.0200 1955.5600 1742.5000 ;
        RECT 1953.9600 1736.5800 1955.5600 1737.0600 ;
        RECT 1953.9600 1731.1400 1955.5600 1731.6200 ;
        RECT 1953.9600 1725.7000 1955.5600 1726.1800 ;
        RECT 1953.9600 1720.2600 1955.5600 1720.7400 ;
        RECT 1953.9600 1714.8200 1955.5600 1715.3000 ;
        RECT 1953.9600 1709.3800 1955.5600 1709.8600 ;
        RECT 1953.9600 1703.9400 1955.5600 1704.4200 ;
        RECT 1953.9600 1698.5000 1955.5600 1698.9800 ;
        RECT 1953.9600 1693.0600 1955.5600 1693.5400 ;
        RECT 1953.9600 1687.6200 1955.5600 1688.1000 ;
        RECT 1953.9600 1682.1800 1955.5600 1682.6600 ;
        RECT 1953.9600 1676.7400 1955.5600 1677.2200 ;
        RECT 1953.9600 1671.3000 1955.5600 1671.7800 ;
        RECT 1953.9600 1665.8600 1955.5600 1666.3400 ;
        RECT 1953.9600 1660.4200 1955.5600 1660.9000 ;
        RECT 1953.9600 1654.9800 1955.5600 1655.4600 ;
        RECT 1953.9600 1649.5400 1955.5600 1650.0200 ;
        RECT 1953.9600 1644.1000 1955.5600 1644.5800 ;
        RECT 1953.9600 1638.6600 1955.5600 1639.1400 ;
        RECT 1953.9600 1633.2200 1955.5600 1633.7000 ;
        RECT 1953.9600 1627.7800 1955.5600 1628.2600 ;
        RECT 1953.9600 1622.3400 1955.5600 1622.8200 ;
        RECT 1953.9600 1611.4600 1955.5600 1611.9400 ;
        RECT 1953.9600 1606.0200 1955.5600 1606.5000 ;
        RECT 1953.9600 1600.5800 1955.5600 1601.0600 ;
        RECT 1953.9600 1595.1400 1955.5600 1595.6200 ;
        RECT 1953.9600 1589.7000 1955.5600 1590.1800 ;
        RECT 1953.9600 1584.2600 1955.5600 1584.7400 ;
        RECT 1953.9600 1578.8200 1955.5600 1579.3000 ;
        RECT 1953.9600 1573.3800 1955.5600 1573.8600 ;
        RECT 1953.9600 1616.9000 1955.5600 1617.3800 ;
        RECT 2156.6600 1785.5400 2158.2600 1786.0200 ;
        RECT 1953.9600 1785.5400 1955.5600 1786.0200 ;
        RECT 1951.0000 2006.2600 2161.2200 2007.8600 ;
        RECT 1951.0000 1563.8700 2161.2200 1565.4700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 1561.0400 1955.5600 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 2009.2600 1955.5600 2010.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 1561.0400 2158.2600 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 2009.2600 2158.2600 2010.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1563.8700 1952.6000 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1563.8700 2161.2200 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2006.2600 1952.6000 2007.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2006.2600 2161.2200 2007.8600 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1953.9600 1101.7600 1955.5600 1551.5800 ;
        RECT 2156.6600 1101.7600 2158.2600 1551.5800 ;
        RECT 1961.1200 1104.5900 1962.7200 1548.5800 ;
        RECT 2006.1200 1104.5900 2007.7200 1548.5800 ;
        RECT 2051.1200 1104.5900 2052.7200 1548.5800 ;
        RECT 2096.1200 1104.5900 2097.7200 1548.5800 ;
        RECT 2141.1200 1104.5900 2142.7200 1548.5800 ;
      LAYER met3 ;
        RECT 2156.6600 1538.4200 2158.2600 1538.9000 ;
        RECT 2156.6600 1532.9800 2158.2600 1533.4600 ;
        RECT 2156.6600 1527.5400 2158.2600 1528.0200 ;
        RECT 2156.6600 1522.1000 2158.2600 1522.5800 ;
        RECT 2156.6600 1516.6600 2158.2600 1517.1400 ;
        RECT 2156.6600 1511.2200 2158.2600 1511.7000 ;
        RECT 2156.6600 1505.7800 2158.2600 1506.2600 ;
        RECT 2156.6600 1500.3400 2158.2600 1500.8200 ;
        RECT 2156.6600 1489.4600 2158.2600 1489.9400 ;
        RECT 2156.6600 1484.0200 2158.2600 1484.5000 ;
        RECT 2156.6600 1478.5800 2158.2600 1479.0600 ;
        RECT 2156.6600 1473.1400 2158.2600 1473.6200 ;
        RECT 2156.6600 1467.7000 2158.2600 1468.1800 ;
        RECT 2156.6600 1462.2600 2158.2600 1462.7400 ;
        RECT 2156.6600 1456.8200 2158.2600 1457.3000 ;
        RECT 2156.6600 1451.3800 2158.2600 1451.8600 ;
        RECT 2156.6600 1445.9400 2158.2600 1446.4200 ;
        RECT 2156.6600 1440.5000 2158.2600 1440.9800 ;
        RECT 2156.6600 1494.9000 2158.2600 1495.3800 ;
        RECT 2156.6600 1435.0600 2158.2600 1435.5400 ;
        RECT 2156.6600 1429.6200 2158.2600 1430.1000 ;
        RECT 2156.6600 1424.1800 2158.2600 1424.6600 ;
        RECT 2156.6600 1418.7400 2158.2600 1419.2200 ;
        RECT 2156.6600 1413.3000 2158.2600 1413.7800 ;
        RECT 2156.6600 1407.8600 2158.2600 1408.3400 ;
        RECT 2156.6600 1402.4200 2158.2600 1402.9000 ;
        RECT 2156.6600 1396.9800 2158.2600 1397.4600 ;
        RECT 2156.6600 1391.5400 2158.2600 1392.0200 ;
        RECT 2156.6600 1386.1000 2158.2600 1386.5800 ;
        RECT 2156.6600 1380.6600 2158.2600 1381.1400 ;
        RECT 2156.6600 1375.2200 2158.2600 1375.7000 ;
        RECT 2156.6600 1369.7800 2158.2600 1370.2600 ;
        RECT 2156.6600 1364.3400 2158.2600 1364.8200 ;
        RECT 2156.6600 1358.9000 2158.2600 1359.3800 ;
        RECT 2156.6600 1353.4600 2158.2600 1353.9400 ;
        RECT 2156.6600 1348.0200 2158.2600 1348.5000 ;
        RECT 2156.6600 1342.5800 2158.2600 1343.0600 ;
        RECT 2156.6600 1337.1400 2158.2600 1337.6200 ;
        RECT 2156.6600 1331.7000 2158.2600 1332.1800 ;
        RECT 1953.9600 1538.4200 1955.5600 1538.9000 ;
        RECT 1953.9600 1532.9800 1955.5600 1533.4600 ;
        RECT 1953.9600 1527.5400 1955.5600 1528.0200 ;
        RECT 1953.9600 1522.1000 1955.5600 1522.5800 ;
        RECT 1953.9600 1516.6600 1955.5600 1517.1400 ;
        RECT 1953.9600 1511.2200 1955.5600 1511.7000 ;
        RECT 1953.9600 1505.7800 1955.5600 1506.2600 ;
        RECT 1953.9600 1500.3400 1955.5600 1500.8200 ;
        RECT 1953.9600 1489.4600 1955.5600 1489.9400 ;
        RECT 1953.9600 1484.0200 1955.5600 1484.5000 ;
        RECT 1953.9600 1478.5800 1955.5600 1479.0600 ;
        RECT 1953.9600 1473.1400 1955.5600 1473.6200 ;
        RECT 1953.9600 1467.7000 1955.5600 1468.1800 ;
        RECT 1953.9600 1462.2600 1955.5600 1462.7400 ;
        RECT 1953.9600 1456.8200 1955.5600 1457.3000 ;
        RECT 1953.9600 1451.3800 1955.5600 1451.8600 ;
        RECT 1953.9600 1445.9400 1955.5600 1446.4200 ;
        RECT 1953.9600 1440.5000 1955.5600 1440.9800 ;
        RECT 1953.9600 1494.9000 1955.5600 1495.3800 ;
        RECT 1953.9600 1435.0600 1955.5600 1435.5400 ;
        RECT 1953.9600 1429.6200 1955.5600 1430.1000 ;
        RECT 1953.9600 1424.1800 1955.5600 1424.6600 ;
        RECT 1953.9600 1418.7400 1955.5600 1419.2200 ;
        RECT 1953.9600 1413.3000 1955.5600 1413.7800 ;
        RECT 1953.9600 1407.8600 1955.5600 1408.3400 ;
        RECT 1953.9600 1402.4200 1955.5600 1402.9000 ;
        RECT 1953.9600 1396.9800 1955.5600 1397.4600 ;
        RECT 1953.9600 1391.5400 1955.5600 1392.0200 ;
        RECT 1953.9600 1386.1000 1955.5600 1386.5800 ;
        RECT 1953.9600 1380.6600 1955.5600 1381.1400 ;
        RECT 1953.9600 1375.2200 1955.5600 1375.7000 ;
        RECT 1953.9600 1369.7800 1955.5600 1370.2600 ;
        RECT 1953.9600 1364.3400 1955.5600 1364.8200 ;
        RECT 1953.9600 1358.9000 1955.5600 1359.3800 ;
        RECT 1953.9600 1353.4600 1955.5600 1353.9400 ;
        RECT 1953.9600 1348.0200 1955.5600 1348.5000 ;
        RECT 1953.9600 1342.5800 1955.5600 1343.0600 ;
        RECT 1953.9600 1337.1400 1955.5600 1337.6200 ;
        RECT 1953.9600 1331.7000 1955.5600 1332.1800 ;
        RECT 2156.6600 1320.8200 2158.2600 1321.3000 ;
        RECT 2156.6600 1315.3800 2158.2600 1315.8600 ;
        RECT 2156.6600 1309.9400 2158.2600 1310.4200 ;
        RECT 2156.6600 1304.5000 2158.2600 1304.9800 ;
        RECT 2156.6600 1299.0600 2158.2600 1299.5400 ;
        RECT 2156.6600 1293.6200 2158.2600 1294.1000 ;
        RECT 2156.6600 1288.1800 2158.2600 1288.6600 ;
        RECT 2156.6600 1282.7400 2158.2600 1283.2200 ;
        RECT 2156.6600 1277.3000 2158.2600 1277.7800 ;
        RECT 2156.6600 1271.8600 2158.2600 1272.3400 ;
        RECT 2156.6600 1266.4200 2158.2600 1266.9000 ;
        RECT 2156.6600 1260.9800 2158.2600 1261.4600 ;
        RECT 2156.6600 1255.5400 2158.2600 1256.0200 ;
        RECT 2156.6600 1250.1000 2158.2600 1250.5800 ;
        RECT 2156.6600 1244.6600 2158.2600 1245.1400 ;
        RECT 2156.6600 1239.2200 2158.2600 1239.7000 ;
        RECT 2156.6600 1233.7800 2158.2600 1234.2600 ;
        RECT 2156.6600 1228.3400 2158.2600 1228.8200 ;
        RECT 2156.6600 1222.9000 2158.2600 1223.3800 ;
        RECT 2156.6600 1217.4600 2158.2600 1217.9400 ;
        RECT 2156.6600 1212.0200 2158.2600 1212.5000 ;
        RECT 2156.6600 1206.5800 2158.2600 1207.0600 ;
        RECT 2156.6600 1201.1400 2158.2600 1201.6200 ;
        RECT 2156.6600 1195.7000 2158.2600 1196.1800 ;
        RECT 2156.6600 1190.2600 2158.2600 1190.7400 ;
        RECT 2156.6600 1184.8200 2158.2600 1185.3000 ;
        RECT 2156.6600 1179.3800 2158.2600 1179.8600 ;
        RECT 2156.6600 1173.9400 2158.2600 1174.4200 ;
        RECT 2156.6600 1168.5000 2158.2600 1168.9800 ;
        RECT 2156.6600 1163.0600 2158.2600 1163.5400 ;
        RECT 2156.6600 1152.1800 2158.2600 1152.6600 ;
        RECT 2156.6600 1146.7400 2158.2600 1147.2200 ;
        RECT 2156.6600 1141.3000 2158.2600 1141.7800 ;
        RECT 2156.6600 1135.8600 2158.2600 1136.3400 ;
        RECT 2156.6600 1130.4200 2158.2600 1130.9000 ;
        RECT 2156.6600 1124.9800 2158.2600 1125.4600 ;
        RECT 2156.6600 1119.5400 2158.2600 1120.0200 ;
        RECT 2156.6600 1114.1000 2158.2600 1114.5800 ;
        RECT 2156.6600 1157.6200 2158.2600 1158.1000 ;
        RECT 1953.9600 1320.8200 1955.5600 1321.3000 ;
        RECT 1953.9600 1315.3800 1955.5600 1315.8600 ;
        RECT 1953.9600 1309.9400 1955.5600 1310.4200 ;
        RECT 1953.9600 1304.5000 1955.5600 1304.9800 ;
        RECT 1953.9600 1299.0600 1955.5600 1299.5400 ;
        RECT 1953.9600 1293.6200 1955.5600 1294.1000 ;
        RECT 1953.9600 1288.1800 1955.5600 1288.6600 ;
        RECT 1953.9600 1282.7400 1955.5600 1283.2200 ;
        RECT 1953.9600 1277.3000 1955.5600 1277.7800 ;
        RECT 1953.9600 1271.8600 1955.5600 1272.3400 ;
        RECT 1953.9600 1266.4200 1955.5600 1266.9000 ;
        RECT 1953.9600 1260.9800 1955.5600 1261.4600 ;
        RECT 1953.9600 1255.5400 1955.5600 1256.0200 ;
        RECT 1953.9600 1250.1000 1955.5600 1250.5800 ;
        RECT 1953.9600 1244.6600 1955.5600 1245.1400 ;
        RECT 1953.9600 1239.2200 1955.5600 1239.7000 ;
        RECT 1953.9600 1233.7800 1955.5600 1234.2600 ;
        RECT 1953.9600 1228.3400 1955.5600 1228.8200 ;
        RECT 1953.9600 1222.9000 1955.5600 1223.3800 ;
        RECT 1953.9600 1217.4600 1955.5600 1217.9400 ;
        RECT 1953.9600 1212.0200 1955.5600 1212.5000 ;
        RECT 1953.9600 1206.5800 1955.5600 1207.0600 ;
        RECT 1953.9600 1201.1400 1955.5600 1201.6200 ;
        RECT 1953.9600 1195.7000 1955.5600 1196.1800 ;
        RECT 1953.9600 1190.2600 1955.5600 1190.7400 ;
        RECT 1953.9600 1184.8200 1955.5600 1185.3000 ;
        RECT 1953.9600 1179.3800 1955.5600 1179.8600 ;
        RECT 1953.9600 1173.9400 1955.5600 1174.4200 ;
        RECT 1953.9600 1168.5000 1955.5600 1168.9800 ;
        RECT 1953.9600 1163.0600 1955.5600 1163.5400 ;
        RECT 1953.9600 1152.1800 1955.5600 1152.6600 ;
        RECT 1953.9600 1146.7400 1955.5600 1147.2200 ;
        RECT 1953.9600 1141.3000 1955.5600 1141.7800 ;
        RECT 1953.9600 1135.8600 1955.5600 1136.3400 ;
        RECT 1953.9600 1130.4200 1955.5600 1130.9000 ;
        RECT 1953.9600 1124.9800 1955.5600 1125.4600 ;
        RECT 1953.9600 1119.5400 1955.5600 1120.0200 ;
        RECT 1953.9600 1114.1000 1955.5600 1114.5800 ;
        RECT 1953.9600 1157.6200 1955.5600 1158.1000 ;
        RECT 2156.6600 1326.2600 2158.2600 1326.7400 ;
        RECT 1953.9600 1326.2600 1955.5600 1326.7400 ;
        RECT 1951.0000 1546.9800 2161.2200 1548.5800 ;
        RECT 1951.0000 1104.5900 2161.2200 1106.1900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 1101.7600 1955.5600 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 1549.9800 1955.5600 1551.5800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 1101.7600 2158.2600 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 1549.9800 2158.2600 1551.5800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1104.5900 1952.6000 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1104.5900 2161.2200 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1546.9800 1952.6000 1548.5800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1546.9800 2161.2200 1548.5800 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1953.9600 642.4800 1955.5600 1092.3000 ;
        RECT 2156.6600 642.4800 2158.2600 1092.3000 ;
        RECT 1961.1200 645.3100 1962.7200 1089.3000 ;
        RECT 2006.1200 645.3100 2007.7200 1089.3000 ;
        RECT 2051.1200 645.3100 2052.7200 1089.3000 ;
        RECT 2096.1200 645.3100 2097.7200 1089.3000 ;
        RECT 2141.1200 645.3100 2142.7200 1089.3000 ;
      LAYER met3 ;
        RECT 2156.6600 1079.1400 2158.2600 1079.6200 ;
        RECT 2156.6600 1073.7000 2158.2600 1074.1800 ;
        RECT 2156.6600 1068.2600 2158.2600 1068.7400 ;
        RECT 2156.6600 1062.8200 2158.2600 1063.3000 ;
        RECT 2156.6600 1057.3800 2158.2600 1057.8600 ;
        RECT 2156.6600 1051.9400 2158.2600 1052.4200 ;
        RECT 2156.6600 1046.5000 2158.2600 1046.9800 ;
        RECT 2156.6600 1041.0600 2158.2600 1041.5400 ;
        RECT 2156.6600 1030.1800 2158.2600 1030.6600 ;
        RECT 2156.6600 1024.7400 2158.2600 1025.2200 ;
        RECT 2156.6600 1019.3000 2158.2600 1019.7800 ;
        RECT 2156.6600 1013.8600 2158.2600 1014.3400 ;
        RECT 2156.6600 1008.4200 2158.2600 1008.9000 ;
        RECT 2156.6600 1002.9800 2158.2600 1003.4600 ;
        RECT 2156.6600 997.5400 2158.2600 998.0200 ;
        RECT 2156.6600 992.1000 2158.2600 992.5800 ;
        RECT 2156.6600 986.6600 2158.2600 987.1400 ;
        RECT 2156.6600 981.2200 2158.2600 981.7000 ;
        RECT 2156.6600 1035.6200 2158.2600 1036.1000 ;
        RECT 2156.6600 975.7800 2158.2600 976.2600 ;
        RECT 2156.6600 970.3400 2158.2600 970.8200 ;
        RECT 2156.6600 964.9000 2158.2600 965.3800 ;
        RECT 2156.6600 959.4600 2158.2600 959.9400 ;
        RECT 2156.6600 954.0200 2158.2600 954.5000 ;
        RECT 2156.6600 948.5800 2158.2600 949.0600 ;
        RECT 2156.6600 943.1400 2158.2600 943.6200 ;
        RECT 2156.6600 937.7000 2158.2600 938.1800 ;
        RECT 2156.6600 932.2600 2158.2600 932.7400 ;
        RECT 2156.6600 926.8200 2158.2600 927.3000 ;
        RECT 2156.6600 921.3800 2158.2600 921.8600 ;
        RECT 2156.6600 915.9400 2158.2600 916.4200 ;
        RECT 2156.6600 910.5000 2158.2600 910.9800 ;
        RECT 2156.6600 905.0600 2158.2600 905.5400 ;
        RECT 2156.6600 899.6200 2158.2600 900.1000 ;
        RECT 2156.6600 894.1800 2158.2600 894.6600 ;
        RECT 2156.6600 888.7400 2158.2600 889.2200 ;
        RECT 2156.6600 883.3000 2158.2600 883.7800 ;
        RECT 2156.6600 877.8600 2158.2600 878.3400 ;
        RECT 2156.6600 872.4200 2158.2600 872.9000 ;
        RECT 1953.9600 1079.1400 1955.5600 1079.6200 ;
        RECT 1953.9600 1073.7000 1955.5600 1074.1800 ;
        RECT 1953.9600 1068.2600 1955.5600 1068.7400 ;
        RECT 1953.9600 1062.8200 1955.5600 1063.3000 ;
        RECT 1953.9600 1057.3800 1955.5600 1057.8600 ;
        RECT 1953.9600 1051.9400 1955.5600 1052.4200 ;
        RECT 1953.9600 1046.5000 1955.5600 1046.9800 ;
        RECT 1953.9600 1041.0600 1955.5600 1041.5400 ;
        RECT 1953.9600 1030.1800 1955.5600 1030.6600 ;
        RECT 1953.9600 1024.7400 1955.5600 1025.2200 ;
        RECT 1953.9600 1019.3000 1955.5600 1019.7800 ;
        RECT 1953.9600 1013.8600 1955.5600 1014.3400 ;
        RECT 1953.9600 1008.4200 1955.5600 1008.9000 ;
        RECT 1953.9600 1002.9800 1955.5600 1003.4600 ;
        RECT 1953.9600 997.5400 1955.5600 998.0200 ;
        RECT 1953.9600 992.1000 1955.5600 992.5800 ;
        RECT 1953.9600 986.6600 1955.5600 987.1400 ;
        RECT 1953.9600 981.2200 1955.5600 981.7000 ;
        RECT 1953.9600 1035.6200 1955.5600 1036.1000 ;
        RECT 1953.9600 975.7800 1955.5600 976.2600 ;
        RECT 1953.9600 970.3400 1955.5600 970.8200 ;
        RECT 1953.9600 964.9000 1955.5600 965.3800 ;
        RECT 1953.9600 959.4600 1955.5600 959.9400 ;
        RECT 1953.9600 954.0200 1955.5600 954.5000 ;
        RECT 1953.9600 948.5800 1955.5600 949.0600 ;
        RECT 1953.9600 943.1400 1955.5600 943.6200 ;
        RECT 1953.9600 937.7000 1955.5600 938.1800 ;
        RECT 1953.9600 932.2600 1955.5600 932.7400 ;
        RECT 1953.9600 926.8200 1955.5600 927.3000 ;
        RECT 1953.9600 921.3800 1955.5600 921.8600 ;
        RECT 1953.9600 915.9400 1955.5600 916.4200 ;
        RECT 1953.9600 910.5000 1955.5600 910.9800 ;
        RECT 1953.9600 905.0600 1955.5600 905.5400 ;
        RECT 1953.9600 899.6200 1955.5600 900.1000 ;
        RECT 1953.9600 894.1800 1955.5600 894.6600 ;
        RECT 1953.9600 888.7400 1955.5600 889.2200 ;
        RECT 1953.9600 883.3000 1955.5600 883.7800 ;
        RECT 1953.9600 877.8600 1955.5600 878.3400 ;
        RECT 1953.9600 872.4200 1955.5600 872.9000 ;
        RECT 2156.6600 861.5400 2158.2600 862.0200 ;
        RECT 2156.6600 856.1000 2158.2600 856.5800 ;
        RECT 2156.6600 850.6600 2158.2600 851.1400 ;
        RECT 2156.6600 845.2200 2158.2600 845.7000 ;
        RECT 2156.6600 839.7800 2158.2600 840.2600 ;
        RECT 2156.6600 834.3400 2158.2600 834.8200 ;
        RECT 2156.6600 828.9000 2158.2600 829.3800 ;
        RECT 2156.6600 823.4600 2158.2600 823.9400 ;
        RECT 2156.6600 818.0200 2158.2600 818.5000 ;
        RECT 2156.6600 812.5800 2158.2600 813.0600 ;
        RECT 2156.6600 807.1400 2158.2600 807.6200 ;
        RECT 2156.6600 801.7000 2158.2600 802.1800 ;
        RECT 2156.6600 796.2600 2158.2600 796.7400 ;
        RECT 2156.6600 790.8200 2158.2600 791.3000 ;
        RECT 2156.6600 785.3800 2158.2600 785.8600 ;
        RECT 2156.6600 779.9400 2158.2600 780.4200 ;
        RECT 2156.6600 774.5000 2158.2600 774.9800 ;
        RECT 2156.6600 769.0600 2158.2600 769.5400 ;
        RECT 2156.6600 763.6200 2158.2600 764.1000 ;
        RECT 2156.6600 758.1800 2158.2600 758.6600 ;
        RECT 2156.6600 752.7400 2158.2600 753.2200 ;
        RECT 2156.6600 747.3000 2158.2600 747.7800 ;
        RECT 2156.6600 741.8600 2158.2600 742.3400 ;
        RECT 2156.6600 736.4200 2158.2600 736.9000 ;
        RECT 2156.6600 730.9800 2158.2600 731.4600 ;
        RECT 2156.6600 725.5400 2158.2600 726.0200 ;
        RECT 2156.6600 720.1000 2158.2600 720.5800 ;
        RECT 2156.6600 714.6600 2158.2600 715.1400 ;
        RECT 2156.6600 709.2200 2158.2600 709.7000 ;
        RECT 2156.6600 703.7800 2158.2600 704.2600 ;
        RECT 2156.6600 692.9000 2158.2600 693.3800 ;
        RECT 2156.6600 687.4600 2158.2600 687.9400 ;
        RECT 2156.6600 682.0200 2158.2600 682.5000 ;
        RECT 2156.6600 676.5800 2158.2600 677.0600 ;
        RECT 2156.6600 671.1400 2158.2600 671.6200 ;
        RECT 2156.6600 665.7000 2158.2600 666.1800 ;
        RECT 2156.6600 660.2600 2158.2600 660.7400 ;
        RECT 2156.6600 654.8200 2158.2600 655.3000 ;
        RECT 2156.6600 698.3400 2158.2600 698.8200 ;
        RECT 1953.9600 861.5400 1955.5600 862.0200 ;
        RECT 1953.9600 856.1000 1955.5600 856.5800 ;
        RECT 1953.9600 850.6600 1955.5600 851.1400 ;
        RECT 1953.9600 845.2200 1955.5600 845.7000 ;
        RECT 1953.9600 839.7800 1955.5600 840.2600 ;
        RECT 1953.9600 834.3400 1955.5600 834.8200 ;
        RECT 1953.9600 828.9000 1955.5600 829.3800 ;
        RECT 1953.9600 823.4600 1955.5600 823.9400 ;
        RECT 1953.9600 818.0200 1955.5600 818.5000 ;
        RECT 1953.9600 812.5800 1955.5600 813.0600 ;
        RECT 1953.9600 807.1400 1955.5600 807.6200 ;
        RECT 1953.9600 801.7000 1955.5600 802.1800 ;
        RECT 1953.9600 796.2600 1955.5600 796.7400 ;
        RECT 1953.9600 790.8200 1955.5600 791.3000 ;
        RECT 1953.9600 785.3800 1955.5600 785.8600 ;
        RECT 1953.9600 779.9400 1955.5600 780.4200 ;
        RECT 1953.9600 774.5000 1955.5600 774.9800 ;
        RECT 1953.9600 769.0600 1955.5600 769.5400 ;
        RECT 1953.9600 763.6200 1955.5600 764.1000 ;
        RECT 1953.9600 758.1800 1955.5600 758.6600 ;
        RECT 1953.9600 752.7400 1955.5600 753.2200 ;
        RECT 1953.9600 747.3000 1955.5600 747.7800 ;
        RECT 1953.9600 741.8600 1955.5600 742.3400 ;
        RECT 1953.9600 736.4200 1955.5600 736.9000 ;
        RECT 1953.9600 730.9800 1955.5600 731.4600 ;
        RECT 1953.9600 725.5400 1955.5600 726.0200 ;
        RECT 1953.9600 720.1000 1955.5600 720.5800 ;
        RECT 1953.9600 714.6600 1955.5600 715.1400 ;
        RECT 1953.9600 709.2200 1955.5600 709.7000 ;
        RECT 1953.9600 703.7800 1955.5600 704.2600 ;
        RECT 1953.9600 692.9000 1955.5600 693.3800 ;
        RECT 1953.9600 687.4600 1955.5600 687.9400 ;
        RECT 1953.9600 682.0200 1955.5600 682.5000 ;
        RECT 1953.9600 676.5800 1955.5600 677.0600 ;
        RECT 1953.9600 671.1400 1955.5600 671.6200 ;
        RECT 1953.9600 665.7000 1955.5600 666.1800 ;
        RECT 1953.9600 660.2600 1955.5600 660.7400 ;
        RECT 1953.9600 654.8200 1955.5600 655.3000 ;
        RECT 1953.9600 698.3400 1955.5600 698.8200 ;
        RECT 2156.6600 866.9800 2158.2600 867.4600 ;
        RECT 1953.9600 866.9800 1955.5600 867.4600 ;
        RECT 1951.0000 1087.7000 2161.2200 1089.3000 ;
        RECT 1951.0000 645.3100 2161.2200 646.9100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 642.4800 1955.5600 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 1090.7000 1955.5600 1092.3000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 642.4800 2158.2600 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 1090.7000 2158.2600 1092.3000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 645.3100 1952.6000 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 645.3100 2161.2200 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1087.7000 1952.6000 1089.3000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1087.7000 2161.2200 1089.3000 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1953.9600 183.2000 1955.5600 633.0200 ;
        RECT 2156.6600 183.2000 2158.2600 633.0200 ;
        RECT 1961.1200 186.0300 1962.7200 630.0200 ;
        RECT 2006.1200 186.0300 2007.7200 630.0200 ;
        RECT 2051.1200 186.0300 2052.7200 630.0200 ;
        RECT 2096.1200 186.0300 2097.7200 630.0200 ;
        RECT 2141.1200 186.0300 2142.7200 630.0200 ;
      LAYER met3 ;
        RECT 2156.6600 619.8600 2158.2600 620.3400 ;
        RECT 2156.6600 614.4200 2158.2600 614.9000 ;
        RECT 2156.6600 608.9800 2158.2600 609.4600 ;
        RECT 2156.6600 603.5400 2158.2600 604.0200 ;
        RECT 2156.6600 598.1000 2158.2600 598.5800 ;
        RECT 2156.6600 592.6600 2158.2600 593.1400 ;
        RECT 2156.6600 587.2200 2158.2600 587.7000 ;
        RECT 2156.6600 581.7800 2158.2600 582.2600 ;
        RECT 2156.6600 570.9000 2158.2600 571.3800 ;
        RECT 2156.6600 565.4600 2158.2600 565.9400 ;
        RECT 2156.6600 560.0200 2158.2600 560.5000 ;
        RECT 2156.6600 554.5800 2158.2600 555.0600 ;
        RECT 2156.6600 549.1400 2158.2600 549.6200 ;
        RECT 2156.6600 543.7000 2158.2600 544.1800 ;
        RECT 2156.6600 538.2600 2158.2600 538.7400 ;
        RECT 2156.6600 532.8200 2158.2600 533.3000 ;
        RECT 2156.6600 527.3800 2158.2600 527.8600 ;
        RECT 2156.6600 521.9400 2158.2600 522.4200 ;
        RECT 2156.6600 576.3400 2158.2600 576.8200 ;
        RECT 2156.6600 516.5000 2158.2600 516.9800 ;
        RECT 2156.6600 511.0600 2158.2600 511.5400 ;
        RECT 2156.6600 505.6200 2158.2600 506.1000 ;
        RECT 2156.6600 500.1800 2158.2600 500.6600 ;
        RECT 2156.6600 494.7400 2158.2600 495.2200 ;
        RECT 2156.6600 489.3000 2158.2600 489.7800 ;
        RECT 2156.6600 483.8600 2158.2600 484.3400 ;
        RECT 2156.6600 478.4200 2158.2600 478.9000 ;
        RECT 2156.6600 472.9800 2158.2600 473.4600 ;
        RECT 2156.6600 467.5400 2158.2600 468.0200 ;
        RECT 2156.6600 462.1000 2158.2600 462.5800 ;
        RECT 2156.6600 456.6600 2158.2600 457.1400 ;
        RECT 2156.6600 451.2200 2158.2600 451.7000 ;
        RECT 2156.6600 445.7800 2158.2600 446.2600 ;
        RECT 2156.6600 440.3400 2158.2600 440.8200 ;
        RECT 2156.6600 434.9000 2158.2600 435.3800 ;
        RECT 2156.6600 429.4600 2158.2600 429.9400 ;
        RECT 2156.6600 424.0200 2158.2600 424.5000 ;
        RECT 2156.6600 418.5800 2158.2600 419.0600 ;
        RECT 2156.6600 413.1400 2158.2600 413.6200 ;
        RECT 1953.9600 619.8600 1955.5600 620.3400 ;
        RECT 1953.9600 614.4200 1955.5600 614.9000 ;
        RECT 1953.9600 608.9800 1955.5600 609.4600 ;
        RECT 1953.9600 603.5400 1955.5600 604.0200 ;
        RECT 1953.9600 598.1000 1955.5600 598.5800 ;
        RECT 1953.9600 592.6600 1955.5600 593.1400 ;
        RECT 1953.9600 587.2200 1955.5600 587.7000 ;
        RECT 1953.9600 581.7800 1955.5600 582.2600 ;
        RECT 1953.9600 570.9000 1955.5600 571.3800 ;
        RECT 1953.9600 565.4600 1955.5600 565.9400 ;
        RECT 1953.9600 560.0200 1955.5600 560.5000 ;
        RECT 1953.9600 554.5800 1955.5600 555.0600 ;
        RECT 1953.9600 549.1400 1955.5600 549.6200 ;
        RECT 1953.9600 543.7000 1955.5600 544.1800 ;
        RECT 1953.9600 538.2600 1955.5600 538.7400 ;
        RECT 1953.9600 532.8200 1955.5600 533.3000 ;
        RECT 1953.9600 527.3800 1955.5600 527.8600 ;
        RECT 1953.9600 521.9400 1955.5600 522.4200 ;
        RECT 1953.9600 576.3400 1955.5600 576.8200 ;
        RECT 1953.9600 516.5000 1955.5600 516.9800 ;
        RECT 1953.9600 511.0600 1955.5600 511.5400 ;
        RECT 1953.9600 505.6200 1955.5600 506.1000 ;
        RECT 1953.9600 500.1800 1955.5600 500.6600 ;
        RECT 1953.9600 494.7400 1955.5600 495.2200 ;
        RECT 1953.9600 489.3000 1955.5600 489.7800 ;
        RECT 1953.9600 483.8600 1955.5600 484.3400 ;
        RECT 1953.9600 478.4200 1955.5600 478.9000 ;
        RECT 1953.9600 472.9800 1955.5600 473.4600 ;
        RECT 1953.9600 467.5400 1955.5600 468.0200 ;
        RECT 1953.9600 462.1000 1955.5600 462.5800 ;
        RECT 1953.9600 456.6600 1955.5600 457.1400 ;
        RECT 1953.9600 451.2200 1955.5600 451.7000 ;
        RECT 1953.9600 445.7800 1955.5600 446.2600 ;
        RECT 1953.9600 440.3400 1955.5600 440.8200 ;
        RECT 1953.9600 434.9000 1955.5600 435.3800 ;
        RECT 1953.9600 429.4600 1955.5600 429.9400 ;
        RECT 1953.9600 424.0200 1955.5600 424.5000 ;
        RECT 1953.9600 418.5800 1955.5600 419.0600 ;
        RECT 1953.9600 413.1400 1955.5600 413.6200 ;
        RECT 2156.6600 402.2600 2158.2600 402.7400 ;
        RECT 2156.6600 396.8200 2158.2600 397.3000 ;
        RECT 2156.6600 391.3800 2158.2600 391.8600 ;
        RECT 2156.6600 385.9400 2158.2600 386.4200 ;
        RECT 2156.6600 380.5000 2158.2600 380.9800 ;
        RECT 2156.6600 375.0600 2158.2600 375.5400 ;
        RECT 2156.6600 369.6200 2158.2600 370.1000 ;
        RECT 2156.6600 364.1800 2158.2600 364.6600 ;
        RECT 2156.6600 358.7400 2158.2600 359.2200 ;
        RECT 2156.6600 353.3000 2158.2600 353.7800 ;
        RECT 2156.6600 347.8600 2158.2600 348.3400 ;
        RECT 2156.6600 342.4200 2158.2600 342.9000 ;
        RECT 2156.6600 336.9800 2158.2600 337.4600 ;
        RECT 2156.6600 331.5400 2158.2600 332.0200 ;
        RECT 2156.6600 326.1000 2158.2600 326.5800 ;
        RECT 2156.6600 320.6600 2158.2600 321.1400 ;
        RECT 2156.6600 315.2200 2158.2600 315.7000 ;
        RECT 2156.6600 309.7800 2158.2600 310.2600 ;
        RECT 2156.6600 304.3400 2158.2600 304.8200 ;
        RECT 2156.6600 298.9000 2158.2600 299.3800 ;
        RECT 2156.6600 293.4600 2158.2600 293.9400 ;
        RECT 2156.6600 288.0200 2158.2600 288.5000 ;
        RECT 2156.6600 282.5800 2158.2600 283.0600 ;
        RECT 2156.6600 277.1400 2158.2600 277.6200 ;
        RECT 2156.6600 271.7000 2158.2600 272.1800 ;
        RECT 2156.6600 266.2600 2158.2600 266.7400 ;
        RECT 2156.6600 260.8200 2158.2600 261.3000 ;
        RECT 2156.6600 255.3800 2158.2600 255.8600 ;
        RECT 2156.6600 249.9400 2158.2600 250.4200 ;
        RECT 2156.6600 244.5000 2158.2600 244.9800 ;
        RECT 2156.6600 233.6200 2158.2600 234.1000 ;
        RECT 2156.6600 228.1800 2158.2600 228.6600 ;
        RECT 2156.6600 222.7400 2158.2600 223.2200 ;
        RECT 2156.6600 217.3000 2158.2600 217.7800 ;
        RECT 2156.6600 211.8600 2158.2600 212.3400 ;
        RECT 2156.6600 206.4200 2158.2600 206.9000 ;
        RECT 2156.6600 200.9800 2158.2600 201.4600 ;
        RECT 2156.6600 195.5400 2158.2600 196.0200 ;
        RECT 2156.6600 239.0600 2158.2600 239.5400 ;
        RECT 1953.9600 402.2600 1955.5600 402.7400 ;
        RECT 1953.9600 396.8200 1955.5600 397.3000 ;
        RECT 1953.9600 391.3800 1955.5600 391.8600 ;
        RECT 1953.9600 385.9400 1955.5600 386.4200 ;
        RECT 1953.9600 380.5000 1955.5600 380.9800 ;
        RECT 1953.9600 375.0600 1955.5600 375.5400 ;
        RECT 1953.9600 369.6200 1955.5600 370.1000 ;
        RECT 1953.9600 364.1800 1955.5600 364.6600 ;
        RECT 1953.9600 358.7400 1955.5600 359.2200 ;
        RECT 1953.9600 353.3000 1955.5600 353.7800 ;
        RECT 1953.9600 347.8600 1955.5600 348.3400 ;
        RECT 1953.9600 342.4200 1955.5600 342.9000 ;
        RECT 1953.9600 336.9800 1955.5600 337.4600 ;
        RECT 1953.9600 331.5400 1955.5600 332.0200 ;
        RECT 1953.9600 326.1000 1955.5600 326.5800 ;
        RECT 1953.9600 320.6600 1955.5600 321.1400 ;
        RECT 1953.9600 315.2200 1955.5600 315.7000 ;
        RECT 1953.9600 309.7800 1955.5600 310.2600 ;
        RECT 1953.9600 304.3400 1955.5600 304.8200 ;
        RECT 1953.9600 298.9000 1955.5600 299.3800 ;
        RECT 1953.9600 293.4600 1955.5600 293.9400 ;
        RECT 1953.9600 288.0200 1955.5600 288.5000 ;
        RECT 1953.9600 282.5800 1955.5600 283.0600 ;
        RECT 1953.9600 277.1400 1955.5600 277.6200 ;
        RECT 1953.9600 271.7000 1955.5600 272.1800 ;
        RECT 1953.9600 266.2600 1955.5600 266.7400 ;
        RECT 1953.9600 260.8200 1955.5600 261.3000 ;
        RECT 1953.9600 255.3800 1955.5600 255.8600 ;
        RECT 1953.9600 249.9400 1955.5600 250.4200 ;
        RECT 1953.9600 244.5000 1955.5600 244.9800 ;
        RECT 1953.9600 233.6200 1955.5600 234.1000 ;
        RECT 1953.9600 228.1800 1955.5600 228.6600 ;
        RECT 1953.9600 222.7400 1955.5600 223.2200 ;
        RECT 1953.9600 217.3000 1955.5600 217.7800 ;
        RECT 1953.9600 211.8600 1955.5600 212.3400 ;
        RECT 1953.9600 206.4200 1955.5600 206.9000 ;
        RECT 1953.9600 200.9800 1955.5600 201.4600 ;
        RECT 1953.9600 195.5400 1955.5600 196.0200 ;
        RECT 1953.9600 239.0600 1955.5600 239.5400 ;
        RECT 2156.6600 407.7000 2158.2600 408.1800 ;
        RECT 1953.9600 407.7000 1955.5600 408.1800 ;
        RECT 1951.0000 628.4200 2161.2200 630.0200 ;
        RECT 1951.0000 186.0300 2161.2200 187.6300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 183.2000 1955.5600 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1953.9600 631.4200 1955.5600 633.0200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 183.2000 2158.2600 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2156.6600 631.4200 2158.2600 633.0200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 186.0300 1952.6000 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 186.0300 2161.2200 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 628.4200 1952.6000 630.0200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 628.4200 2161.2200 630.0200 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2174.2800 2479.6000 2175.8800 2509.8600 ;
        RECT 2376.7800 2479.6000 2378.3800 2509.8600 ;
      LAYER met3 ;
        RECT 2376.7800 2500.1000 2378.3800 2500.5800 ;
        RECT 2174.2800 2500.1000 2175.8800 2500.5800 ;
        RECT 2376.7800 2489.2200 2378.3800 2489.7000 ;
        RECT 2174.2800 2489.2200 2175.8800 2489.7000 ;
        RECT 2376.7800 2494.6600 2378.3800 2495.1400 ;
        RECT 2174.2800 2494.6600 2175.8800 2495.1400 ;
        RECT 2171.2200 2505.5000 2381.4400 2507.1000 ;
        RECT 2171.2200 2481.1700 2381.4400 2482.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.2800 2479.6000 2175.8800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.2800 2508.2600 2175.8800 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.7800 2479.6000 2378.3800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.7800 2508.2600 2378.3800 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2481.1700 2172.8200 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2481.1700 2381.4400 2482.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2505.5000 2172.8200 2507.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2505.5000 2381.4400 2507.1000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 186.0300 2362.9400 399.3300 ;
        RECT 2316.3400 186.0300 2317.9400 399.3300 ;
        RECT 2271.3400 186.0300 2272.9400 399.3300 ;
        RECT 2226.3400 186.0300 2227.9400 399.3300 ;
        RECT 2181.3400 186.0300 2182.9400 399.3300 ;
        RECT 2376.8800 183.2000 2378.4800 402.8400 ;
        RECT 2174.1800 183.2000 2175.7800 402.8400 ;
      LAYER met3 ;
        RECT 2361.3400 391.3800 2362.9400 391.8600 ;
        RECT 2376.8800 391.3800 2378.4800 391.8600 ;
        RECT 2376.8800 380.5000 2378.4800 380.9800 ;
        RECT 2376.8800 385.9400 2378.4800 386.4200 ;
        RECT 2361.3400 380.5000 2362.9400 380.9800 ;
        RECT 2361.3400 385.9400 2362.9400 386.4200 ;
        RECT 2376.8800 364.1800 2378.4800 364.6600 ;
        RECT 2376.8800 369.6200 2378.4800 370.1000 ;
        RECT 2361.3400 364.1800 2362.9400 364.6600 ;
        RECT 2361.3400 369.6200 2362.9400 370.1000 ;
        RECT 2376.8800 353.3000 2378.4800 353.7800 ;
        RECT 2376.8800 358.7400 2378.4800 359.2200 ;
        RECT 2361.3400 353.3000 2362.9400 353.7800 ;
        RECT 2361.3400 358.7400 2362.9400 359.2200 ;
        RECT 2361.3400 375.0600 2362.9400 375.5400 ;
        RECT 2376.8800 375.0600 2378.4800 375.5400 ;
        RECT 2316.3400 380.5000 2317.9400 380.9800 ;
        RECT 2316.3400 385.9400 2317.9400 386.4200 ;
        RECT 2316.3400 391.3800 2317.9400 391.8600 ;
        RECT 2316.3400 364.1800 2317.9400 364.6600 ;
        RECT 2316.3400 369.6200 2317.9400 370.1000 ;
        RECT 2316.3400 358.7400 2317.9400 359.2200 ;
        RECT 2316.3400 353.3000 2317.9400 353.7800 ;
        RECT 2316.3400 375.0600 2317.9400 375.5400 ;
        RECT 2376.8800 336.9800 2378.4800 337.4600 ;
        RECT 2376.8800 342.4200 2378.4800 342.9000 ;
        RECT 2361.3400 336.9800 2362.9400 337.4600 ;
        RECT 2361.3400 342.4200 2362.9400 342.9000 ;
        RECT 2376.8800 320.6600 2378.4800 321.1400 ;
        RECT 2376.8800 326.1000 2378.4800 326.5800 ;
        RECT 2376.8800 331.5400 2378.4800 332.0200 ;
        RECT 2361.3400 320.6600 2362.9400 321.1400 ;
        RECT 2361.3400 326.1000 2362.9400 326.5800 ;
        RECT 2361.3400 331.5400 2362.9400 332.0200 ;
        RECT 2376.8800 309.7800 2378.4800 310.2600 ;
        RECT 2376.8800 315.2200 2378.4800 315.7000 ;
        RECT 2361.3400 309.7800 2362.9400 310.2600 ;
        RECT 2361.3400 315.2200 2362.9400 315.7000 ;
        RECT 2376.8800 293.4600 2378.4800 293.9400 ;
        RECT 2376.8800 298.9000 2378.4800 299.3800 ;
        RECT 2376.8800 304.3400 2378.4800 304.8200 ;
        RECT 2361.3400 293.4600 2362.9400 293.9400 ;
        RECT 2361.3400 298.9000 2362.9400 299.3800 ;
        RECT 2361.3400 304.3400 2362.9400 304.8200 ;
        RECT 2316.3400 336.9800 2317.9400 337.4600 ;
        RECT 2316.3400 342.4200 2317.9400 342.9000 ;
        RECT 2316.3400 320.6600 2317.9400 321.1400 ;
        RECT 2316.3400 326.1000 2317.9400 326.5800 ;
        RECT 2316.3400 331.5400 2317.9400 332.0200 ;
        RECT 2316.3400 309.7800 2317.9400 310.2600 ;
        RECT 2316.3400 315.2200 2317.9400 315.7000 ;
        RECT 2316.3400 293.4600 2317.9400 293.9400 ;
        RECT 2316.3400 298.9000 2317.9400 299.3800 ;
        RECT 2316.3400 304.3400 2317.9400 304.8200 ;
        RECT 2316.3400 347.8600 2317.9400 348.3400 ;
        RECT 2361.3400 347.8600 2362.9400 348.3400 ;
        RECT 2376.8800 347.8600 2378.4800 348.3400 ;
        RECT 2271.3400 380.5000 2272.9400 380.9800 ;
        RECT 2271.3400 385.9400 2272.9400 386.4200 ;
        RECT 2271.3400 391.3800 2272.9400 391.8600 ;
        RECT 2226.3400 380.5000 2227.9400 380.9800 ;
        RECT 2226.3400 385.9400 2227.9400 386.4200 ;
        RECT 2226.3400 391.3800 2227.9400 391.8600 ;
        RECT 2271.3400 364.1800 2272.9400 364.6600 ;
        RECT 2271.3400 369.6200 2272.9400 370.1000 ;
        RECT 2271.3400 353.3000 2272.9400 353.7800 ;
        RECT 2271.3400 358.7400 2272.9400 359.2200 ;
        RECT 2226.3400 364.1800 2227.9400 364.6600 ;
        RECT 2226.3400 369.6200 2227.9400 370.1000 ;
        RECT 2226.3400 353.3000 2227.9400 353.7800 ;
        RECT 2226.3400 358.7400 2227.9400 359.2200 ;
        RECT 2226.3400 375.0600 2227.9400 375.5400 ;
        RECT 2271.3400 375.0600 2272.9400 375.5400 ;
        RECT 2174.1800 391.3800 2175.7800 391.8600 ;
        RECT 2181.3400 391.3800 2182.9400 391.8600 ;
        RECT 2181.3400 380.5000 2182.9400 380.9800 ;
        RECT 2181.3400 385.9400 2182.9400 386.4200 ;
        RECT 2174.1800 380.5000 2175.7800 380.9800 ;
        RECT 2174.1800 385.9400 2175.7800 386.4200 ;
        RECT 2181.3400 364.1800 2182.9400 364.6600 ;
        RECT 2181.3400 369.6200 2182.9400 370.1000 ;
        RECT 2174.1800 364.1800 2175.7800 364.6600 ;
        RECT 2174.1800 369.6200 2175.7800 370.1000 ;
        RECT 2181.3400 353.3000 2182.9400 353.7800 ;
        RECT 2181.3400 358.7400 2182.9400 359.2200 ;
        RECT 2174.1800 353.3000 2175.7800 353.7800 ;
        RECT 2174.1800 358.7400 2175.7800 359.2200 ;
        RECT 2174.1800 375.0600 2175.7800 375.5400 ;
        RECT 2181.3400 375.0600 2182.9400 375.5400 ;
        RECT 2271.3400 336.9800 2272.9400 337.4600 ;
        RECT 2271.3400 342.4200 2272.9400 342.9000 ;
        RECT 2271.3400 320.6600 2272.9400 321.1400 ;
        RECT 2271.3400 326.1000 2272.9400 326.5800 ;
        RECT 2271.3400 331.5400 2272.9400 332.0200 ;
        RECT 2226.3400 336.9800 2227.9400 337.4600 ;
        RECT 2226.3400 342.4200 2227.9400 342.9000 ;
        RECT 2226.3400 320.6600 2227.9400 321.1400 ;
        RECT 2226.3400 326.1000 2227.9400 326.5800 ;
        RECT 2226.3400 331.5400 2227.9400 332.0200 ;
        RECT 2271.3400 309.7800 2272.9400 310.2600 ;
        RECT 2271.3400 315.2200 2272.9400 315.7000 ;
        RECT 2271.3400 293.4600 2272.9400 293.9400 ;
        RECT 2271.3400 298.9000 2272.9400 299.3800 ;
        RECT 2271.3400 304.3400 2272.9400 304.8200 ;
        RECT 2226.3400 309.7800 2227.9400 310.2600 ;
        RECT 2226.3400 315.2200 2227.9400 315.7000 ;
        RECT 2226.3400 293.4600 2227.9400 293.9400 ;
        RECT 2226.3400 298.9000 2227.9400 299.3800 ;
        RECT 2226.3400 304.3400 2227.9400 304.8200 ;
        RECT 2181.3400 336.9800 2182.9400 337.4600 ;
        RECT 2181.3400 342.4200 2182.9400 342.9000 ;
        RECT 2174.1800 336.9800 2175.7800 337.4600 ;
        RECT 2174.1800 342.4200 2175.7800 342.9000 ;
        RECT 2181.3400 320.6600 2182.9400 321.1400 ;
        RECT 2181.3400 326.1000 2182.9400 326.5800 ;
        RECT 2181.3400 331.5400 2182.9400 332.0200 ;
        RECT 2174.1800 320.6600 2175.7800 321.1400 ;
        RECT 2174.1800 326.1000 2175.7800 326.5800 ;
        RECT 2174.1800 331.5400 2175.7800 332.0200 ;
        RECT 2181.3400 309.7800 2182.9400 310.2600 ;
        RECT 2181.3400 315.2200 2182.9400 315.7000 ;
        RECT 2174.1800 309.7800 2175.7800 310.2600 ;
        RECT 2174.1800 315.2200 2175.7800 315.7000 ;
        RECT 2181.3400 293.4600 2182.9400 293.9400 ;
        RECT 2181.3400 298.9000 2182.9400 299.3800 ;
        RECT 2181.3400 304.3400 2182.9400 304.8200 ;
        RECT 2174.1800 293.4600 2175.7800 293.9400 ;
        RECT 2174.1800 298.9000 2175.7800 299.3800 ;
        RECT 2174.1800 304.3400 2175.7800 304.8200 ;
        RECT 2174.1800 347.8600 2175.7800 348.3400 ;
        RECT 2181.3400 347.8600 2182.9400 348.3400 ;
        RECT 2226.3400 347.8600 2227.9400 348.3400 ;
        RECT 2271.3400 347.8600 2272.9400 348.3400 ;
        RECT 2376.8800 282.5800 2378.4800 283.0600 ;
        RECT 2376.8800 288.0200 2378.4800 288.5000 ;
        RECT 2361.3400 282.5800 2362.9400 283.0600 ;
        RECT 2361.3400 288.0200 2362.9400 288.5000 ;
        RECT 2376.8800 266.2600 2378.4800 266.7400 ;
        RECT 2376.8800 271.7000 2378.4800 272.1800 ;
        RECT 2376.8800 277.1400 2378.4800 277.6200 ;
        RECT 2361.3400 266.2600 2362.9400 266.7400 ;
        RECT 2361.3400 271.7000 2362.9400 272.1800 ;
        RECT 2361.3400 277.1400 2362.9400 277.6200 ;
        RECT 2376.8800 255.3800 2378.4800 255.8600 ;
        RECT 2376.8800 260.8200 2378.4800 261.3000 ;
        RECT 2361.3400 255.3800 2362.9400 255.8600 ;
        RECT 2361.3400 260.8200 2362.9400 261.3000 ;
        RECT 2376.8800 239.0600 2378.4800 239.5400 ;
        RECT 2376.8800 244.5000 2378.4800 244.9800 ;
        RECT 2376.8800 249.9400 2378.4800 250.4200 ;
        RECT 2361.3400 239.0600 2362.9400 239.5400 ;
        RECT 2361.3400 244.5000 2362.9400 244.9800 ;
        RECT 2361.3400 249.9400 2362.9400 250.4200 ;
        RECT 2316.3400 282.5800 2317.9400 283.0600 ;
        RECT 2316.3400 288.0200 2317.9400 288.5000 ;
        RECT 2316.3400 266.2600 2317.9400 266.7400 ;
        RECT 2316.3400 271.7000 2317.9400 272.1800 ;
        RECT 2316.3400 277.1400 2317.9400 277.6200 ;
        RECT 2316.3400 255.3800 2317.9400 255.8600 ;
        RECT 2316.3400 260.8200 2317.9400 261.3000 ;
        RECT 2316.3400 239.0600 2317.9400 239.5400 ;
        RECT 2316.3400 244.5000 2317.9400 244.9800 ;
        RECT 2316.3400 249.9400 2317.9400 250.4200 ;
        RECT 2376.8800 228.1800 2378.4800 228.6600 ;
        RECT 2376.8800 233.6200 2378.4800 234.1000 ;
        RECT 2361.3400 228.1800 2362.9400 228.6600 ;
        RECT 2361.3400 233.6200 2362.9400 234.1000 ;
        RECT 2376.8800 211.8600 2378.4800 212.3400 ;
        RECT 2376.8800 217.3000 2378.4800 217.7800 ;
        RECT 2376.8800 222.7400 2378.4800 223.2200 ;
        RECT 2361.3400 211.8600 2362.9400 212.3400 ;
        RECT 2361.3400 217.3000 2362.9400 217.7800 ;
        RECT 2361.3400 222.7400 2362.9400 223.2200 ;
        RECT 2376.8800 200.9800 2378.4800 201.4600 ;
        RECT 2376.8800 206.4200 2378.4800 206.9000 ;
        RECT 2361.3400 200.9800 2362.9400 201.4600 ;
        RECT 2361.3400 206.4200 2362.9400 206.9000 ;
        RECT 2361.3400 195.5400 2362.9400 196.0200 ;
        RECT 2376.8800 195.5400 2378.4800 196.0200 ;
        RECT 2316.3400 228.1800 2317.9400 228.6600 ;
        RECT 2316.3400 233.6200 2317.9400 234.1000 ;
        RECT 2316.3400 211.8600 2317.9400 212.3400 ;
        RECT 2316.3400 217.3000 2317.9400 217.7800 ;
        RECT 2316.3400 222.7400 2317.9400 223.2200 ;
        RECT 2316.3400 200.9800 2317.9400 201.4600 ;
        RECT 2316.3400 206.4200 2317.9400 206.9000 ;
        RECT 2316.3400 195.5400 2317.9400 196.0200 ;
        RECT 2271.3400 282.5800 2272.9400 283.0600 ;
        RECT 2271.3400 288.0200 2272.9400 288.5000 ;
        RECT 2271.3400 266.2600 2272.9400 266.7400 ;
        RECT 2271.3400 271.7000 2272.9400 272.1800 ;
        RECT 2271.3400 277.1400 2272.9400 277.6200 ;
        RECT 2226.3400 282.5800 2227.9400 283.0600 ;
        RECT 2226.3400 288.0200 2227.9400 288.5000 ;
        RECT 2226.3400 266.2600 2227.9400 266.7400 ;
        RECT 2226.3400 271.7000 2227.9400 272.1800 ;
        RECT 2226.3400 277.1400 2227.9400 277.6200 ;
        RECT 2271.3400 255.3800 2272.9400 255.8600 ;
        RECT 2271.3400 260.8200 2272.9400 261.3000 ;
        RECT 2271.3400 239.0600 2272.9400 239.5400 ;
        RECT 2271.3400 244.5000 2272.9400 244.9800 ;
        RECT 2271.3400 249.9400 2272.9400 250.4200 ;
        RECT 2226.3400 255.3800 2227.9400 255.8600 ;
        RECT 2226.3400 260.8200 2227.9400 261.3000 ;
        RECT 2226.3400 239.0600 2227.9400 239.5400 ;
        RECT 2226.3400 244.5000 2227.9400 244.9800 ;
        RECT 2226.3400 249.9400 2227.9400 250.4200 ;
        RECT 2181.3400 282.5800 2182.9400 283.0600 ;
        RECT 2181.3400 288.0200 2182.9400 288.5000 ;
        RECT 2174.1800 282.5800 2175.7800 283.0600 ;
        RECT 2174.1800 288.0200 2175.7800 288.5000 ;
        RECT 2181.3400 266.2600 2182.9400 266.7400 ;
        RECT 2181.3400 271.7000 2182.9400 272.1800 ;
        RECT 2181.3400 277.1400 2182.9400 277.6200 ;
        RECT 2174.1800 266.2600 2175.7800 266.7400 ;
        RECT 2174.1800 271.7000 2175.7800 272.1800 ;
        RECT 2174.1800 277.1400 2175.7800 277.6200 ;
        RECT 2181.3400 255.3800 2182.9400 255.8600 ;
        RECT 2181.3400 260.8200 2182.9400 261.3000 ;
        RECT 2174.1800 255.3800 2175.7800 255.8600 ;
        RECT 2174.1800 260.8200 2175.7800 261.3000 ;
        RECT 2181.3400 239.0600 2182.9400 239.5400 ;
        RECT 2181.3400 244.5000 2182.9400 244.9800 ;
        RECT 2181.3400 249.9400 2182.9400 250.4200 ;
        RECT 2174.1800 239.0600 2175.7800 239.5400 ;
        RECT 2174.1800 244.5000 2175.7800 244.9800 ;
        RECT 2174.1800 249.9400 2175.7800 250.4200 ;
        RECT 2271.3400 228.1800 2272.9400 228.6600 ;
        RECT 2271.3400 233.6200 2272.9400 234.1000 ;
        RECT 2271.3400 211.8600 2272.9400 212.3400 ;
        RECT 2271.3400 217.3000 2272.9400 217.7800 ;
        RECT 2271.3400 222.7400 2272.9400 223.2200 ;
        RECT 2226.3400 228.1800 2227.9400 228.6600 ;
        RECT 2226.3400 233.6200 2227.9400 234.1000 ;
        RECT 2226.3400 211.8600 2227.9400 212.3400 ;
        RECT 2226.3400 217.3000 2227.9400 217.7800 ;
        RECT 2226.3400 222.7400 2227.9400 223.2200 ;
        RECT 2271.3400 206.4200 2272.9400 206.9000 ;
        RECT 2271.3400 200.9800 2272.9400 201.4600 ;
        RECT 2271.3400 195.5400 2272.9400 196.0200 ;
        RECT 2226.3400 206.4200 2227.9400 206.9000 ;
        RECT 2226.3400 200.9800 2227.9400 201.4600 ;
        RECT 2226.3400 195.5400 2227.9400 196.0200 ;
        RECT 2181.3400 228.1800 2182.9400 228.6600 ;
        RECT 2181.3400 233.6200 2182.9400 234.1000 ;
        RECT 2174.1800 228.1800 2175.7800 228.6600 ;
        RECT 2174.1800 233.6200 2175.7800 234.1000 ;
        RECT 2181.3400 211.8600 2182.9400 212.3400 ;
        RECT 2181.3400 217.3000 2182.9400 217.7800 ;
        RECT 2181.3400 222.7400 2182.9400 223.2200 ;
        RECT 2174.1800 211.8600 2175.7800 212.3400 ;
        RECT 2174.1800 217.3000 2175.7800 217.7800 ;
        RECT 2174.1800 222.7400 2175.7800 223.2200 ;
        RECT 2181.3400 200.9800 2182.9400 201.4600 ;
        RECT 2181.3400 206.4200 2182.9400 206.9000 ;
        RECT 2174.1800 200.9800 2175.7800 201.4600 ;
        RECT 2174.1800 206.4200 2175.7800 206.9000 ;
        RECT 2174.1800 195.5400 2175.7800 196.0200 ;
        RECT 2181.3400 195.5400 2182.9400 196.0200 ;
        RECT 2171.2200 397.7300 2381.4400 399.3300 ;
        RECT 2171.2200 186.0300 2381.4400 187.6300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 183.2000 2175.7800 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 401.2400 2175.7800 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 183.2000 2378.4800 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 401.2400 2378.4800 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 186.0300 2172.8200 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 186.0300 2381.4400 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 397.7300 2172.8200 399.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 397.7300 2381.4400 399.3300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2174.2800 142.9400 2175.8800 173.2000 ;
        RECT 2376.7800 142.9400 2378.3800 173.2000 ;
      LAYER met3 ;
        RECT 2376.7800 163.4400 2378.3800 163.9200 ;
        RECT 2174.2800 163.4400 2175.8800 163.9200 ;
        RECT 2376.7800 152.5600 2378.3800 153.0400 ;
        RECT 2174.2800 152.5600 2175.8800 153.0400 ;
        RECT 2376.7800 158.0000 2378.3800 158.4800 ;
        RECT 2174.2800 158.0000 2175.8800 158.4800 ;
        RECT 2171.2200 168.8400 2381.4400 170.4400 ;
        RECT 2171.2200 144.5100 2381.4400 146.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.2800 142.9400 2175.8800 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.2800 171.6000 2175.8800 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.7800 142.9400 2378.3800 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.7800 171.6000 2378.3800 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 144.5100 2172.8200 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 144.5100 2381.4400 146.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 168.8400 2172.8200 170.4400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 168.8400 2381.4400 170.4400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 2252.7900 2362.9400 2466.0900 ;
        RECT 2316.3400 2252.7900 2317.9400 2466.0900 ;
        RECT 2271.3400 2252.7900 2272.9400 2466.0900 ;
        RECT 2226.3400 2252.7900 2227.9400 2466.0900 ;
        RECT 2181.3400 2252.7900 2182.9400 2466.0900 ;
        RECT 2376.8800 2249.9600 2378.4800 2469.6000 ;
        RECT 2174.1800 2249.9600 2175.7800 2469.6000 ;
      LAYER met3 ;
        RECT 2361.3400 2458.1400 2362.9400 2458.6200 ;
        RECT 2376.8800 2458.1400 2378.4800 2458.6200 ;
        RECT 2376.8800 2447.2600 2378.4800 2447.7400 ;
        RECT 2376.8800 2452.7000 2378.4800 2453.1800 ;
        RECT 2361.3400 2447.2600 2362.9400 2447.7400 ;
        RECT 2361.3400 2452.7000 2362.9400 2453.1800 ;
        RECT 2376.8800 2430.9400 2378.4800 2431.4200 ;
        RECT 2376.8800 2436.3800 2378.4800 2436.8600 ;
        RECT 2361.3400 2430.9400 2362.9400 2431.4200 ;
        RECT 2361.3400 2436.3800 2362.9400 2436.8600 ;
        RECT 2376.8800 2420.0600 2378.4800 2420.5400 ;
        RECT 2376.8800 2425.5000 2378.4800 2425.9800 ;
        RECT 2361.3400 2420.0600 2362.9400 2420.5400 ;
        RECT 2361.3400 2425.5000 2362.9400 2425.9800 ;
        RECT 2361.3400 2441.8200 2362.9400 2442.3000 ;
        RECT 2376.8800 2441.8200 2378.4800 2442.3000 ;
        RECT 2316.3400 2447.2600 2317.9400 2447.7400 ;
        RECT 2316.3400 2452.7000 2317.9400 2453.1800 ;
        RECT 2316.3400 2458.1400 2317.9400 2458.6200 ;
        RECT 2316.3400 2430.9400 2317.9400 2431.4200 ;
        RECT 2316.3400 2436.3800 2317.9400 2436.8600 ;
        RECT 2316.3400 2425.5000 2317.9400 2425.9800 ;
        RECT 2316.3400 2420.0600 2317.9400 2420.5400 ;
        RECT 2316.3400 2441.8200 2317.9400 2442.3000 ;
        RECT 2376.8800 2403.7400 2378.4800 2404.2200 ;
        RECT 2376.8800 2409.1800 2378.4800 2409.6600 ;
        RECT 2361.3400 2403.7400 2362.9400 2404.2200 ;
        RECT 2361.3400 2409.1800 2362.9400 2409.6600 ;
        RECT 2376.8800 2387.4200 2378.4800 2387.9000 ;
        RECT 2376.8800 2392.8600 2378.4800 2393.3400 ;
        RECT 2376.8800 2398.3000 2378.4800 2398.7800 ;
        RECT 2361.3400 2387.4200 2362.9400 2387.9000 ;
        RECT 2361.3400 2392.8600 2362.9400 2393.3400 ;
        RECT 2361.3400 2398.3000 2362.9400 2398.7800 ;
        RECT 2376.8800 2376.5400 2378.4800 2377.0200 ;
        RECT 2376.8800 2381.9800 2378.4800 2382.4600 ;
        RECT 2361.3400 2376.5400 2362.9400 2377.0200 ;
        RECT 2361.3400 2381.9800 2362.9400 2382.4600 ;
        RECT 2376.8800 2360.2200 2378.4800 2360.7000 ;
        RECT 2376.8800 2365.6600 2378.4800 2366.1400 ;
        RECT 2376.8800 2371.1000 2378.4800 2371.5800 ;
        RECT 2361.3400 2360.2200 2362.9400 2360.7000 ;
        RECT 2361.3400 2365.6600 2362.9400 2366.1400 ;
        RECT 2361.3400 2371.1000 2362.9400 2371.5800 ;
        RECT 2316.3400 2403.7400 2317.9400 2404.2200 ;
        RECT 2316.3400 2409.1800 2317.9400 2409.6600 ;
        RECT 2316.3400 2387.4200 2317.9400 2387.9000 ;
        RECT 2316.3400 2392.8600 2317.9400 2393.3400 ;
        RECT 2316.3400 2398.3000 2317.9400 2398.7800 ;
        RECT 2316.3400 2376.5400 2317.9400 2377.0200 ;
        RECT 2316.3400 2381.9800 2317.9400 2382.4600 ;
        RECT 2316.3400 2360.2200 2317.9400 2360.7000 ;
        RECT 2316.3400 2365.6600 2317.9400 2366.1400 ;
        RECT 2316.3400 2371.1000 2317.9400 2371.5800 ;
        RECT 2316.3400 2414.6200 2317.9400 2415.1000 ;
        RECT 2361.3400 2414.6200 2362.9400 2415.1000 ;
        RECT 2376.8800 2414.6200 2378.4800 2415.1000 ;
        RECT 2271.3400 2447.2600 2272.9400 2447.7400 ;
        RECT 2271.3400 2452.7000 2272.9400 2453.1800 ;
        RECT 2271.3400 2458.1400 2272.9400 2458.6200 ;
        RECT 2226.3400 2447.2600 2227.9400 2447.7400 ;
        RECT 2226.3400 2452.7000 2227.9400 2453.1800 ;
        RECT 2226.3400 2458.1400 2227.9400 2458.6200 ;
        RECT 2271.3400 2430.9400 2272.9400 2431.4200 ;
        RECT 2271.3400 2436.3800 2272.9400 2436.8600 ;
        RECT 2271.3400 2420.0600 2272.9400 2420.5400 ;
        RECT 2271.3400 2425.5000 2272.9400 2425.9800 ;
        RECT 2226.3400 2430.9400 2227.9400 2431.4200 ;
        RECT 2226.3400 2436.3800 2227.9400 2436.8600 ;
        RECT 2226.3400 2420.0600 2227.9400 2420.5400 ;
        RECT 2226.3400 2425.5000 2227.9400 2425.9800 ;
        RECT 2226.3400 2441.8200 2227.9400 2442.3000 ;
        RECT 2271.3400 2441.8200 2272.9400 2442.3000 ;
        RECT 2174.1800 2458.1400 2175.7800 2458.6200 ;
        RECT 2181.3400 2458.1400 2182.9400 2458.6200 ;
        RECT 2181.3400 2447.2600 2182.9400 2447.7400 ;
        RECT 2181.3400 2452.7000 2182.9400 2453.1800 ;
        RECT 2174.1800 2447.2600 2175.7800 2447.7400 ;
        RECT 2174.1800 2452.7000 2175.7800 2453.1800 ;
        RECT 2181.3400 2430.9400 2182.9400 2431.4200 ;
        RECT 2181.3400 2436.3800 2182.9400 2436.8600 ;
        RECT 2174.1800 2430.9400 2175.7800 2431.4200 ;
        RECT 2174.1800 2436.3800 2175.7800 2436.8600 ;
        RECT 2181.3400 2420.0600 2182.9400 2420.5400 ;
        RECT 2181.3400 2425.5000 2182.9400 2425.9800 ;
        RECT 2174.1800 2420.0600 2175.7800 2420.5400 ;
        RECT 2174.1800 2425.5000 2175.7800 2425.9800 ;
        RECT 2174.1800 2441.8200 2175.7800 2442.3000 ;
        RECT 2181.3400 2441.8200 2182.9400 2442.3000 ;
        RECT 2271.3400 2403.7400 2272.9400 2404.2200 ;
        RECT 2271.3400 2409.1800 2272.9400 2409.6600 ;
        RECT 2271.3400 2387.4200 2272.9400 2387.9000 ;
        RECT 2271.3400 2392.8600 2272.9400 2393.3400 ;
        RECT 2271.3400 2398.3000 2272.9400 2398.7800 ;
        RECT 2226.3400 2403.7400 2227.9400 2404.2200 ;
        RECT 2226.3400 2409.1800 2227.9400 2409.6600 ;
        RECT 2226.3400 2387.4200 2227.9400 2387.9000 ;
        RECT 2226.3400 2392.8600 2227.9400 2393.3400 ;
        RECT 2226.3400 2398.3000 2227.9400 2398.7800 ;
        RECT 2271.3400 2376.5400 2272.9400 2377.0200 ;
        RECT 2271.3400 2381.9800 2272.9400 2382.4600 ;
        RECT 2271.3400 2360.2200 2272.9400 2360.7000 ;
        RECT 2271.3400 2365.6600 2272.9400 2366.1400 ;
        RECT 2271.3400 2371.1000 2272.9400 2371.5800 ;
        RECT 2226.3400 2376.5400 2227.9400 2377.0200 ;
        RECT 2226.3400 2381.9800 2227.9400 2382.4600 ;
        RECT 2226.3400 2360.2200 2227.9400 2360.7000 ;
        RECT 2226.3400 2365.6600 2227.9400 2366.1400 ;
        RECT 2226.3400 2371.1000 2227.9400 2371.5800 ;
        RECT 2181.3400 2403.7400 2182.9400 2404.2200 ;
        RECT 2181.3400 2409.1800 2182.9400 2409.6600 ;
        RECT 2174.1800 2403.7400 2175.7800 2404.2200 ;
        RECT 2174.1800 2409.1800 2175.7800 2409.6600 ;
        RECT 2181.3400 2387.4200 2182.9400 2387.9000 ;
        RECT 2181.3400 2392.8600 2182.9400 2393.3400 ;
        RECT 2181.3400 2398.3000 2182.9400 2398.7800 ;
        RECT 2174.1800 2387.4200 2175.7800 2387.9000 ;
        RECT 2174.1800 2392.8600 2175.7800 2393.3400 ;
        RECT 2174.1800 2398.3000 2175.7800 2398.7800 ;
        RECT 2181.3400 2376.5400 2182.9400 2377.0200 ;
        RECT 2181.3400 2381.9800 2182.9400 2382.4600 ;
        RECT 2174.1800 2376.5400 2175.7800 2377.0200 ;
        RECT 2174.1800 2381.9800 2175.7800 2382.4600 ;
        RECT 2181.3400 2360.2200 2182.9400 2360.7000 ;
        RECT 2181.3400 2365.6600 2182.9400 2366.1400 ;
        RECT 2181.3400 2371.1000 2182.9400 2371.5800 ;
        RECT 2174.1800 2360.2200 2175.7800 2360.7000 ;
        RECT 2174.1800 2365.6600 2175.7800 2366.1400 ;
        RECT 2174.1800 2371.1000 2175.7800 2371.5800 ;
        RECT 2174.1800 2414.6200 2175.7800 2415.1000 ;
        RECT 2181.3400 2414.6200 2182.9400 2415.1000 ;
        RECT 2226.3400 2414.6200 2227.9400 2415.1000 ;
        RECT 2271.3400 2414.6200 2272.9400 2415.1000 ;
        RECT 2376.8800 2349.3400 2378.4800 2349.8200 ;
        RECT 2376.8800 2354.7800 2378.4800 2355.2600 ;
        RECT 2361.3400 2349.3400 2362.9400 2349.8200 ;
        RECT 2361.3400 2354.7800 2362.9400 2355.2600 ;
        RECT 2376.8800 2333.0200 2378.4800 2333.5000 ;
        RECT 2376.8800 2338.4600 2378.4800 2338.9400 ;
        RECT 2376.8800 2343.9000 2378.4800 2344.3800 ;
        RECT 2361.3400 2333.0200 2362.9400 2333.5000 ;
        RECT 2361.3400 2338.4600 2362.9400 2338.9400 ;
        RECT 2361.3400 2343.9000 2362.9400 2344.3800 ;
        RECT 2376.8800 2322.1400 2378.4800 2322.6200 ;
        RECT 2376.8800 2327.5800 2378.4800 2328.0600 ;
        RECT 2361.3400 2322.1400 2362.9400 2322.6200 ;
        RECT 2361.3400 2327.5800 2362.9400 2328.0600 ;
        RECT 2376.8800 2305.8200 2378.4800 2306.3000 ;
        RECT 2376.8800 2311.2600 2378.4800 2311.7400 ;
        RECT 2376.8800 2316.7000 2378.4800 2317.1800 ;
        RECT 2361.3400 2305.8200 2362.9400 2306.3000 ;
        RECT 2361.3400 2311.2600 2362.9400 2311.7400 ;
        RECT 2361.3400 2316.7000 2362.9400 2317.1800 ;
        RECT 2316.3400 2349.3400 2317.9400 2349.8200 ;
        RECT 2316.3400 2354.7800 2317.9400 2355.2600 ;
        RECT 2316.3400 2333.0200 2317.9400 2333.5000 ;
        RECT 2316.3400 2338.4600 2317.9400 2338.9400 ;
        RECT 2316.3400 2343.9000 2317.9400 2344.3800 ;
        RECT 2316.3400 2322.1400 2317.9400 2322.6200 ;
        RECT 2316.3400 2327.5800 2317.9400 2328.0600 ;
        RECT 2316.3400 2305.8200 2317.9400 2306.3000 ;
        RECT 2316.3400 2311.2600 2317.9400 2311.7400 ;
        RECT 2316.3400 2316.7000 2317.9400 2317.1800 ;
        RECT 2376.8800 2294.9400 2378.4800 2295.4200 ;
        RECT 2376.8800 2300.3800 2378.4800 2300.8600 ;
        RECT 2361.3400 2294.9400 2362.9400 2295.4200 ;
        RECT 2361.3400 2300.3800 2362.9400 2300.8600 ;
        RECT 2376.8800 2278.6200 2378.4800 2279.1000 ;
        RECT 2376.8800 2284.0600 2378.4800 2284.5400 ;
        RECT 2376.8800 2289.5000 2378.4800 2289.9800 ;
        RECT 2361.3400 2278.6200 2362.9400 2279.1000 ;
        RECT 2361.3400 2284.0600 2362.9400 2284.5400 ;
        RECT 2361.3400 2289.5000 2362.9400 2289.9800 ;
        RECT 2376.8800 2267.7400 2378.4800 2268.2200 ;
        RECT 2376.8800 2273.1800 2378.4800 2273.6600 ;
        RECT 2361.3400 2267.7400 2362.9400 2268.2200 ;
        RECT 2361.3400 2273.1800 2362.9400 2273.6600 ;
        RECT 2361.3400 2262.3000 2362.9400 2262.7800 ;
        RECT 2376.8800 2262.3000 2378.4800 2262.7800 ;
        RECT 2316.3400 2294.9400 2317.9400 2295.4200 ;
        RECT 2316.3400 2300.3800 2317.9400 2300.8600 ;
        RECT 2316.3400 2278.6200 2317.9400 2279.1000 ;
        RECT 2316.3400 2284.0600 2317.9400 2284.5400 ;
        RECT 2316.3400 2289.5000 2317.9400 2289.9800 ;
        RECT 2316.3400 2267.7400 2317.9400 2268.2200 ;
        RECT 2316.3400 2273.1800 2317.9400 2273.6600 ;
        RECT 2316.3400 2262.3000 2317.9400 2262.7800 ;
        RECT 2271.3400 2349.3400 2272.9400 2349.8200 ;
        RECT 2271.3400 2354.7800 2272.9400 2355.2600 ;
        RECT 2271.3400 2333.0200 2272.9400 2333.5000 ;
        RECT 2271.3400 2338.4600 2272.9400 2338.9400 ;
        RECT 2271.3400 2343.9000 2272.9400 2344.3800 ;
        RECT 2226.3400 2349.3400 2227.9400 2349.8200 ;
        RECT 2226.3400 2354.7800 2227.9400 2355.2600 ;
        RECT 2226.3400 2333.0200 2227.9400 2333.5000 ;
        RECT 2226.3400 2338.4600 2227.9400 2338.9400 ;
        RECT 2226.3400 2343.9000 2227.9400 2344.3800 ;
        RECT 2271.3400 2322.1400 2272.9400 2322.6200 ;
        RECT 2271.3400 2327.5800 2272.9400 2328.0600 ;
        RECT 2271.3400 2305.8200 2272.9400 2306.3000 ;
        RECT 2271.3400 2311.2600 2272.9400 2311.7400 ;
        RECT 2271.3400 2316.7000 2272.9400 2317.1800 ;
        RECT 2226.3400 2322.1400 2227.9400 2322.6200 ;
        RECT 2226.3400 2327.5800 2227.9400 2328.0600 ;
        RECT 2226.3400 2305.8200 2227.9400 2306.3000 ;
        RECT 2226.3400 2311.2600 2227.9400 2311.7400 ;
        RECT 2226.3400 2316.7000 2227.9400 2317.1800 ;
        RECT 2181.3400 2349.3400 2182.9400 2349.8200 ;
        RECT 2181.3400 2354.7800 2182.9400 2355.2600 ;
        RECT 2174.1800 2349.3400 2175.7800 2349.8200 ;
        RECT 2174.1800 2354.7800 2175.7800 2355.2600 ;
        RECT 2181.3400 2333.0200 2182.9400 2333.5000 ;
        RECT 2181.3400 2338.4600 2182.9400 2338.9400 ;
        RECT 2181.3400 2343.9000 2182.9400 2344.3800 ;
        RECT 2174.1800 2333.0200 2175.7800 2333.5000 ;
        RECT 2174.1800 2338.4600 2175.7800 2338.9400 ;
        RECT 2174.1800 2343.9000 2175.7800 2344.3800 ;
        RECT 2181.3400 2322.1400 2182.9400 2322.6200 ;
        RECT 2181.3400 2327.5800 2182.9400 2328.0600 ;
        RECT 2174.1800 2322.1400 2175.7800 2322.6200 ;
        RECT 2174.1800 2327.5800 2175.7800 2328.0600 ;
        RECT 2181.3400 2305.8200 2182.9400 2306.3000 ;
        RECT 2181.3400 2311.2600 2182.9400 2311.7400 ;
        RECT 2181.3400 2316.7000 2182.9400 2317.1800 ;
        RECT 2174.1800 2305.8200 2175.7800 2306.3000 ;
        RECT 2174.1800 2311.2600 2175.7800 2311.7400 ;
        RECT 2174.1800 2316.7000 2175.7800 2317.1800 ;
        RECT 2271.3400 2294.9400 2272.9400 2295.4200 ;
        RECT 2271.3400 2300.3800 2272.9400 2300.8600 ;
        RECT 2271.3400 2278.6200 2272.9400 2279.1000 ;
        RECT 2271.3400 2284.0600 2272.9400 2284.5400 ;
        RECT 2271.3400 2289.5000 2272.9400 2289.9800 ;
        RECT 2226.3400 2294.9400 2227.9400 2295.4200 ;
        RECT 2226.3400 2300.3800 2227.9400 2300.8600 ;
        RECT 2226.3400 2278.6200 2227.9400 2279.1000 ;
        RECT 2226.3400 2284.0600 2227.9400 2284.5400 ;
        RECT 2226.3400 2289.5000 2227.9400 2289.9800 ;
        RECT 2271.3400 2273.1800 2272.9400 2273.6600 ;
        RECT 2271.3400 2267.7400 2272.9400 2268.2200 ;
        RECT 2271.3400 2262.3000 2272.9400 2262.7800 ;
        RECT 2226.3400 2273.1800 2227.9400 2273.6600 ;
        RECT 2226.3400 2267.7400 2227.9400 2268.2200 ;
        RECT 2226.3400 2262.3000 2227.9400 2262.7800 ;
        RECT 2181.3400 2294.9400 2182.9400 2295.4200 ;
        RECT 2181.3400 2300.3800 2182.9400 2300.8600 ;
        RECT 2174.1800 2294.9400 2175.7800 2295.4200 ;
        RECT 2174.1800 2300.3800 2175.7800 2300.8600 ;
        RECT 2181.3400 2278.6200 2182.9400 2279.1000 ;
        RECT 2181.3400 2284.0600 2182.9400 2284.5400 ;
        RECT 2181.3400 2289.5000 2182.9400 2289.9800 ;
        RECT 2174.1800 2278.6200 2175.7800 2279.1000 ;
        RECT 2174.1800 2284.0600 2175.7800 2284.5400 ;
        RECT 2174.1800 2289.5000 2175.7800 2289.9800 ;
        RECT 2181.3400 2267.7400 2182.9400 2268.2200 ;
        RECT 2181.3400 2273.1800 2182.9400 2273.6600 ;
        RECT 2174.1800 2267.7400 2175.7800 2268.2200 ;
        RECT 2174.1800 2273.1800 2175.7800 2273.6600 ;
        RECT 2174.1800 2262.3000 2175.7800 2262.7800 ;
        RECT 2181.3400 2262.3000 2182.9400 2262.7800 ;
        RECT 2171.2200 2464.4900 2381.4400 2466.0900 ;
        RECT 2171.2200 2252.7900 2381.4400 2254.3900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 2249.9600 2175.7800 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 2468.0000 2175.7800 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 2249.9600 2378.4800 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 2468.0000 2378.4800 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2252.7900 2172.8200 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2252.7900 2381.4400 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2464.4900 2172.8200 2466.0900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2464.4900 2381.4400 2466.0900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 2023.1500 2362.9400 2236.4500 ;
        RECT 2316.3400 2023.1500 2317.9400 2236.4500 ;
        RECT 2271.3400 2023.1500 2272.9400 2236.4500 ;
        RECT 2226.3400 2023.1500 2227.9400 2236.4500 ;
        RECT 2181.3400 2023.1500 2182.9400 2236.4500 ;
        RECT 2376.8800 2020.3200 2378.4800 2239.9600 ;
        RECT 2174.1800 2020.3200 2175.7800 2239.9600 ;
      LAYER met3 ;
        RECT 2361.3400 2228.5000 2362.9400 2228.9800 ;
        RECT 2376.8800 2228.5000 2378.4800 2228.9800 ;
        RECT 2376.8800 2217.6200 2378.4800 2218.1000 ;
        RECT 2376.8800 2223.0600 2378.4800 2223.5400 ;
        RECT 2361.3400 2217.6200 2362.9400 2218.1000 ;
        RECT 2361.3400 2223.0600 2362.9400 2223.5400 ;
        RECT 2376.8800 2201.3000 2378.4800 2201.7800 ;
        RECT 2376.8800 2206.7400 2378.4800 2207.2200 ;
        RECT 2361.3400 2201.3000 2362.9400 2201.7800 ;
        RECT 2361.3400 2206.7400 2362.9400 2207.2200 ;
        RECT 2376.8800 2190.4200 2378.4800 2190.9000 ;
        RECT 2376.8800 2195.8600 2378.4800 2196.3400 ;
        RECT 2361.3400 2190.4200 2362.9400 2190.9000 ;
        RECT 2361.3400 2195.8600 2362.9400 2196.3400 ;
        RECT 2361.3400 2212.1800 2362.9400 2212.6600 ;
        RECT 2376.8800 2212.1800 2378.4800 2212.6600 ;
        RECT 2316.3400 2217.6200 2317.9400 2218.1000 ;
        RECT 2316.3400 2223.0600 2317.9400 2223.5400 ;
        RECT 2316.3400 2228.5000 2317.9400 2228.9800 ;
        RECT 2316.3400 2201.3000 2317.9400 2201.7800 ;
        RECT 2316.3400 2206.7400 2317.9400 2207.2200 ;
        RECT 2316.3400 2195.8600 2317.9400 2196.3400 ;
        RECT 2316.3400 2190.4200 2317.9400 2190.9000 ;
        RECT 2316.3400 2212.1800 2317.9400 2212.6600 ;
        RECT 2376.8800 2174.1000 2378.4800 2174.5800 ;
        RECT 2376.8800 2179.5400 2378.4800 2180.0200 ;
        RECT 2361.3400 2174.1000 2362.9400 2174.5800 ;
        RECT 2361.3400 2179.5400 2362.9400 2180.0200 ;
        RECT 2376.8800 2157.7800 2378.4800 2158.2600 ;
        RECT 2376.8800 2163.2200 2378.4800 2163.7000 ;
        RECT 2376.8800 2168.6600 2378.4800 2169.1400 ;
        RECT 2361.3400 2157.7800 2362.9400 2158.2600 ;
        RECT 2361.3400 2163.2200 2362.9400 2163.7000 ;
        RECT 2361.3400 2168.6600 2362.9400 2169.1400 ;
        RECT 2376.8800 2146.9000 2378.4800 2147.3800 ;
        RECT 2376.8800 2152.3400 2378.4800 2152.8200 ;
        RECT 2361.3400 2146.9000 2362.9400 2147.3800 ;
        RECT 2361.3400 2152.3400 2362.9400 2152.8200 ;
        RECT 2376.8800 2130.5800 2378.4800 2131.0600 ;
        RECT 2376.8800 2136.0200 2378.4800 2136.5000 ;
        RECT 2376.8800 2141.4600 2378.4800 2141.9400 ;
        RECT 2361.3400 2130.5800 2362.9400 2131.0600 ;
        RECT 2361.3400 2136.0200 2362.9400 2136.5000 ;
        RECT 2361.3400 2141.4600 2362.9400 2141.9400 ;
        RECT 2316.3400 2174.1000 2317.9400 2174.5800 ;
        RECT 2316.3400 2179.5400 2317.9400 2180.0200 ;
        RECT 2316.3400 2157.7800 2317.9400 2158.2600 ;
        RECT 2316.3400 2163.2200 2317.9400 2163.7000 ;
        RECT 2316.3400 2168.6600 2317.9400 2169.1400 ;
        RECT 2316.3400 2146.9000 2317.9400 2147.3800 ;
        RECT 2316.3400 2152.3400 2317.9400 2152.8200 ;
        RECT 2316.3400 2130.5800 2317.9400 2131.0600 ;
        RECT 2316.3400 2136.0200 2317.9400 2136.5000 ;
        RECT 2316.3400 2141.4600 2317.9400 2141.9400 ;
        RECT 2316.3400 2184.9800 2317.9400 2185.4600 ;
        RECT 2361.3400 2184.9800 2362.9400 2185.4600 ;
        RECT 2376.8800 2184.9800 2378.4800 2185.4600 ;
        RECT 2271.3400 2217.6200 2272.9400 2218.1000 ;
        RECT 2271.3400 2223.0600 2272.9400 2223.5400 ;
        RECT 2271.3400 2228.5000 2272.9400 2228.9800 ;
        RECT 2226.3400 2217.6200 2227.9400 2218.1000 ;
        RECT 2226.3400 2223.0600 2227.9400 2223.5400 ;
        RECT 2226.3400 2228.5000 2227.9400 2228.9800 ;
        RECT 2271.3400 2201.3000 2272.9400 2201.7800 ;
        RECT 2271.3400 2206.7400 2272.9400 2207.2200 ;
        RECT 2271.3400 2190.4200 2272.9400 2190.9000 ;
        RECT 2271.3400 2195.8600 2272.9400 2196.3400 ;
        RECT 2226.3400 2201.3000 2227.9400 2201.7800 ;
        RECT 2226.3400 2206.7400 2227.9400 2207.2200 ;
        RECT 2226.3400 2190.4200 2227.9400 2190.9000 ;
        RECT 2226.3400 2195.8600 2227.9400 2196.3400 ;
        RECT 2226.3400 2212.1800 2227.9400 2212.6600 ;
        RECT 2271.3400 2212.1800 2272.9400 2212.6600 ;
        RECT 2174.1800 2228.5000 2175.7800 2228.9800 ;
        RECT 2181.3400 2228.5000 2182.9400 2228.9800 ;
        RECT 2181.3400 2217.6200 2182.9400 2218.1000 ;
        RECT 2181.3400 2223.0600 2182.9400 2223.5400 ;
        RECT 2174.1800 2217.6200 2175.7800 2218.1000 ;
        RECT 2174.1800 2223.0600 2175.7800 2223.5400 ;
        RECT 2181.3400 2201.3000 2182.9400 2201.7800 ;
        RECT 2181.3400 2206.7400 2182.9400 2207.2200 ;
        RECT 2174.1800 2201.3000 2175.7800 2201.7800 ;
        RECT 2174.1800 2206.7400 2175.7800 2207.2200 ;
        RECT 2181.3400 2190.4200 2182.9400 2190.9000 ;
        RECT 2181.3400 2195.8600 2182.9400 2196.3400 ;
        RECT 2174.1800 2190.4200 2175.7800 2190.9000 ;
        RECT 2174.1800 2195.8600 2175.7800 2196.3400 ;
        RECT 2174.1800 2212.1800 2175.7800 2212.6600 ;
        RECT 2181.3400 2212.1800 2182.9400 2212.6600 ;
        RECT 2271.3400 2174.1000 2272.9400 2174.5800 ;
        RECT 2271.3400 2179.5400 2272.9400 2180.0200 ;
        RECT 2271.3400 2157.7800 2272.9400 2158.2600 ;
        RECT 2271.3400 2163.2200 2272.9400 2163.7000 ;
        RECT 2271.3400 2168.6600 2272.9400 2169.1400 ;
        RECT 2226.3400 2174.1000 2227.9400 2174.5800 ;
        RECT 2226.3400 2179.5400 2227.9400 2180.0200 ;
        RECT 2226.3400 2157.7800 2227.9400 2158.2600 ;
        RECT 2226.3400 2163.2200 2227.9400 2163.7000 ;
        RECT 2226.3400 2168.6600 2227.9400 2169.1400 ;
        RECT 2271.3400 2146.9000 2272.9400 2147.3800 ;
        RECT 2271.3400 2152.3400 2272.9400 2152.8200 ;
        RECT 2271.3400 2130.5800 2272.9400 2131.0600 ;
        RECT 2271.3400 2136.0200 2272.9400 2136.5000 ;
        RECT 2271.3400 2141.4600 2272.9400 2141.9400 ;
        RECT 2226.3400 2146.9000 2227.9400 2147.3800 ;
        RECT 2226.3400 2152.3400 2227.9400 2152.8200 ;
        RECT 2226.3400 2130.5800 2227.9400 2131.0600 ;
        RECT 2226.3400 2136.0200 2227.9400 2136.5000 ;
        RECT 2226.3400 2141.4600 2227.9400 2141.9400 ;
        RECT 2181.3400 2174.1000 2182.9400 2174.5800 ;
        RECT 2181.3400 2179.5400 2182.9400 2180.0200 ;
        RECT 2174.1800 2174.1000 2175.7800 2174.5800 ;
        RECT 2174.1800 2179.5400 2175.7800 2180.0200 ;
        RECT 2181.3400 2157.7800 2182.9400 2158.2600 ;
        RECT 2181.3400 2163.2200 2182.9400 2163.7000 ;
        RECT 2181.3400 2168.6600 2182.9400 2169.1400 ;
        RECT 2174.1800 2157.7800 2175.7800 2158.2600 ;
        RECT 2174.1800 2163.2200 2175.7800 2163.7000 ;
        RECT 2174.1800 2168.6600 2175.7800 2169.1400 ;
        RECT 2181.3400 2146.9000 2182.9400 2147.3800 ;
        RECT 2181.3400 2152.3400 2182.9400 2152.8200 ;
        RECT 2174.1800 2146.9000 2175.7800 2147.3800 ;
        RECT 2174.1800 2152.3400 2175.7800 2152.8200 ;
        RECT 2181.3400 2130.5800 2182.9400 2131.0600 ;
        RECT 2181.3400 2136.0200 2182.9400 2136.5000 ;
        RECT 2181.3400 2141.4600 2182.9400 2141.9400 ;
        RECT 2174.1800 2130.5800 2175.7800 2131.0600 ;
        RECT 2174.1800 2136.0200 2175.7800 2136.5000 ;
        RECT 2174.1800 2141.4600 2175.7800 2141.9400 ;
        RECT 2174.1800 2184.9800 2175.7800 2185.4600 ;
        RECT 2181.3400 2184.9800 2182.9400 2185.4600 ;
        RECT 2226.3400 2184.9800 2227.9400 2185.4600 ;
        RECT 2271.3400 2184.9800 2272.9400 2185.4600 ;
        RECT 2376.8800 2119.7000 2378.4800 2120.1800 ;
        RECT 2376.8800 2125.1400 2378.4800 2125.6200 ;
        RECT 2361.3400 2119.7000 2362.9400 2120.1800 ;
        RECT 2361.3400 2125.1400 2362.9400 2125.6200 ;
        RECT 2376.8800 2103.3800 2378.4800 2103.8600 ;
        RECT 2376.8800 2108.8200 2378.4800 2109.3000 ;
        RECT 2376.8800 2114.2600 2378.4800 2114.7400 ;
        RECT 2361.3400 2103.3800 2362.9400 2103.8600 ;
        RECT 2361.3400 2108.8200 2362.9400 2109.3000 ;
        RECT 2361.3400 2114.2600 2362.9400 2114.7400 ;
        RECT 2376.8800 2092.5000 2378.4800 2092.9800 ;
        RECT 2376.8800 2097.9400 2378.4800 2098.4200 ;
        RECT 2361.3400 2092.5000 2362.9400 2092.9800 ;
        RECT 2361.3400 2097.9400 2362.9400 2098.4200 ;
        RECT 2376.8800 2076.1800 2378.4800 2076.6600 ;
        RECT 2376.8800 2081.6200 2378.4800 2082.1000 ;
        RECT 2376.8800 2087.0600 2378.4800 2087.5400 ;
        RECT 2361.3400 2076.1800 2362.9400 2076.6600 ;
        RECT 2361.3400 2081.6200 2362.9400 2082.1000 ;
        RECT 2361.3400 2087.0600 2362.9400 2087.5400 ;
        RECT 2316.3400 2119.7000 2317.9400 2120.1800 ;
        RECT 2316.3400 2125.1400 2317.9400 2125.6200 ;
        RECT 2316.3400 2103.3800 2317.9400 2103.8600 ;
        RECT 2316.3400 2108.8200 2317.9400 2109.3000 ;
        RECT 2316.3400 2114.2600 2317.9400 2114.7400 ;
        RECT 2316.3400 2092.5000 2317.9400 2092.9800 ;
        RECT 2316.3400 2097.9400 2317.9400 2098.4200 ;
        RECT 2316.3400 2076.1800 2317.9400 2076.6600 ;
        RECT 2316.3400 2081.6200 2317.9400 2082.1000 ;
        RECT 2316.3400 2087.0600 2317.9400 2087.5400 ;
        RECT 2376.8800 2065.3000 2378.4800 2065.7800 ;
        RECT 2376.8800 2070.7400 2378.4800 2071.2200 ;
        RECT 2361.3400 2065.3000 2362.9400 2065.7800 ;
        RECT 2361.3400 2070.7400 2362.9400 2071.2200 ;
        RECT 2376.8800 2048.9800 2378.4800 2049.4600 ;
        RECT 2376.8800 2054.4200 2378.4800 2054.9000 ;
        RECT 2376.8800 2059.8600 2378.4800 2060.3400 ;
        RECT 2361.3400 2048.9800 2362.9400 2049.4600 ;
        RECT 2361.3400 2054.4200 2362.9400 2054.9000 ;
        RECT 2361.3400 2059.8600 2362.9400 2060.3400 ;
        RECT 2376.8800 2038.1000 2378.4800 2038.5800 ;
        RECT 2376.8800 2043.5400 2378.4800 2044.0200 ;
        RECT 2361.3400 2038.1000 2362.9400 2038.5800 ;
        RECT 2361.3400 2043.5400 2362.9400 2044.0200 ;
        RECT 2361.3400 2032.6600 2362.9400 2033.1400 ;
        RECT 2376.8800 2032.6600 2378.4800 2033.1400 ;
        RECT 2316.3400 2065.3000 2317.9400 2065.7800 ;
        RECT 2316.3400 2070.7400 2317.9400 2071.2200 ;
        RECT 2316.3400 2048.9800 2317.9400 2049.4600 ;
        RECT 2316.3400 2054.4200 2317.9400 2054.9000 ;
        RECT 2316.3400 2059.8600 2317.9400 2060.3400 ;
        RECT 2316.3400 2038.1000 2317.9400 2038.5800 ;
        RECT 2316.3400 2043.5400 2317.9400 2044.0200 ;
        RECT 2316.3400 2032.6600 2317.9400 2033.1400 ;
        RECT 2271.3400 2119.7000 2272.9400 2120.1800 ;
        RECT 2271.3400 2125.1400 2272.9400 2125.6200 ;
        RECT 2271.3400 2103.3800 2272.9400 2103.8600 ;
        RECT 2271.3400 2108.8200 2272.9400 2109.3000 ;
        RECT 2271.3400 2114.2600 2272.9400 2114.7400 ;
        RECT 2226.3400 2119.7000 2227.9400 2120.1800 ;
        RECT 2226.3400 2125.1400 2227.9400 2125.6200 ;
        RECT 2226.3400 2103.3800 2227.9400 2103.8600 ;
        RECT 2226.3400 2108.8200 2227.9400 2109.3000 ;
        RECT 2226.3400 2114.2600 2227.9400 2114.7400 ;
        RECT 2271.3400 2092.5000 2272.9400 2092.9800 ;
        RECT 2271.3400 2097.9400 2272.9400 2098.4200 ;
        RECT 2271.3400 2076.1800 2272.9400 2076.6600 ;
        RECT 2271.3400 2081.6200 2272.9400 2082.1000 ;
        RECT 2271.3400 2087.0600 2272.9400 2087.5400 ;
        RECT 2226.3400 2092.5000 2227.9400 2092.9800 ;
        RECT 2226.3400 2097.9400 2227.9400 2098.4200 ;
        RECT 2226.3400 2076.1800 2227.9400 2076.6600 ;
        RECT 2226.3400 2081.6200 2227.9400 2082.1000 ;
        RECT 2226.3400 2087.0600 2227.9400 2087.5400 ;
        RECT 2181.3400 2119.7000 2182.9400 2120.1800 ;
        RECT 2181.3400 2125.1400 2182.9400 2125.6200 ;
        RECT 2174.1800 2119.7000 2175.7800 2120.1800 ;
        RECT 2174.1800 2125.1400 2175.7800 2125.6200 ;
        RECT 2181.3400 2103.3800 2182.9400 2103.8600 ;
        RECT 2181.3400 2108.8200 2182.9400 2109.3000 ;
        RECT 2181.3400 2114.2600 2182.9400 2114.7400 ;
        RECT 2174.1800 2103.3800 2175.7800 2103.8600 ;
        RECT 2174.1800 2108.8200 2175.7800 2109.3000 ;
        RECT 2174.1800 2114.2600 2175.7800 2114.7400 ;
        RECT 2181.3400 2092.5000 2182.9400 2092.9800 ;
        RECT 2181.3400 2097.9400 2182.9400 2098.4200 ;
        RECT 2174.1800 2092.5000 2175.7800 2092.9800 ;
        RECT 2174.1800 2097.9400 2175.7800 2098.4200 ;
        RECT 2181.3400 2076.1800 2182.9400 2076.6600 ;
        RECT 2181.3400 2081.6200 2182.9400 2082.1000 ;
        RECT 2181.3400 2087.0600 2182.9400 2087.5400 ;
        RECT 2174.1800 2076.1800 2175.7800 2076.6600 ;
        RECT 2174.1800 2081.6200 2175.7800 2082.1000 ;
        RECT 2174.1800 2087.0600 2175.7800 2087.5400 ;
        RECT 2271.3400 2065.3000 2272.9400 2065.7800 ;
        RECT 2271.3400 2070.7400 2272.9400 2071.2200 ;
        RECT 2271.3400 2048.9800 2272.9400 2049.4600 ;
        RECT 2271.3400 2054.4200 2272.9400 2054.9000 ;
        RECT 2271.3400 2059.8600 2272.9400 2060.3400 ;
        RECT 2226.3400 2065.3000 2227.9400 2065.7800 ;
        RECT 2226.3400 2070.7400 2227.9400 2071.2200 ;
        RECT 2226.3400 2048.9800 2227.9400 2049.4600 ;
        RECT 2226.3400 2054.4200 2227.9400 2054.9000 ;
        RECT 2226.3400 2059.8600 2227.9400 2060.3400 ;
        RECT 2271.3400 2043.5400 2272.9400 2044.0200 ;
        RECT 2271.3400 2038.1000 2272.9400 2038.5800 ;
        RECT 2271.3400 2032.6600 2272.9400 2033.1400 ;
        RECT 2226.3400 2043.5400 2227.9400 2044.0200 ;
        RECT 2226.3400 2038.1000 2227.9400 2038.5800 ;
        RECT 2226.3400 2032.6600 2227.9400 2033.1400 ;
        RECT 2181.3400 2065.3000 2182.9400 2065.7800 ;
        RECT 2181.3400 2070.7400 2182.9400 2071.2200 ;
        RECT 2174.1800 2065.3000 2175.7800 2065.7800 ;
        RECT 2174.1800 2070.7400 2175.7800 2071.2200 ;
        RECT 2181.3400 2048.9800 2182.9400 2049.4600 ;
        RECT 2181.3400 2054.4200 2182.9400 2054.9000 ;
        RECT 2181.3400 2059.8600 2182.9400 2060.3400 ;
        RECT 2174.1800 2048.9800 2175.7800 2049.4600 ;
        RECT 2174.1800 2054.4200 2175.7800 2054.9000 ;
        RECT 2174.1800 2059.8600 2175.7800 2060.3400 ;
        RECT 2181.3400 2038.1000 2182.9400 2038.5800 ;
        RECT 2181.3400 2043.5400 2182.9400 2044.0200 ;
        RECT 2174.1800 2038.1000 2175.7800 2038.5800 ;
        RECT 2174.1800 2043.5400 2175.7800 2044.0200 ;
        RECT 2174.1800 2032.6600 2175.7800 2033.1400 ;
        RECT 2181.3400 2032.6600 2182.9400 2033.1400 ;
        RECT 2171.2200 2234.8500 2381.4400 2236.4500 ;
        RECT 2171.2200 2023.1500 2381.4400 2024.7500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 2020.3200 2175.7800 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 2238.3600 2175.7800 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 2020.3200 2378.4800 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 2238.3600 2378.4800 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2023.1500 2172.8200 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2023.1500 2381.4400 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2234.8500 2172.8200 2236.4500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2234.8500 2381.4400 2236.4500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 1793.5100 2362.9400 2006.8100 ;
        RECT 2316.3400 1793.5100 2317.9400 2006.8100 ;
        RECT 2271.3400 1793.5100 2272.9400 2006.8100 ;
        RECT 2226.3400 1793.5100 2227.9400 2006.8100 ;
        RECT 2181.3400 1793.5100 2182.9400 2006.8100 ;
        RECT 2376.8800 1790.6800 2378.4800 2010.3200 ;
        RECT 2174.1800 1790.6800 2175.7800 2010.3200 ;
      LAYER met3 ;
        RECT 2361.3400 1998.8600 2362.9400 1999.3400 ;
        RECT 2376.8800 1998.8600 2378.4800 1999.3400 ;
        RECT 2376.8800 1987.9800 2378.4800 1988.4600 ;
        RECT 2376.8800 1993.4200 2378.4800 1993.9000 ;
        RECT 2361.3400 1987.9800 2362.9400 1988.4600 ;
        RECT 2361.3400 1993.4200 2362.9400 1993.9000 ;
        RECT 2376.8800 1971.6600 2378.4800 1972.1400 ;
        RECT 2376.8800 1977.1000 2378.4800 1977.5800 ;
        RECT 2361.3400 1971.6600 2362.9400 1972.1400 ;
        RECT 2361.3400 1977.1000 2362.9400 1977.5800 ;
        RECT 2376.8800 1960.7800 2378.4800 1961.2600 ;
        RECT 2376.8800 1966.2200 2378.4800 1966.7000 ;
        RECT 2361.3400 1960.7800 2362.9400 1961.2600 ;
        RECT 2361.3400 1966.2200 2362.9400 1966.7000 ;
        RECT 2361.3400 1982.5400 2362.9400 1983.0200 ;
        RECT 2376.8800 1982.5400 2378.4800 1983.0200 ;
        RECT 2316.3400 1987.9800 2317.9400 1988.4600 ;
        RECT 2316.3400 1993.4200 2317.9400 1993.9000 ;
        RECT 2316.3400 1998.8600 2317.9400 1999.3400 ;
        RECT 2316.3400 1971.6600 2317.9400 1972.1400 ;
        RECT 2316.3400 1977.1000 2317.9400 1977.5800 ;
        RECT 2316.3400 1966.2200 2317.9400 1966.7000 ;
        RECT 2316.3400 1960.7800 2317.9400 1961.2600 ;
        RECT 2316.3400 1982.5400 2317.9400 1983.0200 ;
        RECT 2376.8800 1944.4600 2378.4800 1944.9400 ;
        RECT 2376.8800 1949.9000 2378.4800 1950.3800 ;
        RECT 2361.3400 1944.4600 2362.9400 1944.9400 ;
        RECT 2361.3400 1949.9000 2362.9400 1950.3800 ;
        RECT 2376.8800 1928.1400 2378.4800 1928.6200 ;
        RECT 2376.8800 1933.5800 2378.4800 1934.0600 ;
        RECT 2376.8800 1939.0200 2378.4800 1939.5000 ;
        RECT 2361.3400 1928.1400 2362.9400 1928.6200 ;
        RECT 2361.3400 1933.5800 2362.9400 1934.0600 ;
        RECT 2361.3400 1939.0200 2362.9400 1939.5000 ;
        RECT 2376.8800 1917.2600 2378.4800 1917.7400 ;
        RECT 2376.8800 1922.7000 2378.4800 1923.1800 ;
        RECT 2361.3400 1917.2600 2362.9400 1917.7400 ;
        RECT 2361.3400 1922.7000 2362.9400 1923.1800 ;
        RECT 2376.8800 1900.9400 2378.4800 1901.4200 ;
        RECT 2376.8800 1906.3800 2378.4800 1906.8600 ;
        RECT 2376.8800 1911.8200 2378.4800 1912.3000 ;
        RECT 2361.3400 1900.9400 2362.9400 1901.4200 ;
        RECT 2361.3400 1906.3800 2362.9400 1906.8600 ;
        RECT 2361.3400 1911.8200 2362.9400 1912.3000 ;
        RECT 2316.3400 1944.4600 2317.9400 1944.9400 ;
        RECT 2316.3400 1949.9000 2317.9400 1950.3800 ;
        RECT 2316.3400 1928.1400 2317.9400 1928.6200 ;
        RECT 2316.3400 1933.5800 2317.9400 1934.0600 ;
        RECT 2316.3400 1939.0200 2317.9400 1939.5000 ;
        RECT 2316.3400 1917.2600 2317.9400 1917.7400 ;
        RECT 2316.3400 1922.7000 2317.9400 1923.1800 ;
        RECT 2316.3400 1900.9400 2317.9400 1901.4200 ;
        RECT 2316.3400 1906.3800 2317.9400 1906.8600 ;
        RECT 2316.3400 1911.8200 2317.9400 1912.3000 ;
        RECT 2316.3400 1955.3400 2317.9400 1955.8200 ;
        RECT 2361.3400 1955.3400 2362.9400 1955.8200 ;
        RECT 2376.8800 1955.3400 2378.4800 1955.8200 ;
        RECT 2271.3400 1987.9800 2272.9400 1988.4600 ;
        RECT 2271.3400 1993.4200 2272.9400 1993.9000 ;
        RECT 2271.3400 1998.8600 2272.9400 1999.3400 ;
        RECT 2226.3400 1987.9800 2227.9400 1988.4600 ;
        RECT 2226.3400 1993.4200 2227.9400 1993.9000 ;
        RECT 2226.3400 1998.8600 2227.9400 1999.3400 ;
        RECT 2271.3400 1971.6600 2272.9400 1972.1400 ;
        RECT 2271.3400 1977.1000 2272.9400 1977.5800 ;
        RECT 2271.3400 1960.7800 2272.9400 1961.2600 ;
        RECT 2271.3400 1966.2200 2272.9400 1966.7000 ;
        RECT 2226.3400 1971.6600 2227.9400 1972.1400 ;
        RECT 2226.3400 1977.1000 2227.9400 1977.5800 ;
        RECT 2226.3400 1960.7800 2227.9400 1961.2600 ;
        RECT 2226.3400 1966.2200 2227.9400 1966.7000 ;
        RECT 2226.3400 1982.5400 2227.9400 1983.0200 ;
        RECT 2271.3400 1982.5400 2272.9400 1983.0200 ;
        RECT 2174.1800 1998.8600 2175.7800 1999.3400 ;
        RECT 2181.3400 1998.8600 2182.9400 1999.3400 ;
        RECT 2181.3400 1987.9800 2182.9400 1988.4600 ;
        RECT 2181.3400 1993.4200 2182.9400 1993.9000 ;
        RECT 2174.1800 1987.9800 2175.7800 1988.4600 ;
        RECT 2174.1800 1993.4200 2175.7800 1993.9000 ;
        RECT 2181.3400 1971.6600 2182.9400 1972.1400 ;
        RECT 2181.3400 1977.1000 2182.9400 1977.5800 ;
        RECT 2174.1800 1971.6600 2175.7800 1972.1400 ;
        RECT 2174.1800 1977.1000 2175.7800 1977.5800 ;
        RECT 2181.3400 1960.7800 2182.9400 1961.2600 ;
        RECT 2181.3400 1966.2200 2182.9400 1966.7000 ;
        RECT 2174.1800 1960.7800 2175.7800 1961.2600 ;
        RECT 2174.1800 1966.2200 2175.7800 1966.7000 ;
        RECT 2174.1800 1982.5400 2175.7800 1983.0200 ;
        RECT 2181.3400 1982.5400 2182.9400 1983.0200 ;
        RECT 2271.3400 1944.4600 2272.9400 1944.9400 ;
        RECT 2271.3400 1949.9000 2272.9400 1950.3800 ;
        RECT 2271.3400 1928.1400 2272.9400 1928.6200 ;
        RECT 2271.3400 1933.5800 2272.9400 1934.0600 ;
        RECT 2271.3400 1939.0200 2272.9400 1939.5000 ;
        RECT 2226.3400 1944.4600 2227.9400 1944.9400 ;
        RECT 2226.3400 1949.9000 2227.9400 1950.3800 ;
        RECT 2226.3400 1928.1400 2227.9400 1928.6200 ;
        RECT 2226.3400 1933.5800 2227.9400 1934.0600 ;
        RECT 2226.3400 1939.0200 2227.9400 1939.5000 ;
        RECT 2271.3400 1917.2600 2272.9400 1917.7400 ;
        RECT 2271.3400 1922.7000 2272.9400 1923.1800 ;
        RECT 2271.3400 1900.9400 2272.9400 1901.4200 ;
        RECT 2271.3400 1906.3800 2272.9400 1906.8600 ;
        RECT 2271.3400 1911.8200 2272.9400 1912.3000 ;
        RECT 2226.3400 1917.2600 2227.9400 1917.7400 ;
        RECT 2226.3400 1922.7000 2227.9400 1923.1800 ;
        RECT 2226.3400 1900.9400 2227.9400 1901.4200 ;
        RECT 2226.3400 1906.3800 2227.9400 1906.8600 ;
        RECT 2226.3400 1911.8200 2227.9400 1912.3000 ;
        RECT 2181.3400 1944.4600 2182.9400 1944.9400 ;
        RECT 2181.3400 1949.9000 2182.9400 1950.3800 ;
        RECT 2174.1800 1944.4600 2175.7800 1944.9400 ;
        RECT 2174.1800 1949.9000 2175.7800 1950.3800 ;
        RECT 2181.3400 1928.1400 2182.9400 1928.6200 ;
        RECT 2181.3400 1933.5800 2182.9400 1934.0600 ;
        RECT 2181.3400 1939.0200 2182.9400 1939.5000 ;
        RECT 2174.1800 1928.1400 2175.7800 1928.6200 ;
        RECT 2174.1800 1933.5800 2175.7800 1934.0600 ;
        RECT 2174.1800 1939.0200 2175.7800 1939.5000 ;
        RECT 2181.3400 1917.2600 2182.9400 1917.7400 ;
        RECT 2181.3400 1922.7000 2182.9400 1923.1800 ;
        RECT 2174.1800 1917.2600 2175.7800 1917.7400 ;
        RECT 2174.1800 1922.7000 2175.7800 1923.1800 ;
        RECT 2181.3400 1900.9400 2182.9400 1901.4200 ;
        RECT 2181.3400 1906.3800 2182.9400 1906.8600 ;
        RECT 2181.3400 1911.8200 2182.9400 1912.3000 ;
        RECT 2174.1800 1900.9400 2175.7800 1901.4200 ;
        RECT 2174.1800 1906.3800 2175.7800 1906.8600 ;
        RECT 2174.1800 1911.8200 2175.7800 1912.3000 ;
        RECT 2174.1800 1955.3400 2175.7800 1955.8200 ;
        RECT 2181.3400 1955.3400 2182.9400 1955.8200 ;
        RECT 2226.3400 1955.3400 2227.9400 1955.8200 ;
        RECT 2271.3400 1955.3400 2272.9400 1955.8200 ;
        RECT 2376.8800 1890.0600 2378.4800 1890.5400 ;
        RECT 2376.8800 1895.5000 2378.4800 1895.9800 ;
        RECT 2361.3400 1890.0600 2362.9400 1890.5400 ;
        RECT 2361.3400 1895.5000 2362.9400 1895.9800 ;
        RECT 2376.8800 1873.7400 2378.4800 1874.2200 ;
        RECT 2376.8800 1879.1800 2378.4800 1879.6600 ;
        RECT 2376.8800 1884.6200 2378.4800 1885.1000 ;
        RECT 2361.3400 1873.7400 2362.9400 1874.2200 ;
        RECT 2361.3400 1879.1800 2362.9400 1879.6600 ;
        RECT 2361.3400 1884.6200 2362.9400 1885.1000 ;
        RECT 2376.8800 1862.8600 2378.4800 1863.3400 ;
        RECT 2376.8800 1868.3000 2378.4800 1868.7800 ;
        RECT 2361.3400 1862.8600 2362.9400 1863.3400 ;
        RECT 2361.3400 1868.3000 2362.9400 1868.7800 ;
        RECT 2376.8800 1846.5400 2378.4800 1847.0200 ;
        RECT 2376.8800 1851.9800 2378.4800 1852.4600 ;
        RECT 2376.8800 1857.4200 2378.4800 1857.9000 ;
        RECT 2361.3400 1846.5400 2362.9400 1847.0200 ;
        RECT 2361.3400 1851.9800 2362.9400 1852.4600 ;
        RECT 2361.3400 1857.4200 2362.9400 1857.9000 ;
        RECT 2316.3400 1890.0600 2317.9400 1890.5400 ;
        RECT 2316.3400 1895.5000 2317.9400 1895.9800 ;
        RECT 2316.3400 1873.7400 2317.9400 1874.2200 ;
        RECT 2316.3400 1879.1800 2317.9400 1879.6600 ;
        RECT 2316.3400 1884.6200 2317.9400 1885.1000 ;
        RECT 2316.3400 1862.8600 2317.9400 1863.3400 ;
        RECT 2316.3400 1868.3000 2317.9400 1868.7800 ;
        RECT 2316.3400 1846.5400 2317.9400 1847.0200 ;
        RECT 2316.3400 1851.9800 2317.9400 1852.4600 ;
        RECT 2316.3400 1857.4200 2317.9400 1857.9000 ;
        RECT 2376.8800 1835.6600 2378.4800 1836.1400 ;
        RECT 2376.8800 1841.1000 2378.4800 1841.5800 ;
        RECT 2361.3400 1835.6600 2362.9400 1836.1400 ;
        RECT 2361.3400 1841.1000 2362.9400 1841.5800 ;
        RECT 2376.8800 1819.3400 2378.4800 1819.8200 ;
        RECT 2376.8800 1824.7800 2378.4800 1825.2600 ;
        RECT 2376.8800 1830.2200 2378.4800 1830.7000 ;
        RECT 2361.3400 1819.3400 2362.9400 1819.8200 ;
        RECT 2361.3400 1824.7800 2362.9400 1825.2600 ;
        RECT 2361.3400 1830.2200 2362.9400 1830.7000 ;
        RECT 2376.8800 1808.4600 2378.4800 1808.9400 ;
        RECT 2376.8800 1813.9000 2378.4800 1814.3800 ;
        RECT 2361.3400 1808.4600 2362.9400 1808.9400 ;
        RECT 2361.3400 1813.9000 2362.9400 1814.3800 ;
        RECT 2361.3400 1803.0200 2362.9400 1803.5000 ;
        RECT 2376.8800 1803.0200 2378.4800 1803.5000 ;
        RECT 2316.3400 1835.6600 2317.9400 1836.1400 ;
        RECT 2316.3400 1841.1000 2317.9400 1841.5800 ;
        RECT 2316.3400 1819.3400 2317.9400 1819.8200 ;
        RECT 2316.3400 1824.7800 2317.9400 1825.2600 ;
        RECT 2316.3400 1830.2200 2317.9400 1830.7000 ;
        RECT 2316.3400 1808.4600 2317.9400 1808.9400 ;
        RECT 2316.3400 1813.9000 2317.9400 1814.3800 ;
        RECT 2316.3400 1803.0200 2317.9400 1803.5000 ;
        RECT 2271.3400 1890.0600 2272.9400 1890.5400 ;
        RECT 2271.3400 1895.5000 2272.9400 1895.9800 ;
        RECT 2271.3400 1873.7400 2272.9400 1874.2200 ;
        RECT 2271.3400 1879.1800 2272.9400 1879.6600 ;
        RECT 2271.3400 1884.6200 2272.9400 1885.1000 ;
        RECT 2226.3400 1890.0600 2227.9400 1890.5400 ;
        RECT 2226.3400 1895.5000 2227.9400 1895.9800 ;
        RECT 2226.3400 1873.7400 2227.9400 1874.2200 ;
        RECT 2226.3400 1879.1800 2227.9400 1879.6600 ;
        RECT 2226.3400 1884.6200 2227.9400 1885.1000 ;
        RECT 2271.3400 1862.8600 2272.9400 1863.3400 ;
        RECT 2271.3400 1868.3000 2272.9400 1868.7800 ;
        RECT 2271.3400 1846.5400 2272.9400 1847.0200 ;
        RECT 2271.3400 1851.9800 2272.9400 1852.4600 ;
        RECT 2271.3400 1857.4200 2272.9400 1857.9000 ;
        RECT 2226.3400 1862.8600 2227.9400 1863.3400 ;
        RECT 2226.3400 1868.3000 2227.9400 1868.7800 ;
        RECT 2226.3400 1846.5400 2227.9400 1847.0200 ;
        RECT 2226.3400 1851.9800 2227.9400 1852.4600 ;
        RECT 2226.3400 1857.4200 2227.9400 1857.9000 ;
        RECT 2181.3400 1890.0600 2182.9400 1890.5400 ;
        RECT 2181.3400 1895.5000 2182.9400 1895.9800 ;
        RECT 2174.1800 1890.0600 2175.7800 1890.5400 ;
        RECT 2174.1800 1895.5000 2175.7800 1895.9800 ;
        RECT 2181.3400 1873.7400 2182.9400 1874.2200 ;
        RECT 2181.3400 1879.1800 2182.9400 1879.6600 ;
        RECT 2181.3400 1884.6200 2182.9400 1885.1000 ;
        RECT 2174.1800 1873.7400 2175.7800 1874.2200 ;
        RECT 2174.1800 1879.1800 2175.7800 1879.6600 ;
        RECT 2174.1800 1884.6200 2175.7800 1885.1000 ;
        RECT 2181.3400 1862.8600 2182.9400 1863.3400 ;
        RECT 2181.3400 1868.3000 2182.9400 1868.7800 ;
        RECT 2174.1800 1862.8600 2175.7800 1863.3400 ;
        RECT 2174.1800 1868.3000 2175.7800 1868.7800 ;
        RECT 2181.3400 1846.5400 2182.9400 1847.0200 ;
        RECT 2181.3400 1851.9800 2182.9400 1852.4600 ;
        RECT 2181.3400 1857.4200 2182.9400 1857.9000 ;
        RECT 2174.1800 1846.5400 2175.7800 1847.0200 ;
        RECT 2174.1800 1851.9800 2175.7800 1852.4600 ;
        RECT 2174.1800 1857.4200 2175.7800 1857.9000 ;
        RECT 2271.3400 1835.6600 2272.9400 1836.1400 ;
        RECT 2271.3400 1841.1000 2272.9400 1841.5800 ;
        RECT 2271.3400 1819.3400 2272.9400 1819.8200 ;
        RECT 2271.3400 1824.7800 2272.9400 1825.2600 ;
        RECT 2271.3400 1830.2200 2272.9400 1830.7000 ;
        RECT 2226.3400 1835.6600 2227.9400 1836.1400 ;
        RECT 2226.3400 1841.1000 2227.9400 1841.5800 ;
        RECT 2226.3400 1819.3400 2227.9400 1819.8200 ;
        RECT 2226.3400 1824.7800 2227.9400 1825.2600 ;
        RECT 2226.3400 1830.2200 2227.9400 1830.7000 ;
        RECT 2271.3400 1813.9000 2272.9400 1814.3800 ;
        RECT 2271.3400 1808.4600 2272.9400 1808.9400 ;
        RECT 2271.3400 1803.0200 2272.9400 1803.5000 ;
        RECT 2226.3400 1813.9000 2227.9400 1814.3800 ;
        RECT 2226.3400 1808.4600 2227.9400 1808.9400 ;
        RECT 2226.3400 1803.0200 2227.9400 1803.5000 ;
        RECT 2181.3400 1835.6600 2182.9400 1836.1400 ;
        RECT 2181.3400 1841.1000 2182.9400 1841.5800 ;
        RECT 2174.1800 1835.6600 2175.7800 1836.1400 ;
        RECT 2174.1800 1841.1000 2175.7800 1841.5800 ;
        RECT 2181.3400 1819.3400 2182.9400 1819.8200 ;
        RECT 2181.3400 1824.7800 2182.9400 1825.2600 ;
        RECT 2181.3400 1830.2200 2182.9400 1830.7000 ;
        RECT 2174.1800 1819.3400 2175.7800 1819.8200 ;
        RECT 2174.1800 1824.7800 2175.7800 1825.2600 ;
        RECT 2174.1800 1830.2200 2175.7800 1830.7000 ;
        RECT 2181.3400 1808.4600 2182.9400 1808.9400 ;
        RECT 2181.3400 1813.9000 2182.9400 1814.3800 ;
        RECT 2174.1800 1808.4600 2175.7800 1808.9400 ;
        RECT 2174.1800 1813.9000 2175.7800 1814.3800 ;
        RECT 2174.1800 1803.0200 2175.7800 1803.5000 ;
        RECT 2181.3400 1803.0200 2182.9400 1803.5000 ;
        RECT 2171.2200 2005.2100 2381.4400 2006.8100 ;
        RECT 2171.2200 1793.5100 2381.4400 1795.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1790.6800 2175.7800 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 2008.7200 2175.7800 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1790.6800 2378.4800 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 2008.7200 2378.4800 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1793.5100 2172.8200 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1793.5100 2381.4400 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2005.2100 2172.8200 2006.8100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2005.2100 2381.4400 2006.8100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 1563.8700 2362.9400 1777.1700 ;
        RECT 2316.3400 1563.8700 2317.9400 1777.1700 ;
        RECT 2271.3400 1563.8700 2272.9400 1777.1700 ;
        RECT 2226.3400 1563.8700 2227.9400 1777.1700 ;
        RECT 2181.3400 1563.8700 2182.9400 1777.1700 ;
        RECT 2376.8800 1561.0400 2378.4800 1780.6800 ;
        RECT 2174.1800 1561.0400 2175.7800 1780.6800 ;
      LAYER met3 ;
        RECT 2361.3400 1769.2200 2362.9400 1769.7000 ;
        RECT 2376.8800 1769.2200 2378.4800 1769.7000 ;
        RECT 2376.8800 1758.3400 2378.4800 1758.8200 ;
        RECT 2376.8800 1763.7800 2378.4800 1764.2600 ;
        RECT 2361.3400 1758.3400 2362.9400 1758.8200 ;
        RECT 2361.3400 1763.7800 2362.9400 1764.2600 ;
        RECT 2376.8800 1742.0200 2378.4800 1742.5000 ;
        RECT 2376.8800 1747.4600 2378.4800 1747.9400 ;
        RECT 2361.3400 1742.0200 2362.9400 1742.5000 ;
        RECT 2361.3400 1747.4600 2362.9400 1747.9400 ;
        RECT 2376.8800 1731.1400 2378.4800 1731.6200 ;
        RECT 2376.8800 1736.5800 2378.4800 1737.0600 ;
        RECT 2361.3400 1731.1400 2362.9400 1731.6200 ;
        RECT 2361.3400 1736.5800 2362.9400 1737.0600 ;
        RECT 2361.3400 1752.9000 2362.9400 1753.3800 ;
        RECT 2376.8800 1752.9000 2378.4800 1753.3800 ;
        RECT 2316.3400 1758.3400 2317.9400 1758.8200 ;
        RECT 2316.3400 1763.7800 2317.9400 1764.2600 ;
        RECT 2316.3400 1769.2200 2317.9400 1769.7000 ;
        RECT 2316.3400 1742.0200 2317.9400 1742.5000 ;
        RECT 2316.3400 1747.4600 2317.9400 1747.9400 ;
        RECT 2316.3400 1736.5800 2317.9400 1737.0600 ;
        RECT 2316.3400 1731.1400 2317.9400 1731.6200 ;
        RECT 2316.3400 1752.9000 2317.9400 1753.3800 ;
        RECT 2376.8800 1714.8200 2378.4800 1715.3000 ;
        RECT 2376.8800 1720.2600 2378.4800 1720.7400 ;
        RECT 2361.3400 1714.8200 2362.9400 1715.3000 ;
        RECT 2361.3400 1720.2600 2362.9400 1720.7400 ;
        RECT 2376.8800 1698.5000 2378.4800 1698.9800 ;
        RECT 2376.8800 1703.9400 2378.4800 1704.4200 ;
        RECT 2376.8800 1709.3800 2378.4800 1709.8600 ;
        RECT 2361.3400 1698.5000 2362.9400 1698.9800 ;
        RECT 2361.3400 1703.9400 2362.9400 1704.4200 ;
        RECT 2361.3400 1709.3800 2362.9400 1709.8600 ;
        RECT 2376.8800 1687.6200 2378.4800 1688.1000 ;
        RECT 2376.8800 1693.0600 2378.4800 1693.5400 ;
        RECT 2361.3400 1687.6200 2362.9400 1688.1000 ;
        RECT 2361.3400 1693.0600 2362.9400 1693.5400 ;
        RECT 2376.8800 1671.3000 2378.4800 1671.7800 ;
        RECT 2376.8800 1676.7400 2378.4800 1677.2200 ;
        RECT 2376.8800 1682.1800 2378.4800 1682.6600 ;
        RECT 2361.3400 1671.3000 2362.9400 1671.7800 ;
        RECT 2361.3400 1676.7400 2362.9400 1677.2200 ;
        RECT 2361.3400 1682.1800 2362.9400 1682.6600 ;
        RECT 2316.3400 1714.8200 2317.9400 1715.3000 ;
        RECT 2316.3400 1720.2600 2317.9400 1720.7400 ;
        RECT 2316.3400 1698.5000 2317.9400 1698.9800 ;
        RECT 2316.3400 1703.9400 2317.9400 1704.4200 ;
        RECT 2316.3400 1709.3800 2317.9400 1709.8600 ;
        RECT 2316.3400 1687.6200 2317.9400 1688.1000 ;
        RECT 2316.3400 1693.0600 2317.9400 1693.5400 ;
        RECT 2316.3400 1671.3000 2317.9400 1671.7800 ;
        RECT 2316.3400 1676.7400 2317.9400 1677.2200 ;
        RECT 2316.3400 1682.1800 2317.9400 1682.6600 ;
        RECT 2316.3400 1725.7000 2317.9400 1726.1800 ;
        RECT 2361.3400 1725.7000 2362.9400 1726.1800 ;
        RECT 2376.8800 1725.7000 2378.4800 1726.1800 ;
        RECT 2271.3400 1758.3400 2272.9400 1758.8200 ;
        RECT 2271.3400 1763.7800 2272.9400 1764.2600 ;
        RECT 2271.3400 1769.2200 2272.9400 1769.7000 ;
        RECT 2226.3400 1758.3400 2227.9400 1758.8200 ;
        RECT 2226.3400 1763.7800 2227.9400 1764.2600 ;
        RECT 2226.3400 1769.2200 2227.9400 1769.7000 ;
        RECT 2271.3400 1742.0200 2272.9400 1742.5000 ;
        RECT 2271.3400 1747.4600 2272.9400 1747.9400 ;
        RECT 2271.3400 1731.1400 2272.9400 1731.6200 ;
        RECT 2271.3400 1736.5800 2272.9400 1737.0600 ;
        RECT 2226.3400 1742.0200 2227.9400 1742.5000 ;
        RECT 2226.3400 1747.4600 2227.9400 1747.9400 ;
        RECT 2226.3400 1731.1400 2227.9400 1731.6200 ;
        RECT 2226.3400 1736.5800 2227.9400 1737.0600 ;
        RECT 2226.3400 1752.9000 2227.9400 1753.3800 ;
        RECT 2271.3400 1752.9000 2272.9400 1753.3800 ;
        RECT 2174.1800 1769.2200 2175.7800 1769.7000 ;
        RECT 2181.3400 1769.2200 2182.9400 1769.7000 ;
        RECT 2181.3400 1758.3400 2182.9400 1758.8200 ;
        RECT 2181.3400 1763.7800 2182.9400 1764.2600 ;
        RECT 2174.1800 1758.3400 2175.7800 1758.8200 ;
        RECT 2174.1800 1763.7800 2175.7800 1764.2600 ;
        RECT 2181.3400 1742.0200 2182.9400 1742.5000 ;
        RECT 2181.3400 1747.4600 2182.9400 1747.9400 ;
        RECT 2174.1800 1742.0200 2175.7800 1742.5000 ;
        RECT 2174.1800 1747.4600 2175.7800 1747.9400 ;
        RECT 2181.3400 1731.1400 2182.9400 1731.6200 ;
        RECT 2181.3400 1736.5800 2182.9400 1737.0600 ;
        RECT 2174.1800 1731.1400 2175.7800 1731.6200 ;
        RECT 2174.1800 1736.5800 2175.7800 1737.0600 ;
        RECT 2174.1800 1752.9000 2175.7800 1753.3800 ;
        RECT 2181.3400 1752.9000 2182.9400 1753.3800 ;
        RECT 2271.3400 1714.8200 2272.9400 1715.3000 ;
        RECT 2271.3400 1720.2600 2272.9400 1720.7400 ;
        RECT 2271.3400 1698.5000 2272.9400 1698.9800 ;
        RECT 2271.3400 1703.9400 2272.9400 1704.4200 ;
        RECT 2271.3400 1709.3800 2272.9400 1709.8600 ;
        RECT 2226.3400 1714.8200 2227.9400 1715.3000 ;
        RECT 2226.3400 1720.2600 2227.9400 1720.7400 ;
        RECT 2226.3400 1698.5000 2227.9400 1698.9800 ;
        RECT 2226.3400 1703.9400 2227.9400 1704.4200 ;
        RECT 2226.3400 1709.3800 2227.9400 1709.8600 ;
        RECT 2271.3400 1687.6200 2272.9400 1688.1000 ;
        RECT 2271.3400 1693.0600 2272.9400 1693.5400 ;
        RECT 2271.3400 1671.3000 2272.9400 1671.7800 ;
        RECT 2271.3400 1676.7400 2272.9400 1677.2200 ;
        RECT 2271.3400 1682.1800 2272.9400 1682.6600 ;
        RECT 2226.3400 1687.6200 2227.9400 1688.1000 ;
        RECT 2226.3400 1693.0600 2227.9400 1693.5400 ;
        RECT 2226.3400 1671.3000 2227.9400 1671.7800 ;
        RECT 2226.3400 1676.7400 2227.9400 1677.2200 ;
        RECT 2226.3400 1682.1800 2227.9400 1682.6600 ;
        RECT 2181.3400 1714.8200 2182.9400 1715.3000 ;
        RECT 2181.3400 1720.2600 2182.9400 1720.7400 ;
        RECT 2174.1800 1714.8200 2175.7800 1715.3000 ;
        RECT 2174.1800 1720.2600 2175.7800 1720.7400 ;
        RECT 2181.3400 1698.5000 2182.9400 1698.9800 ;
        RECT 2181.3400 1703.9400 2182.9400 1704.4200 ;
        RECT 2181.3400 1709.3800 2182.9400 1709.8600 ;
        RECT 2174.1800 1698.5000 2175.7800 1698.9800 ;
        RECT 2174.1800 1703.9400 2175.7800 1704.4200 ;
        RECT 2174.1800 1709.3800 2175.7800 1709.8600 ;
        RECT 2181.3400 1687.6200 2182.9400 1688.1000 ;
        RECT 2181.3400 1693.0600 2182.9400 1693.5400 ;
        RECT 2174.1800 1687.6200 2175.7800 1688.1000 ;
        RECT 2174.1800 1693.0600 2175.7800 1693.5400 ;
        RECT 2181.3400 1671.3000 2182.9400 1671.7800 ;
        RECT 2181.3400 1676.7400 2182.9400 1677.2200 ;
        RECT 2181.3400 1682.1800 2182.9400 1682.6600 ;
        RECT 2174.1800 1671.3000 2175.7800 1671.7800 ;
        RECT 2174.1800 1676.7400 2175.7800 1677.2200 ;
        RECT 2174.1800 1682.1800 2175.7800 1682.6600 ;
        RECT 2174.1800 1725.7000 2175.7800 1726.1800 ;
        RECT 2181.3400 1725.7000 2182.9400 1726.1800 ;
        RECT 2226.3400 1725.7000 2227.9400 1726.1800 ;
        RECT 2271.3400 1725.7000 2272.9400 1726.1800 ;
        RECT 2376.8800 1660.4200 2378.4800 1660.9000 ;
        RECT 2376.8800 1665.8600 2378.4800 1666.3400 ;
        RECT 2361.3400 1660.4200 2362.9400 1660.9000 ;
        RECT 2361.3400 1665.8600 2362.9400 1666.3400 ;
        RECT 2376.8800 1644.1000 2378.4800 1644.5800 ;
        RECT 2376.8800 1649.5400 2378.4800 1650.0200 ;
        RECT 2376.8800 1654.9800 2378.4800 1655.4600 ;
        RECT 2361.3400 1644.1000 2362.9400 1644.5800 ;
        RECT 2361.3400 1649.5400 2362.9400 1650.0200 ;
        RECT 2361.3400 1654.9800 2362.9400 1655.4600 ;
        RECT 2376.8800 1633.2200 2378.4800 1633.7000 ;
        RECT 2376.8800 1638.6600 2378.4800 1639.1400 ;
        RECT 2361.3400 1633.2200 2362.9400 1633.7000 ;
        RECT 2361.3400 1638.6600 2362.9400 1639.1400 ;
        RECT 2376.8800 1616.9000 2378.4800 1617.3800 ;
        RECT 2376.8800 1622.3400 2378.4800 1622.8200 ;
        RECT 2376.8800 1627.7800 2378.4800 1628.2600 ;
        RECT 2361.3400 1616.9000 2362.9400 1617.3800 ;
        RECT 2361.3400 1622.3400 2362.9400 1622.8200 ;
        RECT 2361.3400 1627.7800 2362.9400 1628.2600 ;
        RECT 2316.3400 1660.4200 2317.9400 1660.9000 ;
        RECT 2316.3400 1665.8600 2317.9400 1666.3400 ;
        RECT 2316.3400 1644.1000 2317.9400 1644.5800 ;
        RECT 2316.3400 1649.5400 2317.9400 1650.0200 ;
        RECT 2316.3400 1654.9800 2317.9400 1655.4600 ;
        RECT 2316.3400 1633.2200 2317.9400 1633.7000 ;
        RECT 2316.3400 1638.6600 2317.9400 1639.1400 ;
        RECT 2316.3400 1616.9000 2317.9400 1617.3800 ;
        RECT 2316.3400 1622.3400 2317.9400 1622.8200 ;
        RECT 2316.3400 1627.7800 2317.9400 1628.2600 ;
        RECT 2376.8800 1606.0200 2378.4800 1606.5000 ;
        RECT 2376.8800 1611.4600 2378.4800 1611.9400 ;
        RECT 2361.3400 1606.0200 2362.9400 1606.5000 ;
        RECT 2361.3400 1611.4600 2362.9400 1611.9400 ;
        RECT 2376.8800 1589.7000 2378.4800 1590.1800 ;
        RECT 2376.8800 1595.1400 2378.4800 1595.6200 ;
        RECT 2376.8800 1600.5800 2378.4800 1601.0600 ;
        RECT 2361.3400 1589.7000 2362.9400 1590.1800 ;
        RECT 2361.3400 1595.1400 2362.9400 1595.6200 ;
        RECT 2361.3400 1600.5800 2362.9400 1601.0600 ;
        RECT 2376.8800 1578.8200 2378.4800 1579.3000 ;
        RECT 2376.8800 1584.2600 2378.4800 1584.7400 ;
        RECT 2361.3400 1578.8200 2362.9400 1579.3000 ;
        RECT 2361.3400 1584.2600 2362.9400 1584.7400 ;
        RECT 2361.3400 1573.3800 2362.9400 1573.8600 ;
        RECT 2376.8800 1573.3800 2378.4800 1573.8600 ;
        RECT 2316.3400 1606.0200 2317.9400 1606.5000 ;
        RECT 2316.3400 1611.4600 2317.9400 1611.9400 ;
        RECT 2316.3400 1589.7000 2317.9400 1590.1800 ;
        RECT 2316.3400 1595.1400 2317.9400 1595.6200 ;
        RECT 2316.3400 1600.5800 2317.9400 1601.0600 ;
        RECT 2316.3400 1578.8200 2317.9400 1579.3000 ;
        RECT 2316.3400 1584.2600 2317.9400 1584.7400 ;
        RECT 2316.3400 1573.3800 2317.9400 1573.8600 ;
        RECT 2271.3400 1660.4200 2272.9400 1660.9000 ;
        RECT 2271.3400 1665.8600 2272.9400 1666.3400 ;
        RECT 2271.3400 1644.1000 2272.9400 1644.5800 ;
        RECT 2271.3400 1649.5400 2272.9400 1650.0200 ;
        RECT 2271.3400 1654.9800 2272.9400 1655.4600 ;
        RECT 2226.3400 1660.4200 2227.9400 1660.9000 ;
        RECT 2226.3400 1665.8600 2227.9400 1666.3400 ;
        RECT 2226.3400 1644.1000 2227.9400 1644.5800 ;
        RECT 2226.3400 1649.5400 2227.9400 1650.0200 ;
        RECT 2226.3400 1654.9800 2227.9400 1655.4600 ;
        RECT 2271.3400 1633.2200 2272.9400 1633.7000 ;
        RECT 2271.3400 1638.6600 2272.9400 1639.1400 ;
        RECT 2271.3400 1616.9000 2272.9400 1617.3800 ;
        RECT 2271.3400 1622.3400 2272.9400 1622.8200 ;
        RECT 2271.3400 1627.7800 2272.9400 1628.2600 ;
        RECT 2226.3400 1633.2200 2227.9400 1633.7000 ;
        RECT 2226.3400 1638.6600 2227.9400 1639.1400 ;
        RECT 2226.3400 1616.9000 2227.9400 1617.3800 ;
        RECT 2226.3400 1622.3400 2227.9400 1622.8200 ;
        RECT 2226.3400 1627.7800 2227.9400 1628.2600 ;
        RECT 2181.3400 1660.4200 2182.9400 1660.9000 ;
        RECT 2181.3400 1665.8600 2182.9400 1666.3400 ;
        RECT 2174.1800 1660.4200 2175.7800 1660.9000 ;
        RECT 2174.1800 1665.8600 2175.7800 1666.3400 ;
        RECT 2181.3400 1644.1000 2182.9400 1644.5800 ;
        RECT 2181.3400 1649.5400 2182.9400 1650.0200 ;
        RECT 2181.3400 1654.9800 2182.9400 1655.4600 ;
        RECT 2174.1800 1644.1000 2175.7800 1644.5800 ;
        RECT 2174.1800 1649.5400 2175.7800 1650.0200 ;
        RECT 2174.1800 1654.9800 2175.7800 1655.4600 ;
        RECT 2181.3400 1633.2200 2182.9400 1633.7000 ;
        RECT 2181.3400 1638.6600 2182.9400 1639.1400 ;
        RECT 2174.1800 1633.2200 2175.7800 1633.7000 ;
        RECT 2174.1800 1638.6600 2175.7800 1639.1400 ;
        RECT 2181.3400 1616.9000 2182.9400 1617.3800 ;
        RECT 2181.3400 1622.3400 2182.9400 1622.8200 ;
        RECT 2181.3400 1627.7800 2182.9400 1628.2600 ;
        RECT 2174.1800 1616.9000 2175.7800 1617.3800 ;
        RECT 2174.1800 1622.3400 2175.7800 1622.8200 ;
        RECT 2174.1800 1627.7800 2175.7800 1628.2600 ;
        RECT 2271.3400 1606.0200 2272.9400 1606.5000 ;
        RECT 2271.3400 1611.4600 2272.9400 1611.9400 ;
        RECT 2271.3400 1589.7000 2272.9400 1590.1800 ;
        RECT 2271.3400 1595.1400 2272.9400 1595.6200 ;
        RECT 2271.3400 1600.5800 2272.9400 1601.0600 ;
        RECT 2226.3400 1606.0200 2227.9400 1606.5000 ;
        RECT 2226.3400 1611.4600 2227.9400 1611.9400 ;
        RECT 2226.3400 1589.7000 2227.9400 1590.1800 ;
        RECT 2226.3400 1595.1400 2227.9400 1595.6200 ;
        RECT 2226.3400 1600.5800 2227.9400 1601.0600 ;
        RECT 2271.3400 1584.2600 2272.9400 1584.7400 ;
        RECT 2271.3400 1578.8200 2272.9400 1579.3000 ;
        RECT 2271.3400 1573.3800 2272.9400 1573.8600 ;
        RECT 2226.3400 1584.2600 2227.9400 1584.7400 ;
        RECT 2226.3400 1578.8200 2227.9400 1579.3000 ;
        RECT 2226.3400 1573.3800 2227.9400 1573.8600 ;
        RECT 2181.3400 1606.0200 2182.9400 1606.5000 ;
        RECT 2181.3400 1611.4600 2182.9400 1611.9400 ;
        RECT 2174.1800 1606.0200 2175.7800 1606.5000 ;
        RECT 2174.1800 1611.4600 2175.7800 1611.9400 ;
        RECT 2181.3400 1589.7000 2182.9400 1590.1800 ;
        RECT 2181.3400 1595.1400 2182.9400 1595.6200 ;
        RECT 2181.3400 1600.5800 2182.9400 1601.0600 ;
        RECT 2174.1800 1589.7000 2175.7800 1590.1800 ;
        RECT 2174.1800 1595.1400 2175.7800 1595.6200 ;
        RECT 2174.1800 1600.5800 2175.7800 1601.0600 ;
        RECT 2181.3400 1578.8200 2182.9400 1579.3000 ;
        RECT 2181.3400 1584.2600 2182.9400 1584.7400 ;
        RECT 2174.1800 1578.8200 2175.7800 1579.3000 ;
        RECT 2174.1800 1584.2600 2175.7800 1584.7400 ;
        RECT 2174.1800 1573.3800 2175.7800 1573.8600 ;
        RECT 2181.3400 1573.3800 2182.9400 1573.8600 ;
        RECT 2171.2200 1775.5700 2381.4400 1777.1700 ;
        RECT 2171.2200 1563.8700 2381.4400 1565.4700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1561.0400 2175.7800 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1779.0800 2175.7800 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1561.0400 2378.4800 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1779.0800 2378.4800 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1563.8700 2172.8200 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1563.8700 2381.4400 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1775.5700 2172.8200 1777.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1775.5700 2381.4400 1777.1700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 1334.2300 2362.9400 1547.5300 ;
        RECT 2316.3400 1334.2300 2317.9400 1547.5300 ;
        RECT 2271.3400 1334.2300 2272.9400 1547.5300 ;
        RECT 2226.3400 1334.2300 2227.9400 1547.5300 ;
        RECT 2181.3400 1334.2300 2182.9400 1547.5300 ;
        RECT 2376.8800 1331.4000 2378.4800 1551.0400 ;
        RECT 2174.1800 1331.4000 2175.7800 1551.0400 ;
      LAYER met3 ;
        RECT 2361.3400 1539.5800 2362.9400 1540.0600 ;
        RECT 2376.8800 1539.5800 2378.4800 1540.0600 ;
        RECT 2376.8800 1528.7000 2378.4800 1529.1800 ;
        RECT 2376.8800 1534.1400 2378.4800 1534.6200 ;
        RECT 2361.3400 1528.7000 2362.9400 1529.1800 ;
        RECT 2361.3400 1534.1400 2362.9400 1534.6200 ;
        RECT 2376.8800 1512.3800 2378.4800 1512.8600 ;
        RECT 2376.8800 1517.8200 2378.4800 1518.3000 ;
        RECT 2361.3400 1512.3800 2362.9400 1512.8600 ;
        RECT 2361.3400 1517.8200 2362.9400 1518.3000 ;
        RECT 2376.8800 1501.5000 2378.4800 1501.9800 ;
        RECT 2376.8800 1506.9400 2378.4800 1507.4200 ;
        RECT 2361.3400 1501.5000 2362.9400 1501.9800 ;
        RECT 2361.3400 1506.9400 2362.9400 1507.4200 ;
        RECT 2361.3400 1523.2600 2362.9400 1523.7400 ;
        RECT 2376.8800 1523.2600 2378.4800 1523.7400 ;
        RECT 2316.3400 1528.7000 2317.9400 1529.1800 ;
        RECT 2316.3400 1534.1400 2317.9400 1534.6200 ;
        RECT 2316.3400 1539.5800 2317.9400 1540.0600 ;
        RECT 2316.3400 1512.3800 2317.9400 1512.8600 ;
        RECT 2316.3400 1517.8200 2317.9400 1518.3000 ;
        RECT 2316.3400 1506.9400 2317.9400 1507.4200 ;
        RECT 2316.3400 1501.5000 2317.9400 1501.9800 ;
        RECT 2316.3400 1523.2600 2317.9400 1523.7400 ;
        RECT 2376.8800 1485.1800 2378.4800 1485.6600 ;
        RECT 2376.8800 1490.6200 2378.4800 1491.1000 ;
        RECT 2361.3400 1485.1800 2362.9400 1485.6600 ;
        RECT 2361.3400 1490.6200 2362.9400 1491.1000 ;
        RECT 2376.8800 1468.8600 2378.4800 1469.3400 ;
        RECT 2376.8800 1474.3000 2378.4800 1474.7800 ;
        RECT 2376.8800 1479.7400 2378.4800 1480.2200 ;
        RECT 2361.3400 1468.8600 2362.9400 1469.3400 ;
        RECT 2361.3400 1474.3000 2362.9400 1474.7800 ;
        RECT 2361.3400 1479.7400 2362.9400 1480.2200 ;
        RECT 2376.8800 1457.9800 2378.4800 1458.4600 ;
        RECT 2376.8800 1463.4200 2378.4800 1463.9000 ;
        RECT 2361.3400 1457.9800 2362.9400 1458.4600 ;
        RECT 2361.3400 1463.4200 2362.9400 1463.9000 ;
        RECT 2376.8800 1441.6600 2378.4800 1442.1400 ;
        RECT 2376.8800 1447.1000 2378.4800 1447.5800 ;
        RECT 2376.8800 1452.5400 2378.4800 1453.0200 ;
        RECT 2361.3400 1441.6600 2362.9400 1442.1400 ;
        RECT 2361.3400 1447.1000 2362.9400 1447.5800 ;
        RECT 2361.3400 1452.5400 2362.9400 1453.0200 ;
        RECT 2316.3400 1485.1800 2317.9400 1485.6600 ;
        RECT 2316.3400 1490.6200 2317.9400 1491.1000 ;
        RECT 2316.3400 1468.8600 2317.9400 1469.3400 ;
        RECT 2316.3400 1474.3000 2317.9400 1474.7800 ;
        RECT 2316.3400 1479.7400 2317.9400 1480.2200 ;
        RECT 2316.3400 1457.9800 2317.9400 1458.4600 ;
        RECT 2316.3400 1463.4200 2317.9400 1463.9000 ;
        RECT 2316.3400 1441.6600 2317.9400 1442.1400 ;
        RECT 2316.3400 1447.1000 2317.9400 1447.5800 ;
        RECT 2316.3400 1452.5400 2317.9400 1453.0200 ;
        RECT 2316.3400 1496.0600 2317.9400 1496.5400 ;
        RECT 2361.3400 1496.0600 2362.9400 1496.5400 ;
        RECT 2376.8800 1496.0600 2378.4800 1496.5400 ;
        RECT 2271.3400 1528.7000 2272.9400 1529.1800 ;
        RECT 2271.3400 1534.1400 2272.9400 1534.6200 ;
        RECT 2271.3400 1539.5800 2272.9400 1540.0600 ;
        RECT 2226.3400 1528.7000 2227.9400 1529.1800 ;
        RECT 2226.3400 1534.1400 2227.9400 1534.6200 ;
        RECT 2226.3400 1539.5800 2227.9400 1540.0600 ;
        RECT 2271.3400 1512.3800 2272.9400 1512.8600 ;
        RECT 2271.3400 1517.8200 2272.9400 1518.3000 ;
        RECT 2271.3400 1501.5000 2272.9400 1501.9800 ;
        RECT 2271.3400 1506.9400 2272.9400 1507.4200 ;
        RECT 2226.3400 1512.3800 2227.9400 1512.8600 ;
        RECT 2226.3400 1517.8200 2227.9400 1518.3000 ;
        RECT 2226.3400 1501.5000 2227.9400 1501.9800 ;
        RECT 2226.3400 1506.9400 2227.9400 1507.4200 ;
        RECT 2226.3400 1523.2600 2227.9400 1523.7400 ;
        RECT 2271.3400 1523.2600 2272.9400 1523.7400 ;
        RECT 2174.1800 1539.5800 2175.7800 1540.0600 ;
        RECT 2181.3400 1539.5800 2182.9400 1540.0600 ;
        RECT 2181.3400 1528.7000 2182.9400 1529.1800 ;
        RECT 2181.3400 1534.1400 2182.9400 1534.6200 ;
        RECT 2174.1800 1528.7000 2175.7800 1529.1800 ;
        RECT 2174.1800 1534.1400 2175.7800 1534.6200 ;
        RECT 2181.3400 1512.3800 2182.9400 1512.8600 ;
        RECT 2181.3400 1517.8200 2182.9400 1518.3000 ;
        RECT 2174.1800 1512.3800 2175.7800 1512.8600 ;
        RECT 2174.1800 1517.8200 2175.7800 1518.3000 ;
        RECT 2181.3400 1501.5000 2182.9400 1501.9800 ;
        RECT 2181.3400 1506.9400 2182.9400 1507.4200 ;
        RECT 2174.1800 1501.5000 2175.7800 1501.9800 ;
        RECT 2174.1800 1506.9400 2175.7800 1507.4200 ;
        RECT 2174.1800 1523.2600 2175.7800 1523.7400 ;
        RECT 2181.3400 1523.2600 2182.9400 1523.7400 ;
        RECT 2271.3400 1485.1800 2272.9400 1485.6600 ;
        RECT 2271.3400 1490.6200 2272.9400 1491.1000 ;
        RECT 2271.3400 1468.8600 2272.9400 1469.3400 ;
        RECT 2271.3400 1474.3000 2272.9400 1474.7800 ;
        RECT 2271.3400 1479.7400 2272.9400 1480.2200 ;
        RECT 2226.3400 1485.1800 2227.9400 1485.6600 ;
        RECT 2226.3400 1490.6200 2227.9400 1491.1000 ;
        RECT 2226.3400 1468.8600 2227.9400 1469.3400 ;
        RECT 2226.3400 1474.3000 2227.9400 1474.7800 ;
        RECT 2226.3400 1479.7400 2227.9400 1480.2200 ;
        RECT 2271.3400 1457.9800 2272.9400 1458.4600 ;
        RECT 2271.3400 1463.4200 2272.9400 1463.9000 ;
        RECT 2271.3400 1441.6600 2272.9400 1442.1400 ;
        RECT 2271.3400 1447.1000 2272.9400 1447.5800 ;
        RECT 2271.3400 1452.5400 2272.9400 1453.0200 ;
        RECT 2226.3400 1457.9800 2227.9400 1458.4600 ;
        RECT 2226.3400 1463.4200 2227.9400 1463.9000 ;
        RECT 2226.3400 1441.6600 2227.9400 1442.1400 ;
        RECT 2226.3400 1447.1000 2227.9400 1447.5800 ;
        RECT 2226.3400 1452.5400 2227.9400 1453.0200 ;
        RECT 2181.3400 1485.1800 2182.9400 1485.6600 ;
        RECT 2181.3400 1490.6200 2182.9400 1491.1000 ;
        RECT 2174.1800 1485.1800 2175.7800 1485.6600 ;
        RECT 2174.1800 1490.6200 2175.7800 1491.1000 ;
        RECT 2181.3400 1468.8600 2182.9400 1469.3400 ;
        RECT 2181.3400 1474.3000 2182.9400 1474.7800 ;
        RECT 2181.3400 1479.7400 2182.9400 1480.2200 ;
        RECT 2174.1800 1468.8600 2175.7800 1469.3400 ;
        RECT 2174.1800 1474.3000 2175.7800 1474.7800 ;
        RECT 2174.1800 1479.7400 2175.7800 1480.2200 ;
        RECT 2181.3400 1457.9800 2182.9400 1458.4600 ;
        RECT 2181.3400 1463.4200 2182.9400 1463.9000 ;
        RECT 2174.1800 1457.9800 2175.7800 1458.4600 ;
        RECT 2174.1800 1463.4200 2175.7800 1463.9000 ;
        RECT 2181.3400 1441.6600 2182.9400 1442.1400 ;
        RECT 2181.3400 1447.1000 2182.9400 1447.5800 ;
        RECT 2181.3400 1452.5400 2182.9400 1453.0200 ;
        RECT 2174.1800 1441.6600 2175.7800 1442.1400 ;
        RECT 2174.1800 1447.1000 2175.7800 1447.5800 ;
        RECT 2174.1800 1452.5400 2175.7800 1453.0200 ;
        RECT 2174.1800 1496.0600 2175.7800 1496.5400 ;
        RECT 2181.3400 1496.0600 2182.9400 1496.5400 ;
        RECT 2226.3400 1496.0600 2227.9400 1496.5400 ;
        RECT 2271.3400 1496.0600 2272.9400 1496.5400 ;
        RECT 2376.8800 1430.7800 2378.4800 1431.2600 ;
        RECT 2376.8800 1436.2200 2378.4800 1436.7000 ;
        RECT 2361.3400 1430.7800 2362.9400 1431.2600 ;
        RECT 2361.3400 1436.2200 2362.9400 1436.7000 ;
        RECT 2376.8800 1414.4600 2378.4800 1414.9400 ;
        RECT 2376.8800 1419.9000 2378.4800 1420.3800 ;
        RECT 2376.8800 1425.3400 2378.4800 1425.8200 ;
        RECT 2361.3400 1414.4600 2362.9400 1414.9400 ;
        RECT 2361.3400 1419.9000 2362.9400 1420.3800 ;
        RECT 2361.3400 1425.3400 2362.9400 1425.8200 ;
        RECT 2376.8800 1403.5800 2378.4800 1404.0600 ;
        RECT 2376.8800 1409.0200 2378.4800 1409.5000 ;
        RECT 2361.3400 1403.5800 2362.9400 1404.0600 ;
        RECT 2361.3400 1409.0200 2362.9400 1409.5000 ;
        RECT 2376.8800 1387.2600 2378.4800 1387.7400 ;
        RECT 2376.8800 1392.7000 2378.4800 1393.1800 ;
        RECT 2376.8800 1398.1400 2378.4800 1398.6200 ;
        RECT 2361.3400 1387.2600 2362.9400 1387.7400 ;
        RECT 2361.3400 1392.7000 2362.9400 1393.1800 ;
        RECT 2361.3400 1398.1400 2362.9400 1398.6200 ;
        RECT 2316.3400 1430.7800 2317.9400 1431.2600 ;
        RECT 2316.3400 1436.2200 2317.9400 1436.7000 ;
        RECT 2316.3400 1414.4600 2317.9400 1414.9400 ;
        RECT 2316.3400 1419.9000 2317.9400 1420.3800 ;
        RECT 2316.3400 1425.3400 2317.9400 1425.8200 ;
        RECT 2316.3400 1403.5800 2317.9400 1404.0600 ;
        RECT 2316.3400 1409.0200 2317.9400 1409.5000 ;
        RECT 2316.3400 1387.2600 2317.9400 1387.7400 ;
        RECT 2316.3400 1392.7000 2317.9400 1393.1800 ;
        RECT 2316.3400 1398.1400 2317.9400 1398.6200 ;
        RECT 2376.8800 1376.3800 2378.4800 1376.8600 ;
        RECT 2376.8800 1381.8200 2378.4800 1382.3000 ;
        RECT 2361.3400 1376.3800 2362.9400 1376.8600 ;
        RECT 2361.3400 1381.8200 2362.9400 1382.3000 ;
        RECT 2376.8800 1360.0600 2378.4800 1360.5400 ;
        RECT 2376.8800 1365.5000 2378.4800 1365.9800 ;
        RECT 2376.8800 1370.9400 2378.4800 1371.4200 ;
        RECT 2361.3400 1360.0600 2362.9400 1360.5400 ;
        RECT 2361.3400 1365.5000 2362.9400 1365.9800 ;
        RECT 2361.3400 1370.9400 2362.9400 1371.4200 ;
        RECT 2376.8800 1349.1800 2378.4800 1349.6600 ;
        RECT 2376.8800 1354.6200 2378.4800 1355.1000 ;
        RECT 2361.3400 1349.1800 2362.9400 1349.6600 ;
        RECT 2361.3400 1354.6200 2362.9400 1355.1000 ;
        RECT 2361.3400 1343.7400 2362.9400 1344.2200 ;
        RECT 2376.8800 1343.7400 2378.4800 1344.2200 ;
        RECT 2316.3400 1376.3800 2317.9400 1376.8600 ;
        RECT 2316.3400 1381.8200 2317.9400 1382.3000 ;
        RECT 2316.3400 1360.0600 2317.9400 1360.5400 ;
        RECT 2316.3400 1365.5000 2317.9400 1365.9800 ;
        RECT 2316.3400 1370.9400 2317.9400 1371.4200 ;
        RECT 2316.3400 1349.1800 2317.9400 1349.6600 ;
        RECT 2316.3400 1354.6200 2317.9400 1355.1000 ;
        RECT 2316.3400 1343.7400 2317.9400 1344.2200 ;
        RECT 2271.3400 1430.7800 2272.9400 1431.2600 ;
        RECT 2271.3400 1436.2200 2272.9400 1436.7000 ;
        RECT 2271.3400 1414.4600 2272.9400 1414.9400 ;
        RECT 2271.3400 1419.9000 2272.9400 1420.3800 ;
        RECT 2271.3400 1425.3400 2272.9400 1425.8200 ;
        RECT 2226.3400 1430.7800 2227.9400 1431.2600 ;
        RECT 2226.3400 1436.2200 2227.9400 1436.7000 ;
        RECT 2226.3400 1414.4600 2227.9400 1414.9400 ;
        RECT 2226.3400 1419.9000 2227.9400 1420.3800 ;
        RECT 2226.3400 1425.3400 2227.9400 1425.8200 ;
        RECT 2271.3400 1403.5800 2272.9400 1404.0600 ;
        RECT 2271.3400 1409.0200 2272.9400 1409.5000 ;
        RECT 2271.3400 1387.2600 2272.9400 1387.7400 ;
        RECT 2271.3400 1392.7000 2272.9400 1393.1800 ;
        RECT 2271.3400 1398.1400 2272.9400 1398.6200 ;
        RECT 2226.3400 1403.5800 2227.9400 1404.0600 ;
        RECT 2226.3400 1409.0200 2227.9400 1409.5000 ;
        RECT 2226.3400 1387.2600 2227.9400 1387.7400 ;
        RECT 2226.3400 1392.7000 2227.9400 1393.1800 ;
        RECT 2226.3400 1398.1400 2227.9400 1398.6200 ;
        RECT 2181.3400 1430.7800 2182.9400 1431.2600 ;
        RECT 2181.3400 1436.2200 2182.9400 1436.7000 ;
        RECT 2174.1800 1430.7800 2175.7800 1431.2600 ;
        RECT 2174.1800 1436.2200 2175.7800 1436.7000 ;
        RECT 2181.3400 1414.4600 2182.9400 1414.9400 ;
        RECT 2181.3400 1419.9000 2182.9400 1420.3800 ;
        RECT 2181.3400 1425.3400 2182.9400 1425.8200 ;
        RECT 2174.1800 1414.4600 2175.7800 1414.9400 ;
        RECT 2174.1800 1419.9000 2175.7800 1420.3800 ;
        RECT 2174.1800 1425.3400 2175.7800 1425.8200 ;
        RECT 2181.3400 1403.5800 2182.9400 1404.0600 ;
        RECT 2181.3400 1409.0200 2182.9400 1409.5000 ;
        RECT 2174.1800 1403.5800 2175.7800 1404.0600 ;
        RECT 2174.1800 1409.0200 2175.7800 1409.5000 ;
        RECT 2181.3400 1387.2600 2182.9400 1387.7400 ;
        RECT 2181.3400 1392.7000 2182.9400 1393.1800 ;
        RECT 2181.3400 1398.1400 2182.9400 1398.6200 ;
        RECT 2174.1800 1387.2600 2175.7800 1387.7400 ;
        RECT 2174.1800 1392.7000 2175.7800 1393.1800 ;
        RECT 2174.1800 1398.1400 2175.7800 1398.6200 ;
        RECT 2271.3400 1376.3800 2272.9400 1376.8600 ;
        RECT 2271.3400 1381.8200 2272.9400 1382.3000 ;
        RECT 2271.3400 1360.0600 2272.9400 1360.5400 ;
        RECT 2271.3400 1365.5000 2272.9400 1365.9800 ;
        RECT 2271.3400 1370.9400 2272.9400 1371.4200 ;
        RECT 2226.3400 1376.3800 2227.9400 1376.8600 ;
        RECT 2226.3400 1381.8200 2227.9400 1382.3000 ;
        RECT 2226.3400 1360.0600 2227.9400 1360.5400 ;
        RECT 2226.3400 1365.5000 2227.9400 1365.9800 ;
        RECT 2226.3400 1370.9400 2227.9400 1371.4200 ;
        RECT 2271.3400 1354.6200 2272.9400 1355.1000 ;
        RECT 2271.3400 1349.1800 2272.9400 1349.6600 ;
        RECT 2271.3400 1343.7400 2272.9400 1344.2200 ;
        RECT 2226.3400 1354.6200 2227.9400 1355.1000 ;
        RECT 2226.3400 1349.1800 2227.9400 1349.6600 ;
        RECT 2226.3400 1343.7400 2227.9400 1344.2200 ;
        RECT 2181.3400 1376.3800 2182.9400 1376.8600 ;
        RECT 2181.3400 1381.8200 2182.9400 1382.3000 ;
        RECT 2174.1800 1376.3800 2175.7800 1376.8600 ;
        RECT 2174.1800 1381.8200 2175.7800 1382.3000 ;
        RECT 2181.3400 1360.0600 2182.9400 1360.5400 ;
        RECT 2181.3400 1365.5000 2182.9400 1365.9800 ;
        RECT 2181.3400 1370.9400 2182.9400 1371.4200 ;
        RECT 2174.1800 1360.0600 2175.7800 1360.5400 ;
        RECT 2174.1800 1365.5000 2175.7800 1365.9800 ;
        RECT 2174.1800 1370.9400 2175.7800 1371.4200 ;
        RECT 2181.3400 1349.1800 2182.9400 1349.6600 ;
        RECT 2181.3400 1354.6200 2182.9400 1355.1000 ;
        RECT 2174.1800 1349.1800 2175.7800 1349.6600 ;
        RECT 2174.1800 1354.6200 2175.7800 1355.1000 ;
        RECT 2174.1800 1343.7400 2175.7800 1344.2200 ;
        RECT 2181.3400 1343.7400 2182.9400 1344.2200 ;
        RECT 2171.2200 1545.9300 2381.4400 1547.5300 ;
        RECT 2171.2200 1334.2300 2381.4400 1335.8300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1331.4000 2175.7800 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1549.4400 2175.7800 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1331.4000 2378.4800 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1549.4400 2378.4800 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1334.2300 2172.8200 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1334.2300 2381.4400 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1545.9300 2172.8200 1547.5300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1545.9300 2381.4400 1547.5300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 1104.5900 2362.9400 1317.8900 ;
        RECT 2316.3400 1104.5900 2317.9400 1317.8900 ;
        RECT 2271.3400 1104.5900 2272.9400 1317.8900 ;
        RECT 2226.3400 1104.5900 2227.9400 1317.8900 ;
        RECT 2181.3400 1104.5900 2182.9400 1317.8900 ;
        RECT 2376.8800 1101.7600 2378.4800 1321.4000 ;
        RECT 2174.1800 1101.7600 2175.7800 1321.4000 ;
      LAYER met3 ;
        RECT 2361.3400 1309.9400 2362.9400 1310.4200 ;
        RECT 2376.8800 1309.9400 2378.4800 1310.4200 ;
        RECT 2376.8800 1299.0600 2378.4800 1299.5400 ;
        RECT 2376.8800 1304.5000 2378.4800 1304.9800 ;
        RECT 2361.3400 1299.0600 2362.9400 1299.5400 ;
        RECT 2361.3400 1304.5000 2362.9400 1304.9800 ;
        RECT 2376.8800 1282.7400 2378.4800 1283.2200 ;
        RECT 2376.8800 1288.1800 2378.4800 1288.6600 ;
        RECT 2361.3400 1282.7400 2362.9400 1283.2200 ;
        RECT 2361.3400 1288.1800 2362.9400 1288.6600 ;
        RECT 2376.8800 1271.8600 2378.4800 1272.3400 ;
        RECT 2376.8800 1277.3000 2378.4800 1277.7800 ;
        RECT 2361.3400 1271.8600 2362.9400 1272.3400 ;
        RECT 2361.3400 1277.3000 2362.9400 1277.7800 ;
        RECT 2361.3400 1293.6200 2362.9400 1294.1000 ;
        RECT 2376.8800 1293.6200 2378.4800 1294.1000 ;
        RECT 2316.3400 1299.0600 2317.9400 1299.5400 ;
        RECT 2316.3400 1304.5000 2317.9400 1304.9800 ;
        RECT 2316.3400 1309.9400 2317.9400 1310.4200 ;
        RECT 2316.3400 1282.7400 2317.9400 1283.2200 ;
        RECT 2316.3400 1288.1800 2317.9400 1288.6600 ;
        RECT 2316.3400 1277.3000 2317.9400 1277.7800 ;
        RECT 2316.3400 1271.8600 2317.9400 1272.3400 ;
        RECT 2316.3400 1293.6200 2317.9400 1294.1000 ;
        RECT 2376.8800 1255.5400 2378.4800 1256.0200 ;
        RECT 2376.8800 1260.9800 2378.4800 1261.4600 ;
        RECT 2361.3400 1255.5400 2362.9400 1256.0200 ;
        RECT 2361.3400 1260.9800 2362.9400 1261.4600 ;
        RECT 2376.8800 1239.2200 2378.4800 1239.7000 ;
        RECT 2376.8800 1244.6600 2378.4800 1245.1400 ;
        RECT 2376.8800 1250.1000 2378.4800 1250.5800 ;
        RECT 2361.3400 1239.2200 2362.9400 1239.7000 ;
        RECT 2361.3400 1244.6600 2362.9400 1245.1400 ;
        RECT 2361.3400 1250.1000 2362.9400 1250.5800 ;
        RECT 2376.8800 1228.3400 2378.4800 1228.8200 ;
        RECT 2376.8800 1233.7800 2378.4800 1234.2600 ;
        RECT 2361.3400 1228.3400 2362.9400 1228.8200 ;
        RECT 2361.3400 1233.7800 2362.9400 1234.2600 ;
        RECT 2376.8800 1212.0200 2378.4800 1212.5000 ;
        RECT 2376.8800 1217.4600 2378.4800 1217.9400 ;
        RECT 2376.8800 1222.9000 2378.4800 1223.3800 ;
        RECT 2361.3400 1212.0200 2362.9400 1212.5000 ;
        RECT 2361.3400 1217.4600 2362.9400 1217.9400 ;
        RECT 2361.3400 1222.9000 2362.9400 1223.3800 ;
        RECT 2316.3400 1255.5400 2317.9400 1256.0200 ;
        RECT 2316.3400 1260.9800 2317.9400 1261.4600 ;
        RECT 2316.3400 1239.2200 2317.9400 1239.7000 ;
        RECT 2316.3400 1244.6600 2317.9400 1245.1400 ;
        RECT 2316.3400 1250.1000 2317.9400 1250.5800 ;
        RECT 2316.3400 1228.3400 2317.9400 1228.8200 ;
        RECT 2316.3400 1233.7800 2317.9400 1234.2600 ;
        RECT 2316.3400 1212.0200 2317.9400 1212.5000 ;
        RECT 2316.3400 1217.4600 2317.9400 1217.9400 ;
        RECT 2316.3400 1222.9000 2317.9400 1223.3800 ;
        RECT 2316.3400 1266.4200 2317.9400 1266.9000 ;
        RECT 2361.3400 1266.4200 2362.9400 1266.9000 ;
        RECT 2376.8800 1266.4200 2378.4800 1266.9000 ;
        RECT 2271.3400 1299.0600 2272.9400 1299.5400 ;
        RECT 2271.3400 1304.5000 2272.9400 1304.9800 ;
        RECT 2271.3400 1309.9400 2272.9400 1310.4200 ;
        RECT 2226.3400 1299.0600 2227.9400 1299.5400 ;
        RECT 2226.3400 1304.5000 2227.9400 1304.9800 ;
        RECT 2226.3400 1309.9400 2227.9400 1310.4200 ;
        RECT 2271.3400 1282.7400 2272.9400 1283.2200 ;
        RECT 2271.3400 1288.1800 2272.9400 1288.6600 ;
        RECT 2271.3400 1271.8600 2272.9400 1272.3400 ;
        RECT 2271.3400 1277.3000 2272.9400 1277.7800 ;
        RECT 2226.3400 1282.7400 2227.9400 1283.2200 ;
        RECT 2226.3400 1288.1800 2227.9400 1288.6600 ;
        RECT 2226.3400 1271.8600 2227.9400 1272.3400 ;
        RECT 2226.3400 1277.3000 2227.9400 1277.7800 ;
        RECT 2226.3400 1293.6200 2227.9400 1294.1000 ;
        RECT 2271.3400 1293.6200 2272.9400 1294.1000 ;
        RECT 2174.1800 1309.9400 2175.7800 1310.4200 ;
        RECT 2181.3400 1309.9400 2182.9400 1310.4200 ;
        RECT 2181.3400 1299.0600 2182.9400 1299.5400 ;
        RECT 2181.3400 1304.5000 2182.9400 1304.9800 ;
        RECT 2174.1800 1299.0600 2175.7800 1299.5400 ;
        RECT 2174.1800 1304.5000 2175.7800 1304.9800 ;
        RECT 2181.3400 1282.7400 2182.9400 1283.2200 ;
        RECT 2181.3400 1288.1800 2182.9400 1288.6600 ;
        RECT 2174.1800 1282.7400 2175.7800 1283.2200 ;
        RECT 2174.1800 1288.1800 2175.7800 1288.6600 ;
        RECT 2181.3400 1271.8600 2182.9400 1272.3400 ;
        RECT 2181.3400 1277.3000 2182.9400 1277.7800 ;
        RECT 2174.1800 1271.8600 2175.7800 1272.3400 ;
        RECT 2174.1800 1277.3000 2175.7800 1277.7800 ;
        RECT 2174.1800 1293.6200 2175.7800 1294.1000 ;
        RECT 2181.3400 1293.6200 2182.9400 1294.1000 ;
        RECT 2271.3400 1255.5400 2272.9400 1256.0200 ;
        RECT 2271.3400 1260.9800 2272.9400 1261.4600 ;
        RECT 2271.3400 1239.2200 2272.9400 1239.7000 ;
        RECT 2271.3400 1244.6600 2272.9400 1245.1400 ;
        RECT 2271.3400 1250.1000 2272.9400 1250.5800 ;
        RECT 2226.3400 1255.5400 2227.9400 1256.0200 ;
        RECT 2226.3400 1260.9800 2227.9400 1261.4600 ;
        RECT 2226.3400 1239.2200 2227.9400 1239.7000 ;
        RECT 2226.3400 1244.6600 2227.9400 1245.1400 ;
        RECT 2226.3400 1250.1000 2227.9400 1250.5800 ;
        RECT 2271.3400 1228.3400 2272.9400 1228.8200 ;
        RECT 2271.3400 1233.7800 2272.9400 1234.2600 ;
        RECT 2271.3400 1212.0200 2272.9400 1212.5000 ;
        RECT 2271.3400 1217.4600 2272.9400 1217.9400 ;
        RECT 2271.3400 1222.9000 2272.9400 1223.3800 ;
        RECT 2226.3400 1228.3400 2227.9400 1228.8200 ;
        RECT 2226.3400 1233.7800 2227.9400 1234.2600 ;
        RECT 2226.3400 1212.0200 2227.9400 1212.5000 ;
        RECT 2226.3400 1217.4600 2227.9400 1217.9400 ;
        RECT 2226.3400 1222.9000 2227.9400 1223.3800 ;
        RECT 2181.3400 1255.5400 2182.9400 1256.0200 ;
        RECT 2181.3400 1260.9800 2182.9400 1261.4600 ;
        RECT 2174.1800 1255.5400 2175.7800 1256.0200 ;
        RECT 2174.1800 1260.9800 2175.7800 1261.4600 ;
        RECT 2181.3400 1239.2200 2182.9400 1239.7000 ;
        RECT 2181.3400 1244.6600 2182.9400 1245.1400 ;
        RECT 2181.3400 1250.1000 2182.9400 1250.5800 ;
        RECT 2174.1800 1239.2200 2175.7800 1239.7000 ;
        RECT 2174.1800 1244.6600 2175.7800 1245.1400 ;
        RECT 2174.1800 1250.1000 2175.7800 1250.5800 ;
        RECT 2181.3400 1228.3400 2182.9400 1228.8200 ;
        RECT 2181.3400 1233.7800 2182.9400 1234.2600 ;
        RECT 2174.1800 1228.3400 2175.7800 1228.8200 ;
        RECT 2174.1800 1233.7800 2175.7800 1234.2600 ;
        RECT 2181.3400 1212.0200 2182.9400 1212.5000 ;
        RECT 2181.3400 1217.4600 2182.9400 1217.9400 ;
        RECT 2181.3400 1222.9000 2182.9400 1223.3800 ;
        RECT 2174.1800 1212.0200 2175.7800 1212.5000 ;
        RECT 2174.1800 1217.4600 2175.7800 1217.9400 ;
        RECT 2174.1800 1222.9000 2175.7800 1223.3800 ;
        RECT 2174.1800 1266.4200 2175.7800 1266.9000 ;
        RECT 2181.3400 1266.4200 2182.9400 1266.9000 ;
        RECT 2226.3400 1266.4200 2227.9400 1266.9000 ;
        RECT 2271.3400 1266.4200 2272.9400 1266.9000 ;
        RECT 2376.8800 1201.1400 2378.4800 1201.6200 ;
        RECT 2376.8800 1206.5800 2378.4800 1207.0600 ;
        RECT 2361.3400 1201.1400 2362.9400 1201.6200 ;
        RECT 2361.3400 1206.5800 2362.9400 1207.0600 ;
        RECT 2376.8800 1184.8200 2378.4800 1185.3000 ;
        RECT 2376.8800 1190.2600 2378.4800 1190.7400 ;
        RECT 2376.8800 1195.7000 2378.4800 1196.1800 ;
        RECT 2361.3400 1184.8200 2362.9400 1185.3000 ;
        RECT 2361.3400 1190.2600 2362.9400 1190.7400 ;
        RECT 2361.3400 1195.7000 2362.9400 1196.1800 ;
        RECT 2376.8800 1173.9400 2378.4800 1174.4200 ;
        RECT 2376.8800 1179.3800 2378.4800 1179.8600 ;
        RECT 2361.3400 1173.9400 2362.9400 1174.4200 ;
        RECT 2361.3400 1179.3800 2362.9400 1179.8600 ;
        RECT 2376.8800 1157.6200 2378.4800 1158.1000 ;
        RECT 2376.8800 1163.0600 2378.4800 1163.5400 ;
        RECT 2376.8800 1168.5000 2378.4800 1168.9800 ;
        RECT 2361.3400 1157.6200 2362.9400 1158.1000 ;
        RECT 2361.3400 1163.0600 2362.9400 1163.5400 ;
        RECT 2361.3400 1168.5000 2362.9400 1168.9800 ;
        RECT 2316.3400 1201.1400 2317.9400 1201.6200 ;
        RECT 2316.3400 1206.5800 2317.9400 1207.0600 ;
        RECT 2316.3400 1184.8200 2317.9400 1185.3000 ;
        RECT 2316.3400 1190.2600 2317.9400 1190.7400 ;
        RECT 2316.3400 1195.7000 2317.9400 1196.1800 ;
        RECT 2316.3400 1173.9400 2317.9400 1174.4200 ;
        RECT 2316.3400 1179.3800 2317.9400 1179.8600 ;
        RECT 2316.3400 1157.6200 2317.9400 1158.1000 ;
        RECT 2316.3400 1163.0600 2317.9400 1163.5400 ;
        RECT 2316.3400 1168.5000 2317.9400 1168.9800 ;
        RECT 2376.8800 1146.7400 2378.4800 1147.2200 ;
        RECT 2376.8800 1152.1800 2378.4800 1152.6600 ;
        RECT 2361.3400 1146.7400 2362.9400 1147.2200 ;
        RECT 2361.3400 1152.1800 2362.9400 1152.6600 ;
        RECT 2376.8800 1130.4200 2378.4800 1130.9000 ;
        RECT 2376.8800 1135.8600 2378.4800 1136.3400 ;
        RECT 2376.8800 1141.3000 2378.4800 1141.7800 ;
        RECT 2361.3400 1130.4200 2362.9400 1130.9000 ;
        RECT 2361.3400 1135.8600 2362.9400 1136.3400 ;
        RECT 2361.3400 1141.3000 2362.9400 1141.7800 ;
        RECT 2376.8800 1119.5400 2378.4800 1120.0200 ;
        RECT 2376.8800 1124.9800 2378.4800 1125.4600 ;
        RECT 2361.3400 1119.5400 2362.9400 1120.0200 ;
        RECT 2361.3400 1124.9800 2362.9400 1125.4600 ;
        RECT 2361.3400 1114.1000 2362.9400 1114.5800 ;
        RECT 2376.8800 1114.1000 2378.4800 1114.5800 ;
        RECT 2316.3400 1146.7400 2317.9400 1147.2200 ;
        RECT 2316.3400 1152.1800 2317.9400 1152.6600 ;
        RECT 2316.3400 1130.4200 2317.9400 1130.9000 ;
        RECT 2316.3400 1135.8600 2317.9400 1136.3400 ;
        RECT 2316.3400 1141.3000 2317.9400 1141.7800 ;
        RECT 2316.3400 1119.5400 2317.9400 1120.0200 ;
        RECT 2316.3400 1124.9800 2317.9400 1125.4600 ;
        RECT 2316.3400 1114.1000 2317.9400 1114.5800 ;
        RECT 2271.3400 1201.1400 2272.9400 1201.6200 ;
        RECT 2271.3400 1206.5800 2272.9400 1207.0600 ;
        RECT 2271.3400 1184.8200 2272.9400 1185.3000 ;
        RECT 2271.3400 1190.2600 2272.9400 1190.7400 ;
        RECT 2271.3400 1195.7000 2272.9400 1196.1800 ;
        RECT 2226.3400 1201.1400 2227.9400 1201.6200 ;
        RECT 2226.3400 1206.5800 2227.9400 1207.0600 ;
        RECT 2226.3400 1184.8200 2227.9400 1185.3000 ;
        RECT 2226.3400 1190.2600 2227.9400 1190.7400 ;
        RECT 2226.3400 1195.7000 2227.9400 1196.1800 ;
        RECT 2271.3400 1173.9400 2272.9400 1174.4200 ;
        RECT 2271.3400 1179.3800 2272.9400 1179.8600 ;
        RECT 2271.3400 1157.6200 2272.9400 1158.1000 ;
        RECT 2271.3400 1163.0600 2272.9400 1163.5400 ;
        RECT 2271.3400 1168.5000 2272.9400 1168.9800 ;
        RECT 2226.3400 1173.9400 2227.9400 1174.4200 ;
        RECT 2226.3400 1179.3800 2227.9400 1179.8600 ;
        RECT 2226.3400 1157.6200 2227.9400 1158.1000 ;
        RECT 2226.3400 1163.0600 2227.9400 1163.5400 ;
        RECT 2226.3400 1168.5000 2227.9400 1168.9800 ;
        RECT 2181.3400 1201.1400 2182.9400 1201.6200 ;
        RECT 2181.3400 1206.5800 2182.9400 1207.0600 ;
        RECT 2174.1800 1201.1400 2175.7800 1201.6200 ;
        RECT 2174.1800 1206.5800 2175.7800 1207.0600 ;
        RECT 2181.3400 1184.8200 2182.9400 1185.3000 ;
        RECT 2181.3400 1190.2600 2182.9400 1190.7400 ;
        RECT 2181.3400 1195.7000 2182.9400 1196.1800 ;
        RECT 2174.1800 1184.8200 2175.7800 1185.3000 ;
        RECT 2174.1800 1190.2600 2175.7800 1190.7400 ;
        RECT 2174.1800 1195.7000 2175.7800 1196.1800 ;
        RECT 2181.3400 1173.9400 2182.9400 1174.4200 ;
        RECT 2181.3400 1179.3800 2182.9400 1179.8600 ;
        RECT 2174.1800 1173.9400 2175.7800 1174.4200 ;
        RECT 2174.1800 1179.3800 2175.7800 1179.8600 ;
        RECT 2181.3400 1157.6200 2182.9400 1158.1000 ;
        RECT 2181.3400 1163.0600 2182.9400 1163.5400 ;
        RECT 2181.3400 1168.5000 2182.9400 1168.9800 ;
        RECT 2174.1800 1157.6200 2175.7800 1158.1000 ;
        RECT 2174.1800 1163.0600 2175.7800 1163.5400 ;
        RECT 2174.1800 1168.5000 2175.7800 1168.9800 ;
        RECT 2271.3400 1146.7400 2272.9400 1147.2200 ;
        RECT 2271.3400 1152.1800 2272.9400 1152.6600 ;
        RECT 2271.3400 1130.4200 2272.9400 1130.9000 ;
        RECT 2271.3400 1135.8600 2272.9400 1136.3400 ;
        RECT 2271.3400 1141.3000 2272.9400 1141.7800 ;
        RECT 2226.3400 1146.7400 2227.9400 1147.2200 ;
        RECT 2226.3400 1152.1800 2227.9400 1152.6600 ;
        RECT 2226.3400 1130.4200 2227.9400 1130.9000 ;
        RECT 2226.3400 1135.8600 2227.9400 1136.3400 ;
        RECT 2226.3400 1141.3000 2227.9400 1141.7800 ;
        RECT 2271.3400 1124.9800 2272.9400 1125.4600 ;
        RECT 2271.3400 1119.5400 2272.9400 1120.0200 ;
        RECT 2271.3400 1114.1000 2272.9400 1114.5800 ;
        RECT 2226.3400 1124.9800 2227.9400 1125.4600 ;
        RECT 2226.3400 1119.5400 2227.9400 1120.0200 ;
        RECT 2226.3400 1114.1000 2227.9400 1114.5800 ;
        RECT 2181.3400 1146.7400 2182.9400 1147.2200 ;
        RECT 2181.3400 1152.1800 2182.9400 1152.6600 ;
        RECT 2174.1800 1146.7400 2175.7800 1147.2200 ;
        RECT 2174.1800 1152.1800 2175.7800 1152.6600 ;
        RECT 2181.3400 1130.4200 2182.9400 1130.9000 ;
        RECT 2181.3400 1135.8600 2182.9400 1136.3400 ;
        RECT 2181.3400 1141.3000 2182.9400 1141.7800 ;
        RECT 2174.1800 1130.4200 2175.7800 1130.9000 ;
        RECT 2174.1800 1135.8600 2175.7800 1136.3400 ;
        RECT 2174.1800 1141.3000 2175.7800 1141.7800 ;
        RECT 2181.3400 1119.5400 2182.9400 1120.0200 ;
        RECT 2181.3400 1124.9800 2182.9400 1125.4600 ;
        RECT 2174.1800 1119.5400 2175.7800 1120.0200 ;
        RECT 2174.1800 1124.9800 2175.7800 1125.4600 ;
        RECT 2174.1800 1114.1000 2175.7800 1114.5800 ;
        RECT 2181.3400 1114.1000 2182.9400 1114.5800 ;
        RECT 2171.2200 1316.2900 2381.4400 1317.8900 ;
        RECT 2171.2200 1104.5900 2381.4400 1106.1900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1101.7600 2175.7800 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1319.8000 2175.7800 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1101.7600 2378.4800 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1319.8000 2378.4800 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1104.5900 2172.8200 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1104.5900 2381.4400 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1316.2900 2172.8200 1317.8900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1316.2900 2381.4400 1317.8900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 874.9500 2362.9400 1088.2500 ;
        RECT 2316.3400 874.9500 2317.9400 1088.2500 ;
        RECT 2271.3400 874.9500 2272.9400 1088.2500 ;
        RECT 2226.3400 874.9500 2227.9400 1088.2500 ;
        RECT 2181.3400 874.9500 2182.9400 1088.2500 ;
        RECT 2376.8800 872.1200 2378.4800 1091.7600 ;
        RECT 2174.1800 872.1200 2175.7800 1091.7600 ;
      LAYER met3 ;
        RECT 2361.3400 1080.3000 2362.9400 1080.7800 ;
        RECT 2376.8800 1080.3000 2378.4800 1080.7800 ;
        RECT 2376.8800 1069.4200 2378.4800 1069.9000 ;
        RECT 2376.8800 1074.8600 2378.4800 1075.3400 ;
        RECT 2361.3400 1069.4200 2362.9400 1069.9000 ;
        RECT 2361.3400 1074.8600 2362.9400 1075.3400 ;
        RECT 2376.8800 1053.1000 2378.4800 1053.5800 ;
        RECT 2376.8800 1058.5400 2378.4800 1059.0200 ;
        RECT 2361.3400 1053.1000 2362.9400 1053.5800 ;
        RECT 2361.3400 1058.5400 2362.9400 1059.0200 ;
        RECT 2376.8800 1042.2200 2378.4800 1042.7000 ;
        RECT 2376.8800 1047.6600 2378.4800 1048.1400 ;
        RECT 2361.3400 1042.2200 2362.9400 1042.7000 ;
        RECT 2361.3400 1047.6600 2362.9400 1048.1400 ;
        RECT 2361.3400 1063.9800 2362.9400 1064.4600 ;
        RECT 2376.8800 1063.9800 2378.4800 1064.4600 ;
        RECT 2316.3400 1069.4200 2317.9400 1069.9000 ;
        RECT 2316.3400 1074.8600 2317.9400 1075.3400 ;
        RECT 2316.3400 1080.3000 2317.9400 1080.7800 ;
        RECT 2316.3400 1053.1000 2317.9400 1053.5800 ;
        RECT 2316.3400 1058.5400 2317.9400 1059.0200 ;
        RECT 2316.3400 1047.6600 2317.9400 1048.1400 ;
        RECT 2316.3400 1042.2200 2317.9400 1042.7000 ;
        RECT 2316.3400 1063.9800 2317.9400 1064.4600 ;
        RECT 2376.8800 1025.9000 2378.4800 1026.3800 ;
        RECT 2376.8800 1031.3400 2378.4800 1031.8200 ;
        RECT 2361.3400 1025.9000 2362.9400 1026.3800 ;
        RECT 2361.3400 1031.3400 2362.9400 1031.8200 ;
        RECT 2376.8800 1009.5800 2378.4800 1010.0600 ;
        RECT 2376.8800 1015.0200 2378.4800 1015.5000 ;
        RECT 2376.8800 1020.4600 2378.4800 1020.9400 ;
        RECT 2361.3400 1009.5800 2362.9400 1010.0600 ;
        RECT 2361.3400 1015.0200 2362.9400 1015.5000 ;
        RECT 2361.3400 1020.4600 2362.9400 1020.9400 ;
        RECT 2376.8800 998.7000 2378.4800 999.1800 ;
        RECT 2376.8800 1004.1400 2378.4800 1004.6200 ;
        RECT 2361.3400 998.7000 2362.9400 999.1800 ;
        RECT 2361.3400 1004.1400 2362.9400 1004.6200 ;
        RECT 2376.8800 982.3800 2378.4800 982.8600 ;
        RECT 2376.8800 987.8200 2378.4800 988.3000 ;
        RECT 2376.8800 993.2600 2378.4800 993.7400 ;
        RECT 2361.3400 982.3800 2362.9400 982.8600 ;
        RECT 2361.3400 987.8200 2362.9400 988.3000 ;
        RECT 2361.3400 993.2600 2362.9400 993.7400 ;
        RECT 2316.3400 1025.9000 2317.9400 1026.3800 ;
        RECT 2316.3400 1031.3400 2317.9400 1031.8200 ;
        RECT 2316.3400 1009.5800 2317.9400 1010.0600 ;
        RECT 2316.3400 1015.0200 2317.9400 1015.5000 ;
        RECT 2316.3400 1020.4600 2317.9400 1020.9400 ;
        RECT 2316.3400 998.7000 2317.9400 999.1800 ;
        RECT 2316.3400 1004.1400 2317.9400 1004.6200 ;
        RECT 2316.3400 982.3800 2317.9400 982.8600 ;
        RECT 2316.3400 987.8200 2317.9400 988.3000 ;
        RECT 2316.3400 993.2600 2317.9400 993.7400 ;
        RECT 2316.3400 1036.7800 2317.9400 1037.2600 ;
        RECT 2361.3400 1036.7800 2362.9400 1037.2600 ;
        RECT 2376.8800 1036.7800 2378.4800 1037.2600 ;
        RECT 2271.3400 1069.4200 2272.9400 1069.9000 ;
        RECT 2271.3400 1074.8600 2272.9400 1075.3400 ;
        RECT 2271.3400 1080.3000 2272.9400 1080.7800 ;
        RECT 2226.3400 1069.4200 2227.9400 1069.9000 ;
        RECT 2226.3400 1074.8600 2227.9400 1075.3400 ;
        RECT 2226.3400 1080.3000 2227.9400 1080.7800 ;
        RECT 2271.3400 1053.1000 2272.9400 1053.5800 ;
        RECT 2271.3400 1058.5400 2272.9400 1059.0200 ;
        RECT 2271.3400 1042.2200 2272.9400 1042.7000 ;
        RECT 2271.3400 1047.6600 2272.9400 1048.1400 ;
        RECT 2226.3400 1053.1000 2227.9400 1053.5800 ;
        RECT 2226.3400 1058.5400 2227.9400 1059.0200 ;
        RECT 2226.3400 1042.2200 2227.9400 1042.7000 ;
        RECT 2226.3400 1047.6600 2227.9400 1048.1400 ;
        RECT 2226.3400 1063.9800 2227.9400 1064.4600 ;
        RECT 2271.3400 1063.9800 2272.9400 1064.4600 ;
        RECT 2174.1800 1080.3000 2175.7800 1080.7800 ;
        RECT 2181.3400 1080.3000 2182.9400 1080.7800 ;
        RECT 2181.3400 1069.4200 2182.9400 1069.9000 ;
        RECT 2181.3400 1074.8600 2182.9400 1075.3400 ;
        RECT 2174.1800 1069.4200 2175.7800 1069.9000 ;
        RECT 2174.1800 1074.8600 2175.7800 1075.3400 ;
        RECT 2181.3400 1053.1000 2182.9400 1053.5800 ;
        RECT 2181.3400 1058.5400 2182.9400 1059.0200 ;
        RECT 2174.1800 1053.1000 2175.7800 1053.5800 ;
        RECT 2174.1800 1058.5400 2175.7800 1059.0200 ;
        RECT 2181.3400 1042.2200 2182.9400 1042.7000 ;
        RECT 2181.3400 1047.6600 2182.9400 1048.1400 ;
        RECT 2174.1800 1042.2200 2175.7800 1042.7000 ;
        RECT 2174.1800 1047.6600 2175.7800 1048.1400 ;
        RECT 2174.1800 1063.9800 2175.7800 1064.4600 ;
        RECT 2181.3400 1063.9800 2182.9400 1064.4600 ;
        RECT 2271.3400 1025.9000 2272.9400 1026.3800 ;
        RECT 2271.3400 1031.3400 2272.9400 1031.8200 ;
        RECT 2271.3400 1009.5800 2272.9400 1010.0600 ;
        RECT 2271.3400 1015.0200 2272.9400 1015.5000 ;
        RECT 2271.3400 1020.4600 2272.9400 1020.9400 ;
        RECT 2226.3400 1025.9000 2227.9400 1026.3800 ;
        RECT 2226.3400 1031.3400 2227.9400 1031.8200 ;
        RECT 2226.3400 1009.5800 2227.9400 1010.0600 ;
        RECT 2226.3400 1015.0200 2227.9400 1015.5000 ;
        RECT 2226.3400 1020.4600 2227.9400 1020.9400 ;
        RECT 2271.3400 998.7000 2272.9400 999.1800 ;
        RECT 2271.3400 1004.1400 2272.9400 1004.6200 ;
        RECT 2271.3400 982.3800 2272.9400 982.8600 ;
        RECT 2271.3400 987.8200 2272.9400 988.3000 ;
        RECT 2271.3400 993.2600 2272.9400 993.7400 ;
        RECT 2226.3400 998.7000 2227.9400 999.1800 ;
        RECT 2226.3400 1004.1400 2227.9400 1004.6200 ;
        RECT 2226.3400 982.3800 2227.9400 982.8600 ;
        RECT 2226.3400 987.8200 2227.9400 988.3000 ;
        RECT 2226.3400 993.2600 2227.9400 993.7400 ;
        RECT 2181.3400 1025.9000 2182.9400 1026.3800 ;
        RECT 2181.3400 1031.3400 2182.9400 1031.8200 ;
        RECT 2174.1800 1025.9000 2175.7800 1026.3800 ;
        RECT 2174.1800 1031.3400 2175.7800 1031.8200 ;
        RECT 2181.3400 1009.5800 2182.9400 1010.0600 ;
        RECT 2181.3400 1015.0200 2182.9400 1015.5000 ;
        RECT 2181.3400 1020.4600 2182.9400 1020.9400 ;
        RECT 2174.1800 1009.5800 2175.7800 1010.0600 ;
        RECT 2174.1800 1015.0200 2175.7800 1015.5000 ;
        RECT 2174.1800 1020.4600 2175.7800 1020.9400 ;
        RECT 2181.3400 998.7000 2182.9400 999.1800 ;
        RECT 2181.3400 1004.1400 2182.9400 1004.6200 ;
        RECT 2174.1800 998.7000 2175.7800 999.1800 ;
        RECT 2174.1800 1004.1400 2175.7800 1004.6200 ;
        RECT 2181.3400 982.3800 2182.9400 982.8600 ;
        RECT 2181.3400 987.8200 2182.9400 988.3000 ;
        RECT 2181.3400 993.2600 2182.9400 993.7400 ;
        RECT 2174.1800 982.3800 2175.7800 982.8600 ;
        RECT 2174.1800 987.8200 2175.7800 988.3000 ;
        RECT 2174.1800 993.2600 2175.7800 993.7400 ;
        RECT 2174.1800 1036.7800 2175.7800 1037.2600 ;
        RECT 2181.3400 1036.7800 2182.9400 1037.2600 ;
        RECT 2226.3400 1036.7800 2227.9400 1037.2600 ;
        RECT 2271.3400 1036.7800 2272.9400 1037.2600 ;
        RECT 2376.8800 971.5000 2378.4800 971.9800 ;
        RECT 2376.8800 976.9400 2378.4800 977.4200 ;
        RECT 2361.3400 971.5000 2362.9400 971.9800 ;
        RECT 2361.3400 976.9400 2362.9400 977.4200 ;
        RECT 2376.8800 955.1800 2378.4800 955.6600 ;
        RECT 2376.8800 960.6200 2378.4800 961.1000 ;
        RECT 2376.8800 966.0600 2378.4800 966.5400 ;
        RECT 2361.3400 955.1800 2362.9400 955.6600 ;
        RECT 2361.3400 960.6200 2362.9400 961.1000 ;
        RECT 2361.3400 966.0600 2362.9400 966.5400 ;
        RECT 2376.8800 944.3000 2378.4800 944.7800 ;
        RECT 2376.8800 949.7400 2378.4800 950.2200 ;
        RECT 2361.3400 944.3000 2362.9400 944.7800 ;
        RECT 2361.3400 949.7400 2362.9400 950.2200 ;
        RECT 2376.8800 927.9800 2378.4800 928.4600 ;
        RECT 2376.8800 933.4200 2378.4800 933.9000 ;
        RECT 2376.8800 938.8600 2378.4800 939.3400 ;
        RECT 2361.3400 927.9800 2362.9400 928.4600 ;
        RECT 2361.3400 933.4200 2362.9400 933.9000 ;
        RECT 2361.3400 938.8600 2362.9400 939.3400 ;
        RECT 2316.3400 971.5000 2317.9400 971.9800 ;
        RECT 2316.3400 976.9400 2317.9400 977.4200 ;
        RECT 2316.3400 955.1800 2317.9400 955.6600 ;
        RECT 2316.3400 960.6200 2317.9400 961.1000 ;
        RECT 2316.3400 966.0600 2317.9400 966.5400 ;
        RECT 2316.3400 944.3000 2317.9400 944.7800 ;
        RECT 2316.3400 949.7400 2317.9400 950.2200 ;
        RECT 2316.3400 927.9800 2317.9400 928.4600 ;
        RECT 2316.3400 933.4200 2317.9400 933.9000 ;
        RECT 2316.3400 938.8600 2317.9400 939.3400 ;
        RECT 2376.8800 917.1000 2378.4800 917.5800 ;
        RECT 2376.8800 922.5400 2378.4800 923.0200 ;
        RECT 2361.3400 917.1000 2362.9400 917.5800 ;
        RECT 2361.3400 922.5400 2362.9400 923.0200 ;
        RECT 2376.8800 900.7800 2378.4800 901.2600 ;
        RECT 2376.8800 906.2200 2378.4800 906.7000 ;
        RECT 2376.8800 911.6600 2378.4800 912.1400 ;
        RECT 2361.3400 900.7800 2362.9400 901.2600 ;
        RECT 2361.3400 906.2200 2362.9400 906.7000 ;
        RECT 2361.3400 911.6600 2362.9400 912.1400 ;
        RECT 2376.8800 889.9000 2378.4800 890.3800 ;
        RECT 2376.8800 895.3400 2378.4800 895.8200 ;
        RECT 2361.3400 889.9000 2362.9400 890.3800 ;
        RECT 2361.3400 895.3400 2362.9400 895.8200 ;
        RECT 2361.3400 884.4600 2362.9400 884.9400 ;
        RECT 2376.8800 884.4600 2378.4800 884.9400 ;
        RECT 2316.3400 917.1000 2317.9400 917.5800 ;
        RECT 2316.3400 922.5400 2317.9400 923.0200 ;
        RECT 2316.3400 900.7800 2317.9400 901.2600 ;
        RECT 2316.3400 906.2200 2317.9400 906.7000 ;
        RECT 2316.3400 911.6600 2317.9400 912.1400 ;
        RECT 2316.3400 889.9000 2317.9400 890.3800 ;
        RECT 2316.3400 895.3400 2317.9400 895.8200 ;
        RECT 2316.3400 884.4600 2317.9400 884.9400 ;
        RECT 2271.3400 971.5000 2272.9400 971.9800 ;
        RECT 2271.3400 976.9400 2272.9400 977.4200 ;
        RECT 2271.3400 955.1800 2272.9400 955.6600 ;
        RECT 2271.3400 960.6200 2272.9400 961.1000 ;
        RECT 2271.3400 966.0600 2272.9400 966.5400 ;
        RECT 2226.3400 971.5000 2227.9400 971.9800 ;
        RECT 2226.3400 976.9400 2227.9400 977.4200 ;
        RECT 2226.3400 955.1800 2227.9400 955.6600 ;
        RECT 2226.3400 960.6200 2227.9400 961.1000 ;
        RECT 2226.3400 966.0600 2227.9400 966.5400 ;
        RECT 2271.3400 944.3000 2272.9400 944.7800 ;
        RECT 2271.3400 949.7400 2272.9400 950.2200 ;
        RECT 2271.3400 927.9800 2272.9400 928.4600 ;
        RECT 2271.3400 933.4200 2272.9400 933.9000 ;
        RECT 2271.3400 938.8600 2272.9400 939.3400 ;
        RECT 2226.3400 944.3000 2227.9400 944.7800 ;
        RECT 2226.3400 949.7400 2227.9400 950.2200 ;
        RECT 2226.3400 927.9800 2227.9400 928.4600 ;
        RECT 2226.3400 933.4200 2227.9400 933.9000 ;
        RECT 2226.3400 938.8600 2227.9400 939.3400 ;
        RECT 2181.3400 971.5000 2182.9400 971.9800 ;
        RECT 2181.3400 976.9400 2182.9400 977.4200 ;
        RECT 2174.1800 971.5000 2175.7800 971.9800 ;
        RECT 2174.1800 976.9400 2175.7800 977.4200 ;
        RECT 2181.3400 955.1800 2182.9400 955.6600 ;
        RECT 2181.3400 960.6200 2182.9400 961.1000 ;
        RECT 2181.3400 966.0600 2182.9400 966.5400 ;
        RECT 2174.1800 955.1800 2175.7800 955.6600 ;
        RECT 2174.1800 960.6200 2175.7800 961.1000 ;
        RECT 2174.1800 966.0600 2175.7800 966.5400 ;
        RECT 2181.3400 944.3000 2182.9400 944.7800 ;
        RECT 2181.3400 949.7400 2182.9400 950.2200 ;
        RECT 2174.1800 944.3000 2175.7800 944.7800 ;
        RECT 2174.1800 949.7400 2175.7800 950.2200 ;
        RECT 2181.3400 927.9800 2182.9400 928.4600 ;
        RECT 2181.3400 933.4200 2182.9400 933.9000 ;
        RECT 2181.3400 938.8600 2182.9400 939.3400 ;
        RECT 2174.1800 927.9800 2175.7800 928.4600 ;
        RECT 2174.1800 933.4200 2175.7800 933.9000 ;
        RECT 2174.1800 938.8600 2175.7800 939.3400 ;
        RECT 2271.3400 917.1000 2272.9400 917.5800 ;
        RECT 2271.3400 922.5400 2272.9400 923.0200 ;
        RECT 2271.3400 900.7800 2272.9400 901.2600 ;
        RECT 2271.3400 906.2200 2272.9400 906.7000 ;
        RECT 2271.3400 911.6600 2272.9400 912.1400 ;
        RECT 2226.3400 917.1000 2227.9400 917.5800 ;
        RECT 2226.3400 922.5400 2227.9400 923.0200 ;
        RECT 2226.3400 900.7800 2227.9400 901.2600 ;
        RECT 2226.3400 906.2200 2227.9400 906.7000 ;
        RECT 2226.3400 911.6600 2227.9400 912.1400 ;
        RECT 2271.3400 895.3400 2272.9400 895.8200 ;
        RECT 2271.3400 889.9000 2272.9400 890.3800 ;
        RECT 2271.3400 884.4600 2272.9400 884.9400 ;
        RECT 2226.3400 895.3400 2227.9400 895.8200 ;
        RECT 2226.3400 889.9000 2227.9400 890.3800 ;
        RECT 2226.3400 884.4600 2227.9400 884.9400 ;
        RECT 2181.3400 917.1000 2182.9400 917.5800 ;
        RECT 2181.3400 922.5400 2182.9400 923.0200 ;
        RECT 2174.1800 917.1000 2175.7800 917.5800 ;
        RECT 2174.1800 922.5400 2175.7800 923.0200 ;
        RECT 2181.3400 900.7800 2182.9400 901.2600 ;
        RECT 2181.3400 906.2200 2182.9400 906.7000 ;
        RECT 2181.3400 911.6600 2182.9400 912.1400 ;
        RECT 2174.1800 900.7800 2175.7800 901.2600 ;
        RECT 2174.1800 906.2200 2175.7800 906.7000 ;
        RECT 2174.1800 911.6600 2175.7800 912.1400 ;
        RECT 2181.3400 889.9000 2182.9400 890.3800 ;
        RECT 2181.3400 895.3400 2182.9400 895.8200 ;
        RECT 2174.1800 889.9000 2175.7800 890.3800 ;
        RECT 2174.1800 895.3400 2175.7800 895.8200 ;
        RECT 2174.1800 884.4600 2175.7800 884.9400 ;
        RECT 2181.3400 884.4600 2182.9400 884.9400 ;
        RECT 2171.2200 1086.6500 2381.4400 1088.2500 ;
        RECT 2171.2200 874.9500 2381.4400 876.5500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 872.1200 2175.7800 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 1090.1600 2175.7800 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 872.1200 2378.4800 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 1090.1600 2378.4800 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 874.9500 2172.8200 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 874.9500 2381.4400 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1086.6500 2172.8200 1088.2500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1086.6500 2381.4400 1088.2500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 645.3100 2362.9400 858.6100 ;
        RECT 2316.3400 645.3100 2317.9400 858.6100 ;
        RECT 2271.3400 645.3100 2272.9400 858.6100 ;
        RECT 2226.3400 645.3100 2227.9400 858.6100 ;
        RECT 2181.3400 645.3100 2182.9400 858.6100 ;
        RECT 2376.8800 642.4800 2378.4800 862.1200 ;
        RECT 2174.1800 642.4800 2175.7800 862.1200 ;
      LAYER met3 ;
        RECT 2361.3400 850.6600 2362.9400 851.1400 ;
        RECT 2376.8800 850.6600 2378.4800 851.1400 ;
        RECT 2376.8800 839.7800 2378.4800 840.2600 ;
        RECT 2376.8800 845.2200 2378.4800 845.7000 ;
        RECT 2361.3400 839.7800 2362.9400 840.2600 ;
        RECT 2361.3400 845.2200 2362.9400 845.7000 ;
        RECT 2376.8800 823.4600 2378.4800 823.9400 ;
        RECT 2376.8800 828.9000 2378.4800 829.3800 ;
        RECT 2361.3400 823.4600 2362.9400 823.9400 ;
        RECT 2361.3400 828.9000 2362.9400 829.3800 ;
        RECT 2376.8800 812.5800 2378.4800 813.0600 ;
        RECT 2376.8800 818.0200 2378.4800 818.5000 ;
        RECT 2361.3400 812.5800 2362.9400 813.0600 ;
        RECT 2361.3400 818.0200 2362.9400 818.5000 ;
        RECT 2361.3400 834.3400 2362.9400 834.8200 ;
        RECT 2376.8800 834.3400 2378.4800 834.8200 ;
        RECT 2316.3400 839.7800 2317.9400 840.2600 ;
        RECT 2316.3400 845.2200 2317.9400 845.7000 ;
        RECT 2316.3400 850.6600 2317.9400 851.1400 ;
        RECT 2316.3400 823.4600 2317.9400 823.9400 ;
        RECT 2316.3400 828.9000 2317.9400 829.3800 ;
        RECT 2316.3400 818.0200 2317.9400 818.5000 ;
        RECT 2316.3400 812.5800 2317.9400 813.0600 ;
        RECT 2316.3400 834.3400 2317.9400 834.8200 ;
        RECT 2376.8800 796.2600 2378.4800 796.7400 ;
        RECT 2376.8800 801.7000 2378.4800 802.1800 ;
        RECT 2361.3400 796.2600 2362.9400 796.7400 ;
        RECT 2361.3400 801.7000 2362.9400 802.1800 ;
        RECT 2376.8800 779.9400 2378.4800 780.4200 ;
        RECT 2376.8800 785.3800 2378.4800 785.8600 ;
        RECT 2376.8800 790.8200 2378.4800 791.3000 ;
        RECT 2361.3400 779.9400 2362.9400 780.4200 ;
        RECT 2361.3400 785.3800 2362.9400 785.8600 ;
        RECT 2361.3400 790.8200 2362.9400 791.3000 ;
        RECT 2376.8800 769.0600 2378.4800 769.5400 ;
        RECT 2376.8800 774.5000 2378.4800 774.9800 ;
        RECT 2361.3400 769.0600 2362.9400 769.5400 ;
        RECT 2361.3400 774.5000 2362.9400 774.9800 ;
        RECT 2376.8800 752.7400 2378.4800 753.2200 ;
        RECT 2376.8800 758.1800 2378.4800 758.6600 ;
        RECT 2376.8800 763.6200 2378.4800 764.1000 ;
        RECT 2361.3400 752.7400 2362.9400 753.2200 ;
        RECT 2361.3400 758.1800 2362.9400 758.6600 ;
        RECT 2361.3400 763.6200 2362.9400 764.1000 ;
        RECT 2316.3400 796.2600 2317.9400 796.7400 ;
        RECT 2316.3400 801.7000 2317.9400 802.1800 ;
        RECT 2316.3400 779.9400 2317.9400 780.4200 ;
        RECT 2316.3400 785.3800 2317.9400 785.8600 ;
        RECT 2316.3400 790.8200 2317.9400 791.3000 ;
        RECT 2316.3400 769.0600 2317.9400 769.5400 ;
        RECT 2316.3400 774.5000 2317.9400 774.9800 ;
        RECT 2316.3400 752.7400 2317.9400 753.2200 ;
        RECT 2316.3400 758.1800 2317.9400 758.6600 ;
        RECT 2316.3400 763.6200 2317.9400 764.1000 ;
        RECT 2316.3400 807.1400 2317.9400 807.6200 ;
        RECT 2361.3400 807.1400 2362.9400 807.6200 ;
        RECT 2376.8800 807.1400 2378.4800 807.6200 ;
        RECT 2271.3400 839.7800 2272.9400 840.2600 ;
        RECT 2271.3400 845.2200 2272.9400 845.7000 ;
        RECT 2271.3400 850.6600 2272.9400 851.1400 ;
        RECT 2226.3400 839.7800 2227.9400 840.2600 ;
        RECT 2226.3400 845.2200 2227.9400 845.7000 ;
        RECT 2226.3400 850.6600 2227.9400 851.1400 ;
        RECT 2271.3400 823.4600 2272.9400 823.9400 ;
        RECT 2271.3400 828.9000 2272.9400 829.3800 ;
        RECT 2271.3400 812.5800 2272.9400 813.0600 ;
        RECT 2271.3400 818.0200 2272.9400 818.5000 ;
        RECT 2226.3400 823.4600 2227.9400 823.9400 ;
        RECT 2226.3400 828.9000 2227.9400 829.3800 ;
        RECT 2226.3400 812.5800 2227.9400 813.0600 ;
        RECT 2226.3400 818.0200 2227.9400 818.5000 ;
        RECT 2226.3400 834.3400 2227.9400 834.8200 ;
        RECT 2271.3400 834.3400 2272.9400 834.8200 ;
        RECT 2174.1800 850.6600 2175.7800 851.1400 ;
        RECT 2181.3400 850.6600 2182.9400 851.1400 ;
        RECT 2181.3400 839.7800 2182.9400 840.2600 ;
        RECT 2181.3400 845.2200 2182.9400 845.7000 ;
        RECT 2174.1800 839.7800 2175.7800 840.2600 ;
        RECT 2174.1800 845.2200 2175.7800 845.7000 ;
        RECT 2181.3400 823.4600 2182.9400 823.9400 ;
        RECT 2181.3400 828.9000 2182.9400 829.3800 ;
        RECT 2174.1800 823.4600 2175.7800 823.9400 ;
        RECT 2174.1800 828.9000 2175.7800 829.3800 ;
        RECT 2181.3400 812.5800 2182.9400 813.0600 ;
        RECT 2181.3400 818.0200 2182.9400 818.5000 ;
        RECT 2174.1800 812.5800 2175.7800 813.0600 ;
        RECT 2174.1800 818.0200 2175.7800 818.5000 ;
        RECT 2174.1800 834.3400 2175.7800 834.8200 ;
        RECT 2181.3400 834.3400 2182.9400 834.8200 ;
        RECT 2271.3400 796.2600 2272.9400 796.7400 ;
        RECT 2271.3400 801.7000 2272.9400 802.1800 ;
        RECT 2271.3400 779.9400 2272.9400 780.4200 ;
        RECT 2271.3400 785.3800 2272.9400 785.8600 ;
        RECT 2271.3400 790.8200 2272.9400 791.3000 ;
        RECT 2226.3400 796.2600 2227.9400 796.7400 ;
        RECT 2226.3400 801.7000 2227.9400 802.1800 ;
        RECT 2226.3400 779.9400 2227.9400 780.4200 ;
        RECT 2226.3400 785.3800 2227.9400 785.8600 ;
        RECT 2226.3400 790.8200 2227.9400 791.3000 ;
        RECT 2271.3400 769.0600 2272.9400 769.5400 ;
        RECT 2271.3400 774.5000 2272.9400 774.9800 ;
        RECT 2271.3400 752.7400 2272.9400 753.2200 ;
        RECT 2271.3400 758.1800 2272.9400 758.6600 ;
        RECT 2271.3400 763.6200 2272.9400 764.1000 ;
        RECT 2226.3400 769.0600 2227.9400 769.5400 ;
        RECT 2226.3400 774.5000 2227.9400 774.9800 ;
        RECT 2226.3400 752.7400 2227.9400 753.2200 ;
        RECT 2226.3400 758.1800 2227.9400 758.6600 ;
        RECT 2226.3400 763.6200 2227.9400 764.1000 ;
        RECT 2181.3400 796.2600 2182.9400 796.7400 ;
        RECT 2181.3400 801.7000 2182.9400 802.1800 ;
        RECT 2174.1800 796.2600 2175.7800 796.7400 ;
        RECT 2174.1800 801.7000 2175.7800 802.1800 ;
        RECT 2181.3400 779.9400 2182.9400 780.4200 ;
        RECT 2181.3400 785.3800 2182.9400 785.8600 ;
        RECT 2181.3400 790.8200 2182.9400 791.3000 ;
        RECT 2174.1800 779.9400 2175.7800 780.4200 ;
        RECT 2174.1800 785.3800 2175.7800 785.8600 ;
        RECT 2174.1800 790.8200 2175.7800 791.3000 ;
        RECT 2181.3400 769.0600 2182.9400 769.5400 ;
        RECT 2181.3400 774.5000 2182.9400 774.9800 ;
        RECT 2174.1800 769.0600 2175.7800 769.5400 ;
        RECT 2174.1800 774.5000 2175.7800 774.9800 ;
        RECT 2181.3400 752.7400 2182.9400 753.2200 ;
        RECT 2181.3400 758.1800 2182.9400 758.6600 ;
        RECT 2181.3400 763.6200 2182.9400 764.1000 ;
        RECT 2174.1800 752.7400 2175.7800 753.2200 ;
        RECT 2174.1800 758.1800 2175.7800 758.6600 ;
        RECT 2174.1800 763.6200 2175.7800 764.1000 ;
        RECT 2174.1800 807.1400 2175.7800 807.6200 ;
        RECT 2181.3400 807.1400 2182.9400 807.6200 ;
        RECT 2226.3400 807.1400 2227.9400 807.6200 ;
        RECT 2271.3400 807.1400 2272.9400 807.6200 ;
        RECT 2376.8800 741.8600 2378.4800 742.3400 ;
        RECT 2376.8800 747.3000 2378.4800 747.7800 ;
        RECT 2361.3400 741.8600 2362.9400 742.3400 ;
        RECT 2361.3400 747.3000 2362.9400 747.7800 ;
        RECT 2376.8800 725.5400 2378.4800 726.0200 ;
        RECT 2376.8800 730.9800 2378.4800 731.4600 ;
        RECT 2376.8800 736.4200 2378.4800 736.9000 ;
        RECT 2361.3400 725.5400 2362.9400 726.0200 ;
        RECT 2361.3400 730.9800 2362.9400 731.4600 ;
        RECT 2361.3400 736.4200 2362.9400 736.9000 ;
        RECT 2376.8800 714.6600 2378.4800 715.1400 ;
        RECT 2376.8800 720.1000 2378.4800 720.5800 ;
        RECT 2361.3400 714.6600 2362.9400 715.1400 ;
        RECT 2361.3400 720.1000 2362.9400 720.5800 ;
        RECT 2376.8800 698.3400 2378.4800 698.8200 ;
        RECT 2376.8800 703.7800 2378.4800 704.2600 ;
        RECT 2376.8800 709.2200 2378.4800 709.7000 ;
        RECT 2361.3400 698.3400 2362.9400 698.8200 ;
        RECT 2361.3400 703.7800 2362.9400 704.2600 ;
        RECT 2361.3400 709.2200 2362.9400 709.7000 ;
        RECT 2316.3400 741.8600 2317.9400 742.3400 ;
        RECT 2316.3400 747.3000 2317.9400 747.7800 ;
        RECT 2316.3400 725.5400 2317.9400 726.0200 ;
        RECT 2316.3400 730.9800 2317.9400 731.4600 ;
        RECT 2316.3400 736.4200 2317.9400 736.9000 ;
        RECT 2316.3400 714.6600 2317.9400 715.1400 ;
        RECT 2316.3400 720.1000 2317.9400 720.5800 ;
        RECT 2316.3400 698.3400 2317.9400 698.8200 ;
        RECT 2316.3400 703.7800 2317.9400 704.2600 ;
        RECT 2316.3400 709.2200 2317.9400 709.7000 ;
        RECT 2376.8800 687.4600 2378.4800 687.9400 ;
        RECT 2376.8800 692.9000 2378.4800 693.3800 ;
        RECT 2361.3400 687.4600 2362.9400 687.9400 ;
        RECT 2361.3400 692.9000 2362.9400 693.3800 ;
        RECT 2376.8800 671.1400 2378.4800 671.6200 ;
        RECT 2376.8800 676.5800 2378.4800 677.0600 ;
        RECT 2376.8800 682.0200 2378.4800 682.5000 ;
        RECT 2361.3400 671.1400 2362.9400 671.6200 ;
        RECT 2361.3400 676.5800 2362.9400 677.0600 ;
        RECT 2361.3400 682.0200 2362.9400 682.5000 ;
        RECT 2376.8800 660.2600 2378.4800 660.7400 ;
        RECT 2376.8800 665.7000 2378.4800 666.1800 ;
        RECT 2361.3400 660.2600 2362.9400 660.7400 ;
        RECT 2361.3400 665.7000 2362.9400 666.1800 ;
        RECT 2361.3400 654.8200 2362.9400 655.3000 ;
        RECT 2376.8800 654.8200 2378.4800 655.3000 ;
        RECT 2316.3400 687.4600 2317.9400 687.9400 ;
        RECT 2316.3400 692.9000 2317.9400 693.3800 ;
        RECT 2316.3400 671.1400 2317.9400 671.6200 ;
        RECT 2316.3400 676.5800 2317.9400 677.0600 ;
        RECT 2316.3400 682.0200 2317.9400 682.5000 ;
        RECT 2316.3400 660.2600 2317.9400 660.7400 ;
        RECT 2316.3400 665.7000 2317.9400 666.1800 ;
        RECT 2316.3400 654.8200 2317.9400 655.3000 ;
        RECT 2271.3400 741.8600 2272.9400 742.3400 ;
        RECT 2271.3400 747.3000 2272.9400 747.7800 ;
        RECT 2271.3400 725.5400 2272.9400 726.0200 ;
        RECT 2271.3400 730.9800 2272.9400 731.4600 ;
        RECT 2271.3400 736.4200 2272.9400 736.9000 ;
        RECT 2226.3400 741.8600 2227.9400 742.3400 ;
        RECT 2226.3400 747.3000 2227.9400 747.7800 ;
        RECT 2226.3400 725.5400 2227.9400 726.0200 ;
        RECT 2226.3400 730.9800 2227.9400 731.4600 ;
        RECT 2226.3400 736.4200 2227.9400 736.9000 ;
        RECT 2271.3400 714.6600 2272.9400 715.1400 ;
        RECT 2271.3400 720.1000 2272.9400 720.5800 ;
        RECT 2271.3400 698.3400 2272.9400 698.8200 ;
        RECT 2271.3400 703.7800 2272.9400 704.2600 ;
        RECT 2271.3400 709.2200 2272.9400 709.7000 ;
        RECT 2226.3400 714.6600 2227.9400 715.1400 ;
        RECT 2226.3400 720.1000 2227.9400 720.5800 ;
        RECT 2226.3400 698.3400 2227.9400 698.8200 ;
        RECT 2226.3400 703.7800 2227.9400 704.2600 ;
        RECT 2226.3400 709.2200 2227.9400 709.7000 ;
        RECT 2181.3400 741.8600 2182.9400 742.3400 ;
        RECT 2181.3400 747.3000 2182.9400 747.7800 ;
        RECT 2174.1800 741.8600 2175.7800 742.3400 ;
        RECT 2174.1800 747.3000 2175.7800 747.7800 ;
        RECT 2181.3400 725.5400 2182.9400 726.0200 ;
        RECT 2181.3400 730.9800 2182.9400 731.4600 ;
        RECT 2181.3400 736.4200 2182.9400 736.9000 ;
        RECT 2174.1800 725.5400 2175.7800 726.0200 ;
        RECT 2174.1800 730.9800 2175.7800 731.4600 ;
        RECT 2174.1800 736.4200 2175.7800 736.9000 ;
        RECT 2181.3400 714.6600 2182.9400 715.1400 ;
        RECT 2181.3400 720.1000 2182.9400 720.5800 ;
        RECT 2174.1800 714.6600 2175.7800 715.1400 ;
        RECT 2174.1800 720.1000 2175.7800 720.5800 ;
        RECT 2181.3400 698.3400 2182.9400 698.8200 ;
        RECT 2181.3400 703.7800 2182.9400 704.2600 ;
        RECT 2181.3400 709.2200 2182.9400 709.7000 ;
        RECT 2174.1800 698.3400 2175.7800 698.8200 ;
        RECT 2174.1800 703.7800 2175.7800 704.2600 ;
        RECT 2174.1800 709.2200 2175.7800 709.7000 ;
        RECT 2271.3400 687.4600 2272.9400 687.9400 ;
        RECT 2271.3400 692.9000 2272.9400 693.3800 ;
        RECT 2271.3400 671.1400 2272.9400 671.6200 ;
        RECT 2271.3400 676.5800 2272.9400 677.0600 ;
        RECT 2271.3400 682.0200 2272.9400 682.5000 ;
        RECT 2226.3400 687.4600 2227.9400 687.9400 ;
        RECT 2226.3400 692.9000 2227.9400 693.3800 ;
        RECT 2226.3400 671.1400 2227.9400 671.6200 ;
        RECT 2226.3400 676.5800 2227.9400 677.0600 ;
        RECT 2226.3400 682.0200 2227.9400 682.5000 ;
        RECT 2271.3400 665.7000 2272.9400 666.1800 ;
        RECT 2271.3400 660.2600 2272.9400 660.7400 ;
        RECT 2271.3400 654.8200 2272.9400 655.3000 ;
        RECT 2226.3400 665.7000 2227.9400 666.1800 ;
        RECT 2226.3400 660.2600 2227.9400 660.7400 ;
        RECT 2226.3400 654.8200 2227.9400 655.3000 ;
        RECT 2181.3400 687.4600 2182.9400 687.9400 ;
        RECT 2181.3400 692.9000 2182.9400 693.3800 ;
        RECT 2174.1800 687.4600 2175.7800 687.9400 ;
        RECT 2174.1800 692.9000 2175.7800 693.3800 ;
        RECT 2181.3400 671.1400 2182.9400 671.6200 ;
        RECT 2181.3400 676.5800 2182.9400 677.0600 ;
        RECT 2181.3400 682.0200 2182.9400 682.5000 ;
        RECT 2174.1800 671.1400 2175.7800 671.6200 ;
        RECT 2174.1800 676.5800 2175.7800 677.0600 ;
        RECT 2174.1800 682.0200 2175.7800 682.5000 ;
        RECT 2181.3400 660.2600 2182.9400 660.7400 ;
        RECT 2181.3400 665.7000 2182.9400 666.1800 ;
        RECT 2174.1800 660.2600 2175.7800 660.7400 ;
        RECT 2174.1800 665.7000 2175.7800 666.1800 ;
        RECT 2174.1800 654.8200 2175.7800 655.3000 ;
        RECT 2181.3400 654.8200 2182.9400 655.3000 ;
        RECT 2171.2200 857.0100 2381.4400 858.6100 ;
        RECT 2171.2200 645.3100 2381.4400 646.9100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 642.4800 2175.7800 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 860.5200 2175.7800 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 642.4800 2378.4800 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 860.5200 2378.4800 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 645.3100 2172.8200 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 645.3100 2381.4400 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 857.0100 2172.8200 858.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 857.0100 2381.4400 858.6100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2361.3400 415.6700 2362.9400 628.9700 ;
        RECT 2316.3400 415.6700 2317.9400 628.9700 ;
        RECT 2271.3400 415.6700 2272.9400 628.9700 ;
        RECT 2226.3400 415.6700 2227.9400 628.9700 ;
        RECT 2181.3400 415.6700 2182.9400 628.9700 ;
        RECT 2376.8800 412.8400 2378.4800 632.4800 ;
        RECT 2174.1800 412.8400 2175.7800 632.4800 ;
      LAYER met3 ;
        RECT 2361.3400 621.0200 2362.9400 621.5000 ;
        RECT 2376.8800 621.0200 2378.4800 621.5000 ;
        RECT 2376.8800 610.1400 2378.4800 610.6200 ;
        RECT 2376.8800 615.5800 2378.4800 616.0600 ;
        RECT 2361.3400 610.1400 2362.9400 610.6200 ;
        RECT 2361.3400 615.5800 2362.9400 616.0600 ;
        RECT 2376.8800 593.8200 2378.4800 594.3000 ;
        RECT 2376.8800 599.2600 2378.4800 599.7400 ;
        RECT 2361.3400 593.8200 2362.9400 594.3000 ;
        RECT 2361.3400 599.2600 2362.9400 599.7400 ;
        RECT 2376.8800 582.9400 2378.4800 583.4200 ;
        RECT 2376.8800 588.3800 2378.4800 588.8600 ;
        RECT 2361.3400 582.9400 2362.9400 583.4200 ;
        RECT 2361.3400 588.3800 2362.9400 588.8600 ;
        RECT 2361.3400 604.7000 2362.9400 605.1800 ;
        RECT 2376.8800 604.7000 2378.4800 605.1800 ;
        RECT 2316.3400 610.1400 2317.9400 610.6200 ;
        RECT 2316.3400 615.5800 2317.9400 616.0600 ;
        RECT 2316.3400 621.0200 2317.9400 621.5000 ;
        RECT 2316.3400 593.8200 2317.9400 594.3000 ;
        RECT 2316.3400 599.2600 2317.9400 599.7400 ;
        RECT 2316.3400 588.3800 2317.9400 588.8600 ;
        RECT 2316.3400 582.9400 2317.9400 583.4200 ;
        RECT 2316.3400 604.7000 2317.9400 605.1800 ;
        RECT 2376.8800 566.6200 2378.4800 567.1000 ;
        RECT 2376.8800 572.0600 2378.4800 572.5400 ;
        RECT 2361.3400 566.6200 2362.9400 567.1000 ;
        RECT 2361.3400 572.0600 2362.9400 572.5400 ;
        RECT 2376.8800 550.3000 2378.4800 550.7800 ;
        RECT 2376.8800 555.7400 2378.4800 556.2200 ;
        RECT 2376.8800 561.1800 2378.4800 561.6600 ;
        RECT 2361.3400 550.3000 2362.9400 550.7800 ;
        RECT 2361.3400 555.7400 2362.9400 556.2200 ;
        RECT 2361.3400 561.1800 2362.9400 561.6600 ;
        RECT 2376.8800 539.4200 2378.4800 539.9000 ;
        RECT 2376.8800 544.8600 2378.4800 545.3400 ;
        RECT 2361.3400 539.4200 2362.9400 539.9000 ;
        RECT 2361.3400 544.8600 2362.9400 545.3400 ;
        RECT 2376.8800 523.1000 2378.4800 523.5800 ;
        RECT 2376.8800 528.5400 2378.4800 529.0200 ;
        RECT 2376.8800 533.9800 2378.4800 534.4600 ;
        RECT 2361.3400 523.1000 2362.9400 523.5800 ;
        RECT 2361.3400 528.5400 2362.9400 529.0200 ;
        RECT 2361.3400 533.9800 2362.9400 534.4600 ;
        RECT 2316.3400 566.6200 2317.9400 567.1000 ;
        RECT 2316.3400 572.0600 2317.9400 572.5400 ;
        RECT 2316.3400 550.3000 2317.9400 550.7800 ;
        RECT 2316.3400 555.7400 2317.9400 556.2200 ;
        RECT 2316.3400 561.1800 2317.9400 561.6600 ;
        RECT 2316.3400 539.4200 2317.9400 539.9000 ;
        RECT 2316.3400 544.8600 2317.9400 545.3400 ;
        RECT 2316.3400 523.1000 2317.9400 523.5800 ;
        RECT 2316.3400 528.5400 2317.9400 529.0200 ;
        RECT 2316.3400 533.9800 2317.9400 534.4600 ;
        RECT 2316.3400 577.5000 2317.9400 577.9800 ;
        RECT 2361.3400 577.5000 2362.9400 577.9800 ;
        RECT 2376.8800 577.5000 2378.4800 577.9800 ;
        RECT 2271.3400 610.1400 2272.9400 610.6200 ;
        RECT 2271.3400 615.5800 2272.9400 616.0600 ;
        RECT 2271.3400 621.0200 2272.9400 621.5000 ;
        RECT 2226.3400 610.1400 2227.9400 610.6200 ;
        RECT 2226.3400 615.5800 2227.9400 616.0600 ;
        RECT 2226.3400 621.0200 2227.9400 621.5000 ;
        RECT 2271.3400 593.8200 2272.9400 594.3000 ;
        RECT 2271.3400 599.2600 2272.9400 599.7400 ;
        RECT 2271.3400 582.9400 2272.9400 583.4200 ;
        RECT 2271.3400 588.3800 2272.9400 588.8600 ;
        RECT 2226.3400 593.8200 2227.9400 594.3000 ;
        RECT 2226.3400 599.2600 2227.9400 599.7400 ;
        RECT 2226.3400 582.9400 2227.9400 583.4200 ;
        RECT 2226.3400 588.3800 2227.9400 588.8600 ;
        RECT 2226.3400 604.7000 2227.9400 605.1800 ;
        RECT 2271.3400 604.7000 2272.9400 605.1800 ;
        RECT 2174.1800 621.0200 2175.7800 621.5000 ;
        RECT 2181.3400 621.0200 2182.9400 621.5000 ;
        RECT 2181.3400 610.1400 2182.9400 610.6200 ;
        RECT 2181.3400 615.5800 2182.9400 616.0600 ;
        RECT 2174.1800 610.1400 2175.7800 610.6200 ;
        RECT 2174.1800 615.5800 2175.7800 616.0600 ;
        RECT 2181.3400 593.8200 2182.9400 594.3000 ;
        RECT 2181.3400 599.2600 2182.9400 599.7400 ;
        RECT 2174.1800 593.8200 2175.7800 594.3000 ;
        RECT 2174.1800 599.2600 2175.7800 599.7400 ;
        RECT 2181.3400 582.9400 2182.9400 583.4200 ;
        RECT 2181.3400 588.3800 2182.9400 588.8600 ;
        RECT 2174.1800 582.9400 2175.7800 583.4200 ;
        RECT 2174.1800 588.3800 2175.7800 588.8600 ;
        RECT 2174.1800 604.7000 2175.7800 605.1800 ;
        RECT 2181.3400 604.7000 2182.9400 605.1800 ;
        RECT 2271.3400 566.6200 2272.9400 567.1000 ;
        RECT 2271.3400 572.0600 2272.9400 572.5400 ;
        RECT 2271.3400 550.3000 2272.9400 550.7800 ;
        RECT 2271.3400 555.7400 2272.9400 556.2200 ;
        RECT 2271.3400 561.1800 2272.9400 561.6600 ;
        RECT 2226.3400 566.6200 2227.9400 567.1000 ;
        RECT 2226.3400 572.0600 2227.9400 572.5400 ;
        RECT 2226.3400 550.3000 2227.9400 550.7800 ;
        RECT 2226.3400 555.7400 2227.9400 556.2200 ;
        RECT 2226.3400 561.1800 2227.9400 561.6600 ;
        RECT 2271.3400 539.4200 2272.9400 539.9000 ;
        RECT 2271.3400 544.8600 2272.9400 545.3400 ;
        RECT 2271.3400 523.1000 2272.9400 523.5800 ;
        RECT 2271.3400 528.5400 2272.9400 529.0200 ;
        RECT 2271.3400 533.9800 2272.9400 534.4600 ;
        RECT 2226.3400 539.4200 2227.9400 539.9000 ;
        RECT 2226.3400 544.8600 2227.9400 545.3400 ;
        RECT 2226.3400 523.1000 2227.9400 523.5800 ;
        RECT 2226.3400 528.5400 2227.9400 529.0200 ;
        RECT 2226.3400 533.9800 2227.9400 534.4600 ;
        RECT 2181.3400 566.6200 2182.9400 567.1000 ;
        RECT 2181.3400 572.0600 2182.9400 572.5400 ;
        RECT 2174.1800 566.6200 2175.7800 567.1000 ;
        RECT 2174.1800 572.0600 2175.7800 572.5400 ;
        RECT 2181.3400 550.3000 2182.9400 550.7800 ;
        RECT 2181.3400 555.7400 2182.9400 556.2200 ;
        RECT 2181.3400 561.1800 2182.9400 561.6600 ;
        RECT 2174.1800 550.3000 2175.7800 550.7800 ;
        RECT 2174.1800 555.7400 2175.7800 556.2200 ;
        RECT 2174.1800 561.1800 2175.7800 561.6600 ;
        RECT 2181.3400 539.4200 2182.9400 539.9000 ;
        RECT 2181.3400 544.8600 2182.9400 545.3400 ;
        RECT 2174.1800 539.4200 2175.7800 539.9000 ;
        RECT 2174.1800 544.8600 2175.7800 545.3400 ;
        RECT 2181.3400 523.1000 2182.9400 523.5800 ;
        RECT 2181.3400 528.5400 2182.9400 529.0200 ;
        RECT 2181.3400 533.9800 2182.9400 534.4600 ;
        RECT 2174.1800 523.1000 2175.7800 523.5800 ;
        RECT 2174.1800 528.5400 2175.7800 529.0200 ;
        RECT 2174.1800 533.9800 2175.7800 534.4600 ;
        RECT 2174.1800 577.5000 2175.7800 577.9800 ;
        RECT 2181.3400 577.5000 2182.9400 577.9800 ;
        RECT 2226.3400 577.5000 2227.9400 577.9800 ;
        RECT 2271.3400 577.5000 2272.9400 577.9800 ;
        RECT 2376.8800 512.2200 2378.4800 512.7000 ;
        RECT 2376.8800 517.6600 2378.4800 518.1400 ;
        RECT 2361.3400 512.2200 2362.9400 512.7000 ;
        RECT 2361.3400 517.6600 2362.9400 518.1400 ;
        RECT 2376.8800 495.9000 2378.4800 496.3800 ;
        RECT 2376.8800 501.3400 2378.4800 501.8200 ;
        RECT 2376.8800 506.7800 2378.4800 507.2600 ;
        RECT 2361.3400 495.9000 2362.9400 496.3800 ;
        RECT 2361.3400 501.3400 2362.9400 501.8200 ;
        RECT 2361.3400 506.7800 2362.9400 507.2600 ;
        RECT 2376.8800 485.0200 2378.4800 485.5000 ;
        RECT 2376.8800 490.4600 2378.4800 490.9400 ;
        RECT 2361.3400 485.0200 2362.9400 485.5000 ;
        RECT 2361.3400 490.4600 2362.9400 490.9400 ;
        RECT 2376.8800 468.7000 2378.4800 469.1800 ;
        RECT 2376.8800 474.1400 2378.4800 474.6200 ;
        RECT 2376.8800 479.5800 2378.4800 480.0600 ;
        RECT 2361.3400 468.7000 2362.9400 469.1800 ;
        RECT 2361.3400 474.1400 2362.9400 474.6200 ;
        RECT 2361.3400 479.5800 2362.9400 480.0600 ;
        RECT 2316.3400 512.2200 2317.9400 512.7000 ;
        RECT 2316.3400 517.6600 2317.9400 518.1400 ;
        RECT 2316.3400 495.9000 2317.9400 496.3800 ;
        RECT 2316.3400 501.3400 2317.9400 501.8200 ;
        RECT 2316.3400 506.7800 2317.9400 507.2600 ;
        RECT 2316.3400 485.0200 2317.9400 485.5000 ;
        RECT 2316.3400 490.4600 2317.9400 490.9400 ;
        RECT 2316.3400 468.7000 2317.9400 469.1800 ;
        RECT 2316.3400 474.1400 2317.9400 474.6200 ;
        RECT 2316.3400 479.5800 2317.9400 480.0600 ;
        RECT 2376.8800 457.8200 2378.4800 458.3000 ;
        RECT 2376.8800 463.2600 2378.4800 463.7400 ;
        RECT 2361.3400 457.8200 2362.9400 458.3000 ;
        RECT 2361.3400 463.2600 2362.9400 463.7400 ;
        RECT 2376.8800 441.5000 2378.4800 441.9800 ;
        RECT 2376.8800 446.9400 2378.4800 447.4200 ;
        RECT 2376.8800 452.3800 2378.4800 452.8600 ;
        RECT 2361.3400 441.5000 2362.9400 441.9800 ;
        RECT 2361.3400 446.9400 2362.9400 447.4200 ;
        RECT 2361.3400 452.3800 2362.9400 452.8600 ;
        RECT 2376.8800 430.6200 2378.4800 431.1000 ;
        RECT 2376.8800 436.0600 2378.4800 436.5400 ;
        RECT 2361.3400 430.6200 2362.9400 431.1000 ;
        RECT 2361.3400 436.0600 2362.9400 436.5400 ;
        RECT 2361.3400 425.1800 2362.9400 425.6600 ;
        RECT 2376.8800 425.1800 2378.4800 425.6600 ;
        RECT 2316.3400 457.8200 2317.9400 458.3000 ;
        RECT 2316.3400 463.2600 2317.9400 463.7400 ;
        RECT 2316.3400 441.5000 2317.9400 441.9800 ;
        RECT 2316.3400 446.9400 2317.9400 447.4200 ;
        RECT 2316.3400 452.3800 2317.9400 452.8600 ;
        RECT 2316.3400 430.6200 2317.9400 431.1000 ;
        RECT 2316.3400 436.0600 2317.9400 436.5400 ;
        RECT 2316.3400 425.1800 2317.9400 425.6600 ;
        RECT 2271.3400 512.2200 2272.9400 512.7000 ;
        RECT 2271.3400 517.6600 2272.9400 518.1400 ;
        RECT 2271.3400 495.9000 2272.9400 496.3800 ;
        RECT 2271.3400 501.3400 2272.9400 501.8200 ;
        RECT 2271.3400 506.7800 2272.9400 507.2600 ;
        RECT 2226.3400 512.2200 2227.9400 512.7000 ;
        RECT 2226.3400 517.6600 2227.9400 518.1400 ;
        RECT 2226.3400 495.9000 2227.9400 496.3800 ;
        RECT 2226.3400 501.3400 2227.9400 501.8200 ;
        RECT 2226.3400 506.7800 2227.9400 507.2600 ;
        RECT 2271.3400 485.0200 2272.9400 485.5000 ;
        RECT 2271.3400 490.4600 2272.9400 490.9400 ;
        RECT 2271.3400 468.7000 2272.9400 469.1800 ;
        RECT 2271.3400 474.1400 2272.9400 474.6200 ;
        RECT 2271.3400 479.5800 2272.9400 480.0600 ;
        RECT 2226.3400 485.0200 2227.9400 485.5000 ;
        RECT 2226.3400 490.4600 2227.9400 490.9400 ;
        RECT 2226.3400 468.7000 2227.9400 469.1800 ;
        RECT 2226.3400 474.1400 2227.9400 474.6200 ;
        RECT 2226.3400 479.5800 2227.9400 480.0600 ;
        RECT 2181.3400 512.2200 2182.9400 512.7000 ;
        RECT 2181.3400 517.6600 2182.9400 518.1400 ;
        RECT 2174.1800 512.2200 2175.7800 512.7000 ;
        RECT 2174.1800 517.6600 2175.7800 518.1400 ;
        RECT 2181.3400 495.9000 2182.9400 496.3800 ;
        RECT 2181.3400 501.3400 2182.9400 501.8200 ;
        RECT 2181.3400 506.7800 2182.9400 507.2600 ;
        RECT 2174.1800 495.9000 2175.7800 496.3800 ;
        RECT 2174.1800 501.3400 2175.7800 501.8200 ;
        RECT 2174.1800 506.7800 2175.7800 507.2600 ;
        RECT 2181.3400 485.0200 2182.9400 485.5000 ;
        RECT 2181.3400 490.4600 2182.9400 490.9400 ;
        RECT 2174.1800 485.0200 2175.7800 485.5000 ;
        RECT 2174.1800 490.4600 2175.7800 490.9400 ;
        RECT 2181.3400 468.7000 2182.9400 469.1800 ;
        RECT 2181.3400 474.1400 2182.9400 474.6200 ;
        RECT 2181.3400 479.5800 2182.9400 480.0600 ;
        RECT 2174.1800 468.7000 2175.7800 469.1800 ;
        RECT 2174.1800 474.1400 2175.7800 474.6200 ;
        RECT 2174.1800 479.5800 2175.7800 480.0600 ;
        RECT 2271.3400 457.8200 2272.9400 458.3000 ;
        RECT 2271.3400 463.2600 2272.9400 463.7400 ;
        RECT 2271.3400 441.5000 2272.9400 441.9800 ;
        RECT 2271.3400 446.9400 2272.9400 447.4200 ;
        RECT 2271.3400 452.3800 2272.9400 452.8600 ;
        RECT 2226.3400 457.8200 2227.9400 458.3000 ;
        RECT 2226.3400 463.2600 2227.9400 463.7400 ;
        RECT 2226.3400 441.5000 2227.9400 441.9800 ;
        RECT 2226.3400 446.9400 2227.9400 447.4200 ;
        RECT 2226.3400 452.3800 2227.9400 452.8600 ;
        RECT 2271.3400 436.0600 2272.9400 436.5400 ;
        RECT 2271.3400 430.6200 2272.9400 431.1000 ;
        RECT 2271.3400 425.1800 2272.9400 425.6600 ;
        RECT 2226.3400 436.0600 2227.9400 436.5400 ;
        RECT 2226.3400 430.6200 2227.9400 431.1000 ;
        RECT 2226.3400 425.1800 2227.9400 425.6600 ;
        RECT 2181.3400 457.8200 2182.9400 458.3000 ;
        RECT 2181.3400 463.2600 2182.9400 463.7400 ;
        RECT 2174.1800 457.8200 2175.7800 458.3000 ;
        RECT 2174.1800 463.2600 2175.7800 463.7400 ;
        RECT 2181.3400 441.5000 2182.9400 441.9800 ;
        RECT 2181.3400 446.9400 2182.9400 447.4200 ;
        RECT 2181.3400 452.3800 2182.9400 452.8600 ;
        RECT 2174.1800 441.5000 2175.7800 441.9800 ;
        RECT 2174.1800 446.9400 2175.7800 447.4200 ;
        RECT 2174.1800 452.3800 2175.7800 452.8600 ;
        RECT 2181.3400 430.6200 2182.9400 431.1000 ;
        RECT 2181.3400 436.0600 2182.9400 436.5400 ;
        RECT 2174.1800 430.6200 2175.7800 431.1000 ;
        RECT 2174.1800 436.0600 2175.7800 436.5400 ;
        RECT 2174.1800 425.1800 2175.7800 425.6600 ;
        RECT 2181.3400 425.1800 2182.9400 425.6600 ;
        RECT 2171.2200 627.3700 2381.4400 628.9700 ;
        RECT 2171.2200 415.6700 2381.4400 417.2700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 412.8400 2175.7800 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2174.1800 630.8800 2175.7800 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 412.8400 2378.4800 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.8800 630.8800 2378.4800 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 415.6700 2172.8200 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 415.6700 2381.4400 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 627.3700 2172.8200 628.9700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 627.3700 2381.4400 628.9700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 183.2000 2438.6200 402.8400 ;
        RECT 2394.4000 183.2000 2396.0000 402.8400 ;
      LAYER met3 ;
        RECT 2437.0200 391.3800 2438.6200 391.8600 ;
        RECT 2437.0200 380.5000 2438.6200 380.9800 ;
        RECT 2437.0200 385.9400 2438.6200 386.4200 ;
        RECT 2437.0200 364.1800 2438.6200 364.6600 ;
        RECT 2437.0200 369.6200 2438.6200 370.1000 ;
        RECT 2437.0200 353.3000 2438.6200 353.7800 ;
        RECT 2437.0200 358.7400 2438.6200 359.2200 ;
        RECT 2437.0200 375.0600 2438.6200 375.5400 ;
        RECT 2437.0200 336.9800 2438.6200 337.4600 ;
        RECT 2437.0200 342.4200 2438.6200 342.9000 ;
        RECT 2437.0200 320.6600 2438.6200 321.1400 ;
        RECT 2437.0200 326.1000 2438.6200 326.5800 ;
        RECT 2437.0200 331.5400 2438.6200 332.0200 ;
        RECT 2437.0200 309.7800 2438.6200 310.2600 ;
        RECT 2437.0200 315.2200 2438.6200 315.7000 ;
        RECT 2437.0200 293.4600 2438.6200 293.9400 ;
        RECT 2437.0200 298.9000 2438.6200 299.3800 ;
        RECT 2437.0200 304.3400 2438.6200 304.8200 ;
        RECT 2437.0200 347.8600 2438.6200 348.3400 ;
        RECT 2394.4000 391.3800 2396.0000 391.8600 ;
        RECT 2394.4000 380.5000 2396.0000 380.9800 ;
        RECT 2394.4000 385.9400 2396.0000 386.4200 ;
        RECT 2394.4000 364.1800 2396.0000 364.6600 ;
        RECT 2394.4000 369.6200 2396.0000 370.1000 ;
        RECT 2394.4000 353.3000 2396.0000 353.7800 ;
        RECT 2394.4000 358.7400 2396.0000 359.2200 ;
        RECT 2394.4000 375.0600 2396.0000 375.5400 ;
        RECT 2394.4000 336.9800 2396.0000 337.4600 ;
        RECT 2394.4000 342.4200 2396.0000 342.9000 ;
        RECT 2394.4000 320.6600 2396.0000 321.1400 ;
        RECT 2394.4000 326.1000 2396.0000 326.5800 ;
        RECT 2394.4000 331.5400 2396.0000 332.0200 ;
        RECT 2394.4000 309.7800 2396.0000 310.2600 ;
        RECT 2394.4000 315.2200 2396.0000 315.7000 ;
        RECT 2394.4000 293.4600 2396.0000 293.9400 ;
        RECT 2394.4000 298.9000 2396.0000 299.3800 ;
        RECT 2394.4000 304.3400 2396.0000 304.8200 ;
        RECT 2394.4000 347.8600 2396.0000 348.3400 ;
        RECT 2437.0200 282.5800 2438.6200 283.0600 ;
        RECT 2437.0200 288.0200 2438.6200 288.5000 ;
        RECT 2437.0200 266.2600 2438.6200 266.7400 ;
        RECT 2437.0200 271.7000 2438.6200 272.1800 ;
        RECT 2437.0200 277.1400 2438.6200 277.6200 ;
        RECT 2437.0200 255.3800 2438.6200 255.8600 ;
        RECT 2437.0200 260.8200 2438.6200 261.3000 ;
        RECT 2437.0200 239.0600 2438.6200 239.5400 ;
        RECT 2437.0200 244.5000 2438.6200 244.9800 ;
        RECT 2437.0200 249.9400 2438.6200 250.4200 ;
        RECT 2437.0200 228.1800 2438.6200 228.6600 ;
        RECT 2437.0200 233.6200 2438.6200 234.1000 ;
        RECT 2437.0200 211.8600 2438.6200 212.3400 ;
        RECT 2437.0200 217.3000 2438.6200 217.7800 ;
        RECT 2437.0200 222.7400 2438.6200 223.2200 ;
        RECT 2437.0200 200.9800 2438.6200 201.4600 ;
        RECT 2437.0200 206.4200 2438.6200 206.9000 ;
        RECT 2437.0200 195.5400 2438.6200 196.0200 ;
        RECT 2394.4000 282.5800 2396.0000 283.0600 ;
        RECT 2394.4000 288.0200 2396.0000 288.5000 ;
        RECT 2394.4000 266.2600 2396.0000 266.7400 ;
        RECT 2394.4000 271.7000 2396.0000 272.1800 ;
        RECT 2394.4000 277.1400 2396.0000 277.6200 ;
        RECT 2394.4000 255.3800 2396.0000 255.8600 ;
        RECT 2394.4000 260.8200 2396.0000 261.3000 ;
        RECT 2394.4000 239.0600 2396.0000 239.5400 ;
        RECT 2394.4000 244.5000 2396.0000 244.9800 ;
        RECT 2394.4000 249.9400 2396.0000 250.4200 ;
        RECT 2394.4000 228.1800 2396.0000 228.6600 ;
        RECT 2394.4000 233.6200 2396.0000 234.1000 ;
        RECT 2394.4000 211.8600 2396.0000 212.3400 ;
        RECT 2394.4000 217.3000 2396.0000 217.7800 ;
        RECT 2394.4000 222.7400 2396.0000 223.2200 ;
        RECT 2394.4000 200.9800 2396.0000 201.4600 ;
        RECT 2394.4000 206.4200 2396.0000 206.9000 ;
        RECT 2394.4000 195.5400 2396.0000 196.0200 ;
        RECT 2391.4400 397.7300 2441.5800 399.3300 ;
        RECT 2391.4400 186.0300 2441.5800 187.6300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 183.2000 2396.0000 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 401.2400 2396.0000 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 183.2000 2438.6200 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 401.2400 2438.6200 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 186.0300 2393.0400 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 186.0300 2441.5800 187.6300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 397.7300 2393.0400 399.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 397.7300 2441.5800 399.3300 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 2249.9600 2438.6200 2469.6000 ;
        RECT 2394.4000 2249.9600 2396.0000 2469.6000 ;
      LAYER met3 ;
        RECT 2437.0200 2458.1400 2438.6200 2458.6200 ;
        RECT 2437.0200 2447.2600 2438.6200 2447.7400 ;
        RECT 2437.0200 2452.7000 2438.6200 2453.1800 ;
        RECT 2437.0200 2430.9400 2438.6200 2431.4200 ;
        RECT 2437.0200 2436.3800 2438.6200 2436.8600 ;
        RECT 2437.0200 2420.0600 2438.6200 2420.5400 ;
        RECT 2437.0200 2425.5000 2438.6200 2425.9800 ;
        RECT 2437.0200 2441.8200 2438.6200 2442.3000 ;
        RECT 2437.0200 2403.7400 2438.6200 2404.2200 ;
        RECT 2437.0200 2409.1800 2438.6200 2409.6600 ;
        RECT 2437.0200 2387.4200 2438.6200 2387.9000 ;
        RECT 2437.0200 2392.8600 2438.6200 2393.3400 ;
        RECT 2437.0200 2398.3000 2438.6200 2398.7800 ;
        RECT 2437.0200 2376.5400 2438.6200 2377.0200 ;
        RECT 2437.0200 2381.9800 2438.6200 2382.4600 ;
        RECT 2437.0200 2360.2200 2438.6200 2360.7000 ;
        RECT 2437.0200 2365.6600 2438.6200 2366.1400 ;
        RECT 2437.0200 2371.1000 2438.6200 2371.5800 ;
        RECT 2437.0200 2414.6200 2438.6200 2415.1000 ;
        RECT 2394.4000 2458.1400 2396.0000 2458.6200 ;
        RECT 2394.4000 2447.2600 2396.0000 2447.7400 ;
        RECT 2394.4000 2452.7000 2396.0000 2453.1800 ;
        RECT 2394.4000 2430.9400 2396.0000 2431.4200 ;
        RECT 2394.4000 2436.3800 2396.0000 2436.8600 ;
        RECT 2394.4000 2420.0600 2396.0000 2420.5400 ;
        RECT 2394.4000 2425.5000 2396.0000 2425.9800 ;
        RECT 2394.4000 2441.8200 2396.0000 2442.3000 ;
        RECT 2394.4000 2403.7400 2396.0000 2404.2200 ;
        RECT 2394.4000 2409.1800 2396.0000 2409.6600 ;
        RECT 2394.4000 2387.4200 2396.0000 2387.9000 ;
        RECT 2394.4000 2392.8600 2396.0000 2393.3400 ;
        RECT 2394.4000 2398.3000 2396.0000 2398.7800 ;
        RECT 2394.4000 2376.5400 2396.0000 2377.0200 ;
        RECT 2394.4000 2381.9800 2396.0000 2382.4600 ;
        RECT 2394.4000 2360.2200 2396.0000 2360.7000 ;
        RECT 2394.4000 2365.6600 2396.0000 2366.1400 ;
        RECT 2394.4000 2371.1000 2396.0000 2371.5800 ;
        RECT 2394.4000 2414.6200 2396.0000 2415.1000 ;
        RECT 2437.0200 2349.3400 2438.6200 2349.8200 ;
        RECT 2437.0200 2354.7800 2438.6200 2355.2600 ;
        RECT 2437.0200 2333.0200 2438.6200 2333.5000 ;
        RECT 2437.0200 2338.4600 2438.6200 2338.9400 ;
        RECT 2437.0200 2343.9000 2438.6200 2344.3800 ;
        RECT 2437.0200 2322.1400 2438.6200 2322.6200 ;
        RECT 2437.0200 2327.5800 2438.6200 2328.0600 ;
        RECT 2437.0200 2305.8200 2438.6200 2306.3000 ;
        RECT 2437.0200 2311.2600 2438.6200 2311.7400 ;
        RECT 2437.0200 2316.7000 2438.6200 2317.1800 ;
        RECT 2437.0200 2294.9400 2438.6200 2295.4200 ;
        RECT 2437.0200 2300.3800 2438.6200 2300.8600 ;
        RECT 2437.0200 2278.6200 2438.6200 2279.1000 ;
        RECT 2437.0200 2284.0600 2438.6200 2284.5400 ;
        RECT 2437.0200 2289.5000 2438.6200 2289.9800 ;
        RECT 2437.0200 2267.7400 2438.6200 2268.2200 ;
        RECT 2437.0200 2273.1800 2438.6200 2273.6600 ;
        RECT 2437.0200 2262.3000 2438.6200 2262.7800 ;
        RECT 2394.4000 2349.3400 2396.0000 2349.8200 ;
        RECT 2394.4000 2354.7800 2396.0000 2355.2600 ;
        RECT 2394.4000 2333.0200 2396.0000 2333.5000 ;
        RECT 2394.4000 2338.4600 2396.0000 2338.9400 ;
        RECT 2394.4000 2343.9000 2396.0000 2344.3800 ;
        RECT 2394.4000 2322.1400 2396.0000 2322.6200 ;
        RECT 2394.4000 2327.5800 2396.0000 2328.0600 ;
        RECT 2394.4000 2305.8200 2396.0000 2306.3000 ;
        RECT 2394.4000 2311.2600 2396.0000 2311.7400 ;
        RECT 2394.4000 2316.7000 2396.0000 2317.1800 ;
        RECT 2394.4000 2294.9400 2396.0000 2295.4200 ;
        RECT 2394.4000 2300.3800 2396.0000 2300.8600 ;
        RECT 2394.4000 2278.6200 2396.0000 2279.1000 ;
        RECT 2394.4000 2284.0600 2396.0000 2284.5400 ;
        RECT 2394.4000 2289.5000 2396.0000 2289.9800 ;
        RECT 2394.4000 2267.7400 2396.0000 2268.2200 ;
        RECT 2394.4000 2273.1800 2396.0000 2273.6600 ;
        RECT 2394.4000 2262.3000 2396.0000 2262.7800 ;
        RECT 2391.4400 2464.4900 2441.5800 2466.0900 ;
        RECT 2391.4400 2252.7900 2441.5800 2254.3900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 2249.9600 2396.0000 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 2468.0000 2396.0000 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 2249.9600 2438.6200 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 2468.0000 2438.6200 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2252.7900 2393.0400 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2252.7900 2441.5800 2254.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2464.4900 2393.0400 2466.0900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2464.4900 2441.5800 2466.0900 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 2020.3200 2438.6200 2239.9600 ;
        RECT 2394.4000 2020.3200 2396.0000 2239.9600 ;
      LAYER met3 ;
        RECT 2437.0200 2228.5000 2438.6200 2228.9800 ;
        RECT 2437.0200 2217.6200 2438.6200 2218.1000 ;
        RECT 2437.0200 2223.0600 2438.6200 2223.5400 ;
        RECT 2437.0200 2201.3000 2438.6200 2201.7800 ;
        RECT 2437.0200 2206.7400 2438.6200 2207.2200 ;
        RECT 2437.0200 2190.4200 2438.6200 2190.9000 ;
        RECT 2437.0200 2195.8600 2438.6200 2196.3400 ;
        RECT 2437.0200 2212.1800 2438.6200 2212.6600 ;
        RECT 2437.0200 2174.1000 2438.6200 2174.5800 ;
        RECT 2437.0200 2179.5400 2438.6200 2180.0200 ;
        RECT 2437.0200 2157.7800 2438.6200 2158.2600 ;
        RECT 2437.0200 2163.2200 2438.6200 2163.7000 ;
        RECT 2437.0200 2168.6600 2438.6200 2169.1400 ;
        RECT 2437.0200 2146.9000 2438.6200 2147.3800 ;
        RECT 2437.0200 2152.3400 2438.6200 2152.8200 ;
        RECT 2437.0200 2130.5800 2438.6200 2131.0600 ;
        RECT 2437.0200 2136.0200 2438.6200 2136.5000 ;
        RECT 2437.0200 2141.4600 2438.6200 2141.9400 ;
        RECT 2437.0200 2184.9800 2438.6200 2185.4600 ;
        RECT 2394.4000 2228.5000 2396.0000 2228.9800 ;
        RECT 2394.4000 2217.6200 2396.0000 2218.1000 ;
        RECT 2394.4000 2223.0600 2396.0000 2223.5400 ;
        RECT 2394.4000 2201.3000 2396.0000 2201.7800 ;
        RECT 2394.4000 2206.7400 2396.0000 2207.2200 ;
        RECT 2394.4000 2190.4200 2396.0000 2190.9000 ;
        RECT 2394.4000 2195.8600 2396.0000 2196.3400 ;
        RECT 2394.4000 2212.1800 2396.0000 2212.6600 ;
        RECT 2394.4000 2174.1000 2396.0000 2174.5800 ;
        RECT 2394.4000 2179.5400 2396.0000 2180.0200 ;
        RECT 2394.4000 2157.7800 2396.0000 2158.2600 ;
        RECT 2394.4000 2163.2200 2396.0000 2163.7000 ;
        RECT 2394.4000 2168.6600 2396.0000 2169.1400 ;
        RECT 2394.4000 2146.9000 2396.0000 2147.3800 ;
        RECT 2394.4000 2152.3400 2396.0000 2152.8200 ;
        RECT 2394.4000 2130.5800 2396.0000 2131.0600 ;
        RECT 2394.4000 2136.0200 2396.0000 2136.5000 ;
        RECT 2394.4000 2141.4600 2396.0000 2141.9400 ;
        RECT 2394.4000 2184.9800 2396.0000 2185.4600 ;
        RECT 2437.0200 2119.7000 2438.6200 2120.1800 ;
        RECT 2437.0200 2125.1400 2438.6200 2125.6200 ;
        RECT 2437.0200 2103.3800 2438.6200 2103.8600 ;
        RECT 2437.0200 2108.8200 2438.6200 2109.3000 ;
        RECT 2437.0200 2114.2600 2438.6200 2114.7400 ;
        RECT 2437.0200 2092.5000 2438.6200 2092.9800 ;
        RECT 2437.0200 2097.9400 2438.6200 2098.4200 ;
        RECT 2437.0200 2076.1800 2438.6200 2076.6600 ;
        RECT 2437.0200 2081.6200 2438.6200 2082.1000 ;
        RECT 2437.0200 2087.0600 2438.6200 2087.5400 ;
        RECT 2437.0200 2065.3000 2438.6200 2065.7800 ;
        RECT 2437.0200 2070.7400 2438.6200 2071.2200 ;
        RECT 2437.0200 2048.9800 2438.6200 2049.4600 ;
        RECT 2437.0200 2054.4200 2438.6200 2054.9000 ;
        RECT 2437.0200 2059.8600 2438.6200 2060.3400 ;
        RECT 2437.0200 2038.1000 2438.6200 2038.5800 ;
        RECT 2437.0200 2043.5400 2438.6200 2044.0200 ;
        RECT 2437.0200 2032.6600 2438.6200 2033.1400 ;
        RECT 2394.4000 2119.7000 2396.0000 2120.1800 ;
        RECT 2394.4000 2125.1400 2396.0000 2125.6200 ;
        RECT 2394.4000 2103.3800 2396.0000 2103.8600 ;
        RECT 2394.4000 2108.8200 2396.0000 2109.3000 ;
        RECT 2394.4000 2114.2600 2396.0000 2114.7400 ;
        RECT 2394.4000 2092.5000 2396.0000 2092.9800 ;
        RECT 2394.4000 2097.9400 2396.0000 2098.4200 ;
        RECT 2394.4000 2076.1800 2396.0000 2076.6600 ;
        RECT 2394.4000 2081.6200 2396.0000 2082.1000 ;
        RECT 2394.4000 2087.0600 2396.0000 2087.5400 ;
        RECT 2394.4000 2065.3000 2396.0000 2065.7800 ;
        RECT 2394.4000 2070.7400 2396.0000 2071.2200 ;
        RECT 2394.4000 2048.9800 2396.0000 2049.4600 ;
        RECT 2394.4000 2054.4200 2396.0000 2054.9000 ;
        RECT 2394.4000 2059.8600 2396.0000 2060.3400 ;
        RECT 2394.4000 2038.1000 2396.0000 2038.5800 ;
        RECT 2394.4000 2043.5400 2396.0000 2044.0200 ;
        RECT 2394.4000 2032.6600 2396.0000 2033.1400 ;
        RECT 2391.4400 2234.8500 2441.5800 2236.4500 ;
        RECT 2391.4400 2023.1500 2441.5800 2024.7500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 2020.3200 2396.0000 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 2238.3600 2396.0000 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 2020.3200 2438.6200 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 2238.3600 2438.6200 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2023.1500 2393.0400 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2023.1500 2441.5800 2024.7500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2234.8500 2393.0400 2236.4500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2234.8500 2441.5800 2236.4500 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 1790.6800 2438.6200 2010.3200 ;
        RECT 2394.4000 1790.6800 2396.0000 2010.3200 ;
      LAYER met3 ;
        RECT 2437.0200 1998.8600 2438.6200 1999.3400 ;
        RECT 2437.0200 1987.9800 2438.6200 1988.4600 ;
        RECT 2437.0200 1993.4200 2438.6200 1993.9000 ;
        RECT 2437.0200 1971.6600 2438.6200 1972.1400 ;
        RECT 2437.0200 1977.1000 2438.6200 1977.5800 ;
        RECT 2437.0200 1960.7800 2438.6200 1961.2600 ;
        RECT 2437.0200 1966.2200 2438.6200 1966.7000 ;
        RECT 2437.0200 1982.5400 2438.6200 1983.0200 ;
        RECT 2437.0200 1944.4600 2438.6200 1944.9400 ;
        RECT 2437.0200 1949.9000 2438.6200 1950.3800 ;
        RECT 2437.0200 1928.1400 2438.6200 1928.6200 ;
        RECT 2437.0200 1933.5800 2438.6200 1934.0600 ;
        RECT 2437.0200 1939.0200 2438.6200 1939.5000 ;
        RECT 2437.0200 1917.2600 2438.6200 1917.7400 ;
        RECT 2437.0200 1922.7000 2438.6200 1923.1800 ;
        RECT 2437.0200 1900.9400 2438.6200 1901.4200 ;
        RECT 2437.0200 1906.3800 2438.6200 1906.8600 ;
        RECT 2437.0200 1911.8200 2438.6200 1912.3000 ;
        RECT 2437.0200 1955.3400 2438.6200 1955.8200 ;
        RECT 2394.4000 1998.8600 2396.0000 1999.3400 ;
        RECT 2394.4000 1987.9800 2396.0000 1988.4600 ;
        RECT 2394.4000 1993.4200 2396.0000 1993.9000 ;
        RECT 2394.4000 1971.6600 2396.0000 1972.1400 ;
        RECT 2394.4000 1977.1000 2396.0000 1977.5800 ;
        RECT 2394.4000 1960.7800 2396.0000 1961.2600 ;
        RECT 2394.4000 1966.2200 2396.0000 1966.7000 ;
        RECT 2394.4000 1982.5400 2396.0000 1983.0200 ;
        RECT 2394.4000 1944.4600 2396.0000 1944.9400 ;
        RECT 2394.4000 1949.9000 2396.0000 1950.3800 ;
        RECT 2394.4000 1928.1400 2396.0000 1928.6200 ;
        RECT 2394.4000 1933.5800 2396.0000 1934.0600 ;
        RECT 2394.4000 1939.0200 2396.0000 1939.5000 ;
        RECT 2394.4000 1917.2600 2396.0000 1917.7400 ;
        RECT 2394.4000 1922.7000 2396.0000 1923.1800 ;
        RECT 2394.4000 1900.9400 2396.0000 1901.4200 ;
        RECT 2394.4000 1906.3800 2396.0000 1906.8600 ;
        RECT 2394.4000 1911.8200 2396.0000 1912.3000 ;
        RECT 2394.4000 1955.3400 2396.0000 1955.8200 ;
        RECT 2437.0200 1890.0600 2438.6200 1890.5400 ;
        RECT 2437.0200 1895.5000 2438.6200 1895.9800 ;
        RECT 2437.0200 1873.7400 2438.6200 1874.2200 ;
        RECT 2437.0200 1879.1800 2438.6200 1879.6600 ;
        RECT 2437.0200 1884.6200 2438.6200 1885.1000 ;
        RECT 2437.0200 1862.8600 2438.6200 1863.3400 ;
        RECT 2437.0200 1868.3000 2438.6200 1868.7800 ;
        RECT 2437.0200 1846.5400 2438.6200 1847.0200 ;
        RECT 2437.0200 1851.9800 2438.6200 1852.4600 ;
        RECT 2437.0200 1857.4200 2438.6200 1857.9000 ;
        RECT 2437.0200 1835.6600 2438.6200 1836.1400 ;
        RECT 2437.0200 1841.1000 2438.6200 1841.5800 ;
        RECT 2437.0200 1819.3400 2438.6200 1819.8200 ;
        RECT 2437.0200 1824.7800 2438.6200 1825.2600 ;
        RECT 2437.0200 1830.2200 2438.6200 1830.7000 ;
        RECT 2437.0200 1808.4600 2438.6200 1808.9400 ;
        RECT 2437.0200 1813.9000 2438.6200 1814.3800 ;
        RECT 2437.0200 1803.0200 2438.6200 1803.5000 ;
        RECT 2394.4000 1890.0600 2396.0000 1890.5400 ;
        RECT 2394.4000 1895.5000 2396.0000 1895.9800 ;
        RECT 2394.4000 1873.7400 2396.0000 1874.2200 ;
        RECT 2394.4000 1879.1800 2396.0000 1879.6600 ;
        RECT 2394.4000 1884.6200 2396.0000 1885.1000 ;
        RECT 2394.4000 1862.8600 2396.0000 1863.3400 ;
        RECT 2394.4000 1868.3000 2396.0000 1868.7800 ;
        RECT 2394.4000 1846.5400 2396.0000 1847.0200 ;
        RECT 2394.4000 1851.9800 2396.0000 1852.4600 ;
        RECT 2394.4000 1857.4200 2396.0000 1857.9000 ;
        RECT 2394.4000 1835.6600 2396.0000 1836.1400 ;
        RECT 2394.4000 1841.1000 2396.0000 1841.5800 ;
        RECT 2394.4000 1819.3400 2396.0000 1819.8200 ;
        RECT 2394.4000 1824.7800 2396.0000 1825.2600 ;
        RECT 2394.4000 1830.2200 2396.0000 1830.7000 ;
        RECT 2394.4000 1808.4600 2396.0000 1808.9400 ;
        RECT 2394.4000 1813.9000 2396.0000 1814.3800 ;
        RECT 2394.4000 1803.0200 2396.0000 1803.5000 ;
        RECT 2391.4400 2005.2100 2441.5800 2006.8100 ;
        RECT 2391.4400 1793.5100 2441.5800 1795.1100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1790.6800 2396.0000 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 2008.7200 2396.0000 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1790.6800 2438.6200 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 2008.7200 2438.6200 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1793.5100 2393.0400 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1793.5100 2441.5800 1795.1100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2005.2100 2393.0400 2006.8100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2005.2100 2441.5800 2006.8100 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 1561.0400 2438.6200 1780.6800 ;
        RECT 2394.4000 1561.0400 2396.0000 1780.6800 ;
      LAYER met3 ;
        RECT 2437.0200 1769.2200 2438.6200 1769.7000 ;
        RECT 2437.0200 1758.3400 2438.6200 1758.8200 ;
        RECT 2437.0200 1763.7800 2438.6200 1764.2600 ;
        RECT 2437.0200 1742.0200 2438.6200 1742.5000 ;
        RECT 2437.0200 1747.4600 2438.6200 1747.9400 ;
        RECT 2437.0200 1731.1400 2438.6200 1731.6200 ;
        RECT 2437.0200 1736.5800 2438.6200 1737.0600 ;
        RECT 2437.0200 1752.9000 2438.6200 1753.3800 ;
        RECT 2437.0200 1714.8200 2438.6200 1715.3000 ;
        RECT 2437.0200 1720.2600 2438.6200 1720.7400 ;
        RECT 2437.0200 1698.5000 2438.6200 1698.9800 ;
        RECT 2437.0200 1703.9400 2438.6200 1704.4200 ;
        RECT 2437.0200 1709.3800 2438.6200 1709.8600 ;
        RECT 2437.0200 1687.6200 2438.6200 1688.1000 ;
        RECT 2437.0200 1693.0600 2438.6200 1693.5400 ;
        RECT 2437.0200 1671.3000 2438.6200 1671.7800 ;
        RECT 2437.0200 1676.7400 2438.6200 1677.2200 ;
        RECT 2437.0200 1682.1800 2438.6200 1682.6600 ;
        RECT 2437.0200 1725.7000 2438.6200 1726.1800 ;
        RECT 2394.4000 1769.2200 2396.0000 1769.7000 ;
        RECT 2394.4000 1758.3400 2396.0000 1758.8200 ;
        RECT 2394.4000 1763.7800 2396.0000 1764.2600 ;
        RECT 2394.4000 1742.0200 2396.0000 1742.5000 ;
        RECT 2394.4000 1747.4600 2396.0000 1747.9400 ;
        RECT 2394.4000 1731.1400 2396.0000 1731.6200 ;
        RECT 2394.4000 1736.5800 2396.0000 1737.0600 ;
        RECT 2394.4000 1752.9000 2396.0000 1753.3800 ;
        RECT 2394.4000 1714.8200 2396.0000 1715.3000 ;
        RECT 2394.4000 1720.2600 2396.0000 1720.7400 ;
        RECT 2394.4000 1698.5000 2396.0000 1698.9800 ;
        RECT 2394.4000 1703.9400 2396.0000 1704.4200 ;
        RECT 2394.4000 1709.3800 2396.0000 1709.8600 ;
        RECT 2394.4000 1687.6200 2396.0000 1688.1000 ;
        RECT 2394.4000 1693.0600 2396.0000 1693.5400 ;
        RECT 2394.4000 1671.3000 2396.0000 1671.7800 ;
        RECT 2394.4000 1676.7400 2396.0000 1677.2200 ;
        RECT 2394.4000 1682.1800 2396.0000 1682.6600 ;
        RECT 2394.4000 1725.7000 2396.0000 1726.1800 ;
        RECT 2437.0200 1660.4200 2438.6200 1660.9000 ;
        RECT 2437.0200 1665.8600 2438.6200 1666.3400 ;
        RECT 2437.0200 1644.1000 2438.6200 1644.5800 ;
        RECT 2437.0200 1649.5400 2438.6200 1650.0200 ;
        RECT 2437.0200 1654.9800 2438.6200 1655.4600 ;
        RECT 2437.0200 1633.2200 2438.6200 1633.7000 ;
        RECT 2437.0200 1638.6600 2438.6200 1639.1400 ;
        RECT 2437.0200 1616.9000 2438.6200 1617.3800 ;
        RECT 2437.0200 1622.3400 2438.6200 1622.8200 ;
        RECT 2437.0200 1627.7800 2438.6200 1628.2600 ;
        RECT 2437.0200 1606.0200 2438.6200 1606.5000 ;
        RECT 2437.0200 1611.4600 2438.6200 1611.9400 ;
        RECT 2437.0200 1589.7000 2438.6200 1590.1800 ;
        RECT 2437.0200 1595.1400 2438.6200 1595.6200 ;
        RECT 2437.0200 1600.5800 2438.6200 1601.0600 ;
        RECT 2437.0200 1578.8200 2438.6200 1579.3000 ;
        RECT 2437.0200 1584.2600 2438.6200 1584.7400 ;
        RECT 2437.0200 1573.3800 2438.6200 1573.8600 ;
        RECT 2394.4000 1660.4200 2396.0000 1660.9000 ;
        RECT 2394.4000 1665.8600 2396.0000 1666.3400 ;
        RECT 2394.4000 1644.1000 2396.0000 1644.5800 ;
        RECT 2394.4000 1649.5400 2396.0000 1650.0200 ;
        RECT 2394.4000 1654.9800 2396.0000 1655.4600 ;
        RECT 2394.4000 1633.2200 2396.0000 1633.7000 ;
        RECT 2394.4000 1638.6600 2396.0000 1639.1400 ;
        RECT 2394.4000 1616.9000 2396.0000 1617.3800 ;
        RECT 2394.4000 1622.3400 2396.0000 1622.8200 ;
        RECT 2394.4000 1627.7800 2396.0000 1628.2600 ;
        RECT 2394.4000 1606.0200 2396.0000 1606.5000 ;
        RECT 2394.4000 1611.4600 2396.0000 1611.9400 ;
        RECT 2394.4000 1589.7000 2396.0000 1590.1800 ;
        RECT 2394.4000 1595.1400 2396.0000 1595.6200 ;
        RECT 2394.4000 1600.5800 2396.0000 1601.0600 ;
        RECT 2394.4000 1578.8200 2396.0000 1579.3000 ;
        RECT 2394.4000 1584.2600 2396.0000 1584.7400 ;
        RECT 2394.4000 1573.3800 2396.0000 1573.8600 ;
        RECT 2391.4400 1775.5700 2441.5800 1777.1700 ;
        RECT 2391.4400 1563.8700 2441.5800 1565.4700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1561.0400 2396.0000 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1779.0800 2396.0000 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1561.0400 2438.6200 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1779.0800 2438.6200 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1563.8700 2393.0400 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1563.8700 2441.5800 1565.4700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1775.5700 2393.0400 1777.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1775.5700 2441.5800 1777.1700 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 1331.4000 2438.6200 1551.0400 ;
        RECT 2394.4000 1331.4000 2396.0000 1551.0400 ;
      LAYER met3 ;
        RECT 2437.0200 1539.5800 2438.6200 1540.0600 ;
        RECT 2437.0200 1528.7000 2438.6200 1529.1800 ;
        RECT 2437.0200 1534.1400 2438.6200 1534.6200 ;
        RECT 2437.0200 1512.3800 2438.6200 1512.8600 ;
        RECT 2437.0200 1517.8200 2438.6200 1518.3000 ;
        RECT 2437.0200 1501.5000 2438.6200 1501.9800 ;
        RECT 2437.0200 1506.9400 2438.6200 1507.4200 ;
        RECT 2437.0200 1523.2600 2438.6200 1523.7400 ;
        RECT 2437.0200 1485.1800 2438.6200 1485.6600 ;
        RECT 2437.0200 1490.6200 2438.6200 1491.1000 ;
        RECT 2437.0200 1468.8600 2438.6200 1469.3400 ;
        RECT 2437.0200 1474.3000 2438.6200 1474.7800 ;
        RECT 2437.0200 1479.7400 2438.6200 1480.2200 ;
        RECT 2437.0200 1457.9800 2438.6200 1458.4600 ;
        RECT 2437.0200 1463.4200 2438.6200 1463.9000 ;
        RECT 2437.0200 1441.6600 2438.6200 1442.1400 ;
        RECT 2437.0200 1447.1000 2438.6200 1447.5800 ;
        RECT 2437.0200 1452.5400 2438.6200 1453.0200 ;
        RECT 2437.0200 1496.0600 2438.6200 1496.5400 ;
        RECT 2394.4000 1539.5800 2396.0000 1540.0600 ;
        RECT 2394.4000 1528.7000 2396.0000 1529.1800 ;
        RECT 2394.4000 1534.1400 2396.0000 1534.6200 ;
        RECT 2394.4000 1512.3800 2396.0000 1512.8600 ;
        RECT 2394.4000 1517.8200 2396.0000 1518.3000 ;
        RECT 2394.4000 1501.5000 2396.0000 1501.9800 ;
        RECT 2394.4000 1506.9400 2396.0000 1507.4200 ;
        RECT 2394.4000 1523.2600 2396.0000 1523.7400 ;
        RECT 2394.4000 1485.1800 2396.0000 1485.6600 ;
        RECT 2394.4000 1490.6200 2396.0000 1491.1000 ;
        RECT 2394.4000 1468.8600 2396.0000 1469.3400 ;
        RECT 2394.4000 1474.3000 2396.0000 1474.7800 ;
        RECT 2394.4000 1479.7400 2396.0000 1480.2200 ;
        RECT 2394.4000 1457.9800 2396.0000 1458.4600 ;
        RECT 2394.4000 1463.4200 2396.0000 1463.9000 ;
        RECT 2394.4000 1441.6600 2396.0000 1442.1400 ;
        RECT 2394.4000 1447.1000 2396.0000 1447.5800 ;
        RECT 2394.4000 1452.5400 2396.0000 1453.0200 ;
        RECT 2394.4000 1496.0600 2396.0000 1496.5400 ;
        RECT 2437.0200 1430.7800 2438.6200 1431.2600 ;
        RECT 2437.0200 1436.2200 2438.6200 1436.7000 ;
        RECT 2437.0200 1414.4600 2438.6200 1414.9400 ;
        RECT 2437.0200 1419.9000 2438.6200 1420.3800 ;
        RECT 2437.0200 1425.3400 2438.6200 1425.8200 ;
        RECT 2437.0200 1403.5800 2438.6200 1404.0600 ;
        RECT 2437.0200 1409.0200 2438.6200 1409.5000 ;
        RECT 2437.0200 1387.2600 2438.6200 1387.7400 ;
        RECT 2437.0200 1392.7000 2438.6200 1393.1800 ;
        RECT 2437.0200 1398.1400 2438.6200 1398.6200 ;
        RECT 2437.0200 1376.3800 2438.6200 1376.8600 ;
        RECT 2437.0200 1381.8200 2438.6200 1382.3000 ;
        RECT 2437.0200 1360.0600 2438.6200 1360.5400 ;
        RECT 2437.0200 1365.5000 2438.6200 1365.9800 ;
        RECT 2437.0200 1370.9400 2438.6200 1371.4200 ;
        RECT 2437.0200 1349.1800 2438.6200 1349.6600 ;
        RECT 2437.0200 1354.6200 2438.6200 1355.1000 ;
        RECT 2437.0200 1343.7400 2438.6200 1344.2200 ;
        RECT 2394.4000 1430.7800 2396.0000 1431.2600 ;
        RECT 2394.4000 1436.2200 2396.0000 1436.7000 ;
        RECT 2394.4000 1414.4600 2396.0000 1414.9400 ;
        RECT 2394.4000 1419.9000 2396.0000 1420.3800 ;
        RECT 2394.4000 1425.3400 2396.0000 1425.8200 ;
        RECT 2394.4000 1403.5800 2396.0000 1404.0600 ;
        RECT 2394.4000 1409.0200 2396.0000 1409.5000 ;
        RECT 2394.4000 1387.2600 2396.0000 1387.7400 ;
        RECT 2394.4000 1392.7000 2396.0000 1393.1800 ;
        RECT 2394.4000 1398.1400 2396.0000 1398.6200 ;
        RECT 2394.4000 1376.3800 2396.0000 1376.8600 ;
        RECT 2394.4000 1381.8200 2396.0000 1382.3000 ;
        RECT 2394.4000 1360.0600 2396.0000 1360.5400 ;
        RECT 2394.4000 1365.5000 2396.0000 1365.9800 ;
        RECT 2394.4000 1370.9400 2396.0000 1371.4200 ;
        RECT 2394.4000 1349.1800 2396.0000 1349.6600 ;
        RECT 2394.4000 1354.6200 2396.0000 1355.1000 ;
        RECT 2394.4000 1343.7400 2396.0000 1344.2200 ;
        RECT 2391.4400 1545.9300 2441.5800 1547.5300 ;
        RECT 2391.4400 1334.2300 2441.5800 1335.8300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1331.4000 2396.0000 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1549.4400 2396.0000 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1331.4000 2438.6200 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1549.4400 2438.6200 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1334.2300 2393.0400 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1334.2300 2441.5800 1335.8300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1545.9300 2393.0400 1547.5300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1545.9300 2441.5800 1547.5300 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 1101.7600 2438.6200 1321.4000 ;
        RECT 2394.4000 1101.7600 2396.0000 1321.4000 ;
      LAYER met3 ;
        RECT 2437.0200 1309.9400 2438.6200 1310.4200 ;
        RECT 2437.0200 1299.0600 2438.6200 1299.5400 ;
        RECT 2437.0200 1304.5000 2438.6200 1304.9800 ;
        RECT 2437.0200 1282.7400 2438.6200 1283.2200 ;
        RECT 2437.0200 1288.1800 2438.6200 1288.6600 ;
        RECT 2437.0200 1271.8600 2438.6200 1272.3400 ;
        RECT 2437.0200 1277.3000 2438.6200 1277.7800 ;
        RECT 2437.0200 1293.6200 2438.6200 1294.1000 ;
        RECT 2437.0200 1255.5400 2438.6200 1256.0200 ;
        RECT 2437.0200 1260.9800 2438.6200 1261.4600 ;
        RECT 2437.0200 1239.2200 2438.6200 1239.7000 ;
        RECT 2437.0200 1244.6600 2438.6200 1245.1400 ;
        RECT 2437.0200 1250.1000 2438.6200 1250.5800 ;
        RECT 2437.0200 1228.3400 2438.6200 1228.8200 ;
        RECT 2437.0200 1233.7800 2438.6200 1234.2600 ;
        RECT 2437.0200 1212.0200 2438.6200 1212.5000 ;
        RECT 2437.0200 1217.4600 2438.6200 1217.9400 ;
        RECT 2437.0200 1222.9000 2438.6200 1223.3800 ;
        RECT 2437.0200 1266.4200 2438.6200 1266.9000 ;
        RECT 2394.4000 1309.9400 2396.0000 1310.4200 ;
        RECT 2394.4000 1299.0600 2396.0000 1299.5400 ;
        RECT 2394.4000 1304.5000 2396.0000 1304.9800 ;
        RECT 2394.4000 1282.7400 2396.0000 1283.2200 ;
        RECT 2394.4000 1288.1800 2396.0000 1288.6600 ;
        RECT 2394.4000 1271.8600 2396.0000 1272.3400 ;
        RECT 2394.4000 1277.3000 2396.0000 1277.7800 ;
        RECT 2394.4000 1293.6200 2396.0000 1294.1000 ;
        RECT 2394.4000 1255.5400 2396.0000 1256.0200 ;
        RECT 2394.4000 1260.9800 2396.0000 1261.4600 ;
        RECT 2394.4000 1239.2200 2396.0000 1239.7000 ;
        RECT 2394.4000 1244.6600 2396.0000 1245.1400 ;
        RECT 2394.4000 1250.1000 2396.0000 1250.5800 ;
        RECT 2394.4000 1228.3400 2396.0000 1228.8200 ;
        RECT 2394.4000 1233.7800 2396.0000 1234.2600 ;
        RECT 2394.4000 1212.0200 2396.0000 1212.5000 ;
        RECT 2394.4000 1217.4600 2396.0000 1217.9400 ;
        RECT 2394.4000 1222.9000 2396.0000 1223.3800 ;
        RECT 2394.4000 1266.4200 2396.0000 1266.9000 ;
        RECT 2437.0200 1201.1400 2438.6200 1201.6200 ;
        RECT 2437.0200 1206.5800 2438.6200 1207.0600 ;
        RECT 2437.0200 1184.8200 2438.6200 1185.3000 ;
        RECT 2437.0200 1190.2600 2438.6200 1190.7400 ;
        RECT 2437.0200 1195.7000 2438.6200 1196.1800 ;
        RECT 2437.0200 1173.9400 2438.6200 1174.4200 ;
        RECT 2437.0200 1179.3800 2438.6200 1179.8600 ;
        RECT 2437.0200 1157.6200 2438.6200 1158.1000 ;
        RECT 2437.0200 1163.0600 2438.6200 1163.5400 ;
        RECT 2437.0200 1168.5000 2438.6200 1168.9800 ;
        RECT 2437.0200 1146.7400 2438.6200 1147.2200 ;
        RECT 2437.0200 1152.1800 2438.6200 1152.6600 ;
        RECT 2437.0200 1130.4200 2438.6200 1130.9000 ;
        RECT 2437.0200 1135.8600 2438.6200 1136.3400 ;
        RECT 2437.0200 1141.3000 2438.6200 1141.7800 ;
        RECT 2437.0200 1119.5400 2438.6200 1120.0200 ;
        RECT 2437.0200 1124.9800 2438.6200 1125.4600 ;
        RECT 2437.0200 1114.1000 2438.6200 1114.5800 ;
        RECT 2394.4000 1201.1400 2396.0000 1201.6200 ;
        RECT 2394.4000 1206.5800 2396.0000 1207.0600 ;
        RECT 2394.4000 1184.8200 2396.0000 1185.3000 ;
        RECT 2394.4000 1190.2600 2396.0000 1190.7400 ;
        RECT 2394.4000 1195.7000 2396.0000 1196.1800 ;
        RECT 2394.4000 1173.9400 2396.0000 1174.4200 ;
        RECT 2394.4000 1179.3800 2396.0000 1179.8600 ;
        RECT 2394.4000 1157.6200 2396.0000 1158.1000 ;
        RECT 2394.4000 1163.0600 2396.0000 1163.5400 ;
        RECT 2394.4000 1168.5000 2396.0000 1168.9800 ;
        RECT 2394.4000 1146.7400 2396.0000 1147.2200 ;
        RECT 2394.4000 1152.1800 2396.0000 1152.6600 ;
        RECT 2394.4000 1130.4200 2396.0000 1130.9000 ;
        RECT 2394.4000 1135.8600 2396.0000 1136.3400 ;
        RECT 2394.4000 1141.3000 2396.0000 1141.7800 ;
        RECT 2394.4000 1119.5400 2396.0000 1120.0200 ;
        RECT 2394.4000 1124.9800 2396.0000 1125.4600 ;
        RECT 2394.4000 1114.1000 2396.0000 1114.5800 ;
        RECT 2391.4400 1316.2900 2441.5800 1317.8900 ;
        RECT 2391.4400 1104.5900 2441.5800 1106.1900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1101.7600 2396.0000 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1319.8000 2396.0000 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1101.7600 2438.6200 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1319.8000 2438.6200 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1104.5900 2393.0400 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1104.5900 2441.5800 1106.1900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1316.2900 2393.0400 1317.8900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1316.2900 2441.5800 1317.8900 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 872.1200 2438.6200 1091.7600 ;
        RECT 2394.4000 872.1200 2396.0000 1091.7600 ;
      LAYER met3 ;
        RECT 2437.0200 1080.3000 2438.6200 1080.7800 ;
        RECT 2437.0200 1069.4200 2438.6200 1069.9000 ;
        RECT 2437.0200 1074.8600 2438.6200 1075.3400 ;
        RECT 2437.0200 1053.1000 2438.6200 1053.5800 ;
        RECT 2437.0200 1058.5400 2438.6200 1059.0200 ;
        RECT 2437.0200 1042.2200 2438.6200 1042.7000 ;
        RECT 2437.0200 1047.6600 2438.6200 1048.1400 ;
        RECT 2437.0200 1063.9800 2438.6200 1064.4600 ;
        RECT 2437.0200 1025.9000 2438.6200 1026.3800 ;
        RECT 2437.0200 1031.3400 2438.6200 1031.8200 ;
        RECT 2437.0200 1009.5800 2438.6200 1010.0600 ;
        RECT 2437.0200 1015.0200 2438.6200 1015.5000 ;
        RECT 2437.0200 1020.4600 2438.6200 1020.9400 ;
        RECT 2437.0200 998.7000 2438.6200 999.1800 ;
        RECT 2437.0200 1004.1400 2438.6200 1004.6200 ;
        RECT 2437.0200 982.3800 2438.6200 982.8600 ;
        RECT 2437.0200 987.8200 2438.6200 988.3000 ;
        RECT 2437.0200 993.2600 2438.6200 993.7400 ;
        RECT 2437.0200 1036.7800 2438.6200 1037.2600 ;
        RECT 2394.4000 1080.3000 2396.0000 1080.7800 ;
        RECT 2394.4000 1069.4200 2396.0000 1069.9000 ;
        RECT 2394.4000 1074.8600 2396.0000 1075.3400 ;
        RECT 2394.4000 1053.1000 2396.0000 1053.5800 ;
        RECT 2394.4000 1058.5400 2396.0000 1059.0200 ;
        RECT 2394.4000 1042.2200 2396.0000 1042.7000 ;
        RECT 2394.4000 1047.6600 2396.0000 1048.1400 ;
        RECT 2394.4000 1063.9800 2396.0000 1064.4600 ;
        RECT 2394.4000 1025.9000 2396.0000 1026.3800 ;
        RECT 2394.4000 1031.3400 2396.0000 1031.8200 ;
        RECT 2394.4000 1009.5800 2396.0000 1010.0600 ;
        RECT 2394.4000 1015.0200 2396.0000 1015.5000 ;
        RECT 2394.4000 1020.4600 2396.0000 1020.9400 ;
        RECT 2394.4000 998.7000 2396.0000 999.1800 ;
        RECT 2394.4000 1004.1400 2396.0000 1004.6200 ;
        RECT 2394.4000 982.3800 2396.0000 982.8600 ;
        RECT 2394.4000 987.8200 2396.0000 988.3000 ;
        RECT 2394.4000 993.2600 2396.0000 993.7400 ;
        RECT 2394.4000 1036.7800 2396.0000 1037.2600 ;
        RECT 2437.0200 971.5000 2438.6200 971.9800 ;
        RECT 2437.0200 976.9400 2438.6200 977.4200 ;
        RECT 2437.0200 955.1800 2438.6200 955.6600 ;
        RECT 2437.0200 960.6200 2438.6200 961.1000 ;
        RECT 2437.0200 966.0600 2438.6200 966.5400 ;
        RECT 2437.0200 944.3000 2438.6200 944.7800 ;
        RECT 2437.0200 949.7400 2438.6200 950.2200 ;
        RECT 2437.0200 927.9800 2438.6200 928.4600 ;
        RECT 2437.0200 933.4200 2438.6200 933.9000 ;
        RECT 2437.0200 938.8600 2438.6200 939.3400 ;
        RECT 2437.0200 917.1000 2438.6200 917.5800 ;
        RECT 2437.0200 922.5400 2438.6200 923.0200 ;
        RECT 2437.0200 900.7800 2438.6200 901.2600 ;
        RECT 2437.0200 906.2200 2438.6200 906.7000 ;
        RECT 2437.0200 911.6600 2438.6200 912.1400 ;
        RECT 2437.0200 889.9000 2438.6200 890.3800 ;
        RECT 2437.0200 895.3400 2438.6200 895.8200 ;
        RECT 2437.0200 884.4600 2438.6200 884.9400 ;
        RECT 2394.4000 971.5000 2396.0000 971.9800 ;
        RECT 2394.4000 976.9400 2396.0000 977.4200 ;
        RECT 2394.4000 955.1800 2396.0000 955.6600 ;
        RECT 2394.4000 960.6200 2396.0000 961.1000 ;
        RECT 2394.4000 966.0600 2396.0000 966.5400 ;
        RECT 2394.4000 944.3000 2396.0000 944.7800 ;
        RECT 2394.4000 949.7400 2396.0000 950.2200 ;
        RECT 2394.4000 927.9800 2396.0000 928.4600 ;
        RECT 2394.4000 933.4200 2396.0000 933.9000 ;
        RECT 2394.4000 938.8600 2396.0000 939.3400 ;
        RECT 2394.4000 917.1000 2396.0000 917.5800 ;
        RECT 2394.4000 922.5400 2396.0000 923.0200 ;
        RECT 2394.4000 900.7800 2396.0000 901.2600 ;
        RECT 2394.4000 906.2200 2396.0000 906.7000 ;
        RECT 2394.4000 911.6600 2396.0000 912.1400 ;
        RECT 2394.4000 889.9000 2396.0000 890.3800 ;
        RECT 2394.4000 895.3400 2396.0000 895.8200 ;
        RECT 2394.4000 884.4600 2396.0000 884.9400 ;
        RECT 2391.4400 1086.6500 2441.5800 1088.2500 ;
        RECT 2391.4400 874.9500 2441.5800 876.5500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 872.1200 2396.0000 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 1090.1600 2396.0000 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 872.1200 2438.6200 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 1090.1600 2438.6200 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 874.9500 2393.0400 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 874.9500 2441.5800 876.5500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1086.6500 2393.0400 1088.2500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1086.6500 2441.5800 1088.2500 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 642.4800 2438.6200 862.1200 ;
        RECT 2394.4000 642.4800 2396.0000 862.1200 ;
      LAYER met3 ;
        RECT 2437.0200 850.6600 2438.6200 851.1400 ;
        RECT 2437.0200 839.7800 2438.6200 840.2600 ;
        RECT 2437.0200 845.2200 2438.6200 845.7000 ;
        RECT 2437.0200 823.4600 2438.6200 823.9400 ;
        RECT 2437.0200 828.9000 2438.6200 829.3800 ;
        RECT 2437.0200 812.5800 2438.6200 813.0600 ;
        RECT 2437.0200 818.0200 2438.6200 818.5000 ;
        RECT 2437.0200 834.3400 2438.6200 834.8200 ;
        RECT 2437.0200 796.2600 2438.6200 796.7400 ;
        RECT 2437.0200 801.7000 2438.6200 802.1800 ;
        RECT 2437.0200 779.9400 2438.6200 780.4200 ;
        RECT 2437.0200 785.3800 2438.6200 785.8600 ;
        RECT 2437.0200 790.8200 2438.6200 791.3000 ;
        RECT 2437.0200 769.0600 2438.6200 769.5400 ;
        RECT 2437.0200 774.5000 2438.6200 774.9800 ;
        RECT 2437.0200 752.7400 2438.6200 753.2200 ;
        RECT 2437.0200 758.1800 2438.6200 758.6600 ;
        RECT 2437.0200 763.6200 2438.6200 764.1000 ;
        RECT 2437.0200 807.1400 2438.6200 807.6200 ;
        RECT 2394.4000 850.6600 2396.0000 851.1400 ;
        RECT 2394.4000 839.7800 2396.0000 840.2600 ;
        RECT 2394.4000 845.2200 2396.0000 845.7000 ;
        RECT 2394.4000 823.4600 2396.0000 823.9400 ;
        RECT 2394.4000 828.9000 2396.0000 829.3800 ;
        RECT 2394.4000 812.5800 2396.0000 813.0600 ;
        RECT 2394.4000 818.0200 2396.0000 818.5000 ;
        RECT 2394.4000 834.3400 2396.0000 834.8200 ;
        RECT 2394.4000 796.2600 2396.0000 796.7400 ;
        RECT 2394.4000 801.7000 2396.0000 802.1800 ;
        RECT 2394.4000 779.9400 2396.0000 780.4200 ;
        RECT 2394.4000 785.3800 2396.0000 785.8600 ;
        RECT 2394.4000 790.8200 2396.0000 791.3000 ;
        RECT 2394.4000 769.0600 2396.0000 769.5400 ;
        RECT 2394.4000 774.5000 2396.0000 774.9800 ;
        RECT 2394.4000 752.7400 2396.0000 753.2200 ;
        RECT 2394.4000 758.1800 2396.0000 758.6600 ;
        RECT 2394.4000 763.6200 2396.0000 764.1000 ;
        RECT 2394.4000 807.1400 2396.0000 807.6200 ;
        RECT 2437.0200 741.8600 2438.6200 742.3400 ;
        RECT 2437.0200 747.3000 2438.6200 747.7800 ;
        RECT 2437.0200 725.5400 2438.6200 726.0200 ;
        RECT 2437.0200 730.9800 2438.6200 731.4600 ;
        RECT 2437.0200 736.4200 2438.6200 736.9000 ;
        RECT 2437.0200 714.6600 2438.6200 715.1400 ;
        RECT 2437.0200 720.1000 2438.6200 720.5800 ;
        RECT 2437.0200 698.3400 2438.6200 698.8200 ;
        RECT 2437.0200 703.7800 2438.6200 704.2600 ;
        RECT 2437.0200 709.2200 2438.6200 709.7000 ;
        RECT 2437.0200 687.4600 2438.6200 687.9400 ;
        RECT 2437.0200 692.9000 2438.6200 693.3800 ;
        RECT 2437.0200 671.1400 2438.6200 671.6200 ;
        RECT 2437.0200 676.5800 2438.6200 677.0600 ;
        RECT 2437.0200 682.0200 2438.6200 682.5000 ;
        RECT 2437.0200 660.2600 2438.6200 660.7400 ;
        RECT 2437.0200 665.7000 2438.6200 666.1800 ;
        RECT 2437.0200 654.8200 2438.6200 655.3000 ;
        RECT 2394.4000 741.8600 2396.0000 742.3400 ;
        RECT 2394.4000 747.3000 2396.0000 747.7800 ;
        RECT 2394.4000 725.5400 2396.0000 726.0200 ;
        RECT 2394.4000 730.9800 2396.0000 731.4600 ;
        RECT 2394.4000 736.4200 2396.0000 736.9000 ;
        RECT 2394.4000 714.6600 2396.0000 715.1400 ;
        RECT 2394.4000 720.1000 2396.0000 720.5800 ;
        RECT 2394.4000 698.3400 2396.0000 698.8200 ;
        RECT 2394.4000 703.7800 2396.0000 704.2600 ;
        RECT 2394.4000 709.2200 2396.0000 709.7000 ;
        RECT 2394.4000 687.4600 2396.0000 687.9400 ;
        RECT 2394.4000 692.9000 2396.0000 693.3800 ;
        RECT 2394.4000 671.1400 2396.0000 671.6200 ;
        RECT 2394.4000 676.5800 2396.0000 677.0600 ;
        RECT 2394.4000 682.0200 2396.0000 682.5000 ;
        RECT 2394.4000 660.2600 2396.0000 660.7400 ;
        RECT 2394.4000 665.7000 2396.0000 666.1800 ;
        RECT 2394.4000 654.8200 2396.0000 655.3000 ;
        RECT 2391.4400 857.0100 2441.5800 858.6100 ;
        RECT 2391.4400 645.3100 2441.5800 646.9100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 642.4800 2396.0000 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 860.5200 2396.0000 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 642.4800 2438.6200 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 860.5200 2438.6200 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 645.3100 2393.0400 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 645.3100 2441.5800 646.9100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 857.0100 2393.0400 858.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 857.0100 2441.5800 858.6100 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2437.0200 412.8400 2438.6200 632.4800 ;
        RECT 2394.4000 412.8400 2396.0000 632.4800 ;
      LAYER met3 ;
        RECT 2437.0200 621.0200 2438.6200 621.5000 ;
        RECT 2437.0200 610.1400 2438.6200 610.6200 ;
        RECT 2437.0200 615.5800 2438.6200 616.0600 ;
        RECT 2437.0200 593.8200 2438.6200 594.3000 ;
        RECT 2437.0200 599.2600 2438.6200 599.7400 ;
        RECT 2437.0200 582.9400 2438.6200 583.4200 ;
        RECT 2437.0200 588.3800 2438.6200 588.8600 ;
        RECT 2437.0200 604.7000 2438.6200 605.1800 ;
        RECT 2437.0200 566.6200 2438.6200 567.1000 ;
        RECT 2437.0200 572.0600 2438.6200 572.5400 ;
        RECT 2437.0200 550.3000 2438.6200 550.7800 ;
        RECT 2437.0200 555.7400 2438.6200 556.2200 ;
        RECT 2437.0200 561.1800 2438.6200 561.6600 ;
        RECT 2437.0200 539.4200 2438.6200 539.9000 ;
        RECT 2437.0200 544.8600 2438.6200 545.3400 ;
        RECT 2437.0200 523.1000 2438.6200 523.5800 ;
        RECT 2437.0200 528.5400 2438.6200 529.0200 ;
        RECT 2437.0200 533.9800 2438.6200 534.4600 ;
        RECT 2437.0200 577.5000 2438.6200 577.9800 ;
        RECT 2394.4000 621.0200 2396.0000 621.5000 ;
        RECT 2394.4000 610.1400 2396.0000 610.6200 ;
        RECT 2394.4000 615.5800 2396.0000 616.0600 ;
        RECT 2394.4000 593.8200 2396.0000 594.3000 ;
        RECT 2394.4000 599.2600 2396.0000 599.7400 ;
        RECT 2394.4000 582.9400 2396.0000 583.4200 ;
        RECT 2394.4000 588.3800 2396.0000 588.8600 ;
        RECT 2394.4000 604.7000 2396.0000 605.1800 ;
        RECT 2394.4000 566.6200 2396.0000 567.1000 ;
        RECT 2394.4000 572.0600 2396.0000 572.5400 ;
        RECT 2394.4000 550.3000 2396.0000 550.7800 ;
        RECT 2394.4000 555.7400 2396.0000 556.2200 ;
        RECT 2394.4000 561.1800 2396.0000 561.6600 ;
        RECT 2394.4000 539.4200 2396.0000 539.9000 ;
        RECT 2394.4000 544.8600 2396.0000 545.3400 ;
        RECT 2394.4000 523.1000 2396.0000 523.5800 ;
        RECT 2394.4000 528.5400 2396.0000 529.0200 ;
        RECT 2394.4000 533.9800 2396.0000 534.4600 ;
        RECT 2394.4000 577.5000 2396.0000 577.9800 ;
        RECT 2437.0200 512.2200 2438.6200 512.7000 ;
        RECT 2437.0200 517.6600 2438.6200 518.1400 ;
        RECT 2437.0200 495.9000 2438.6200 496.3800 ;
        RECT 2437.0200 501.3400 2438.6200 501.8200 ;
        RECT 2437.0200 506.7800 2438.6200 507.2600 ;
        RECT 2437.0200 485.0200 2438.6200 485.5000 ;
        RECT 2437.0200 490.4600 2438.6200 490.9400 ;
        RECT 2437.0200 468.7000 2438.6200 469.1800 ;
        RECT 2437.0200 474.1400 2438.6200 474.6200 ;
        RECT 2437.0200 479.5800 2438.6200 480.0600 ;
        RECT 2437.0200 457.8200 2438.6200 458.3000 ;
        RECT 2437.0200 463.2600 2438.6200 463.7400 ;
        RECT 2437.0200 441.5000 2438.6200 441.9800 ;
        RECT 2437.0200 446.9400 2438.6200 447.4200 ;
        RECT 2437.0200 452.3800 2438.6200 452.8600 ;
        RECT 2437.0200 430.6200 2438.6200 431.1000 ;
        RECT 2437.0200 436.0600 2438.6200 436.5400 ;
        RECT 2437.0200 425.1800 2438.6200 425.6600 ;
        RECT 2394.4000 512.2200 2396.0000 512.7000 ;
        RECT 2394.4000 517.6600 2396.0000 518.1400 ;
        RECT 2394.4000 495.9000 2396.0000 496.3800 ;
        RECT 2394.4000 501.3400 2396.0000 501.8200 ;
        RECT 2394.4000 506.7800 2396.0000 507.2600 ;
        RECT 2394.4000 485.0200 2396.0000 485.5000 ;
        RECT 2394.4000 490.4600 2396.0000 490.9400 ;
        RECT 2394.4000 468.7000 2396.0000 469.1800 ;
        RECT 2394.4000 474.1400 2396.0000 474.6200 ;
        RECT 2394.4000 479.5800 2396.0000 480.0600 ;
        RECT 2394.4000 457.8200 2396.0000 458.3000 ;
        RECT 2394.4000 463.2600 2396.0000 463.7400 ;
        RECT 2394.4000 441.5000 2396.0000 441.9800 ;
        RECT 2394.4000 446.9400 2396.0000 447.4200 ;
        RECT 2394.4000 452.3800 2396.0000 452.8600 ;
        RECT 2394.4000 430.6200 2396.0000 431.1000 ;
        RECT 2394.4000 436.0600 2396.0000 436.5400 ;
        RECT 2394.4000 425.1800 2396.0000 425.6600 ;
        RECT 2391.4400 627.3700 2441.5800 628.9700 ;
        RECT 2391.4400 415.6700 2441.5800 417.2700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 412.8400 2396.0000 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.4000 630.8800 2396.0000 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 412.8400 2438.6200 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.0200 630.8800 2438.6200 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 415.6700 2393.0400 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 415.6700 2441.5800 417.2700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 627.3700 2393.0400 628.9700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 627.3700 2441.5800 628.9700 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'wb_mem_split'
    PORT
      LAYER met4 ;
        RECT 521.1600 457.2200 649.4800 458.8200 ;
    END
# end of P/G pin shape extracted from block 'wb_mem_split'

  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER met3 ;
        RECT 2.0000 2.0000 3368.4200 5.0000 ;
        RECT 1283.3400 178.6000 2446.1800 180.2000 ;
        RECT 1283.3400 138.3400 2386.0400 139.9400 ;
        RECT 1283.3400 408.2400 1945.6000 409.8400 ;
        RECT 1283.3400 867.5200 1945.6000 869.1200 ;
        RECT 1283.3400 637.8800 2446.1800 639.4800 ;
        RECT 1283.3400 1097.1600 2446.1800 1098.7600 ;
        RECT 2.0000 178.8600 1285.0800 180.4600 ;
        RECT 656.8450 408.5000 1064.8600 410.1000 ;
        RECT 2.0000 408.5000 516.5150 410.1000 ;
        RECT 1063.2600 138.6000 1285.0800 140.2000 ;
        RECT 1005.5200 188.7900 1010.9200 190.3900 ;
        RECT 1063.2600 147.1700 1071.0600 148.7700 ;
        RECT 1063.2600 166.7000 1071.0600 168.3000 ;
        RECT 1075.8200 193.0800 1077.4200 193.3200 ;
        RECT 1063.2600 188.8900 1071.0600 190.4900 ;
        RECT 1059.4600 188.7900 1064.8600 190.3900 ;
        RECT 1005.5200 395.4900 1010.9200 397.0900 ;
        RECT 1005.5200 418.4300 1010.9200 420.0300 ;
        RECT 1059.4600 395.4900 1064.8600 397.0900 ;
        RECT 1059.4600 418.4300 1064.8600 420.0300 ;
        RECT 1283.3400 146.9100 1291.1400 148.5100 ;
        RECT 1279.6800 147.1700 1285.0800 148.7700 ;
        RECT 1279.6800 166.7000 1285.0800 168.3000 ;
        RECT 1283.3400 166.4400 1291.1400 168.0400 ;
        RECT 1283.3400 188.6300 1291.1400 190.2300 ;
        RECT 1295.9000 192.8200 1297.5000 193.0600 ;
        RECT 1279.6800 188.8900 1285.0800 190.4900 ;
        RECT 1499.7600 146.9100 1505.1600 148.5100 ;
        RECT 1503.5600 146.9100 1511.3600 148.5100 ;
        RECT 1503.5600 166.4400 1511.3600 168.0400 ;
        RECT 1499.7600 166.4400 1505.1600 168.0400 ;
        RECT 1503.5600 188.6300 1511.3600 190.2300 ;
        RECT 1516.1200 192.8200 1517.7200 193.0600 ;
        RECT 1295.9000 422.4600 1297.5000 422.7000 ;
        RECT 1283.3400 395.1300 1291.1400 396.7300 ;
        RECT 1283.3400 418.2700 1291.1400 419.8700 ;
        RECT 1503.5600 395.1300 1511.3600 396.7300 ;
        RECT 1499.7600 395.1300 1505.1600 396.7300 ;
        RECT 1499.7600 418.2700 1505.1600 419.8700 ;
        RECT 1516.1200 422.4600 1517.7200 422.7000 ;
        RECT 1503.5600 418.2700 1511.3600 419.8700 ;
        RECT 2.0000 638.1400 1285.0800 639.7400 ;
        RECT 2.0000 867.7800 167.1150 869.3800 ;
        RECT 2.0000 1097.4200 167.1150 1099.0200 ;
        RECT 1005.5200 625.1300 1010.9200 626.7300 ;
        RECT 1005.5200 648.0700 1010.9200 649.6700 ;
        RECT 1063.2600 626.0800 1071.0600 627.6800 ;
        RECT 1059.4600 625.1300 1064.8600 626.7300 ;
        RECT 1059.4600 648.0700 1064.8600 649.6700 ;
        RECT 1075.8200 652.3600 1077.4200 652.6000 ;
        RECT 1063.2600 648.1700 1071.0600 649.7700 ;
        RECT 1005.5200 854.7700 1010.9200 856.3700 ;
        RECT 1059.4600 854.7700 1064.8600 856.3700 ;
        RECT 1279.6800 626.0800 1285.0800 627.6800 ;
        RECT 1283.3400 624.7700 1291.1400 626.3700 ;
        RECT 1283.3400 647.9100 1291.1400 649.5100 ;
        RECT 1279.6800 648.1700 1285.0800 649.7700 ;
        RECT 1295.9000 652.1000 1297.5000 652.3400 ;
        RECT 1499.7600 624.7700 1505.1600 626.3700 ;
        RECT 1503.5600 624.7700 1511.3600 626.3700 ;
        RECT 1499.7600 647.9100 1505.1600 649.5100 ;
        RECT 1503.5600 647.9100 1511.3600 649.5100 ;
        RECT 1516.1200 652.1000 1517.7200 652.3400 ;
        RECT 1499.7600 854.4100 1505.1600 856.0100 ;
        RECT 1503.5600 854.4100 1511.3600 856.0100 ;
        RECT 1283.3400 854.4100 1291.1400 856.0100 ;
        RECT 953.4450 1097.4200 1285.0800 1099.0200 ;
        RECT 953.4450 867.7800 1064.8600 869.3800 ;
        RECT 1005.5200 877.7100 1010.9200 879.3100 ;
        RECT 1059.4600 877.7100 1064.8600 879.3100 ;
        RECT 1005.5200 1107.3500 1010.9200 1108.9500 ;
        RECT 1005.5200 1084.4100 1010.9200 1086.0100 ;
        RECT 1063.2600 1085.3600 1071.0600 1086.9600 ;
        RECT 1059.4600 1084.4100 1064.8600 1086.0100 ;
        RECT 1063.2600 1107.4500 1071.0600 1109.0500 ;
        RECT 1075.8200 1111.6400 1077.4200 1111.8800 ;
        RECT 1059.4600 1107.3500 1064.8600 1108.9500 ;
        RECT 1283.3400 877.5500 1291.1400 879.1500 ;
        RECT 1295.9000 881.7400 1297.5000 881.9800 ;
        RECT 1499.7600 877.5500 1505.1600 879.1500 ;
        RECT 1503.5600 877.5500 1511.3600 879.1500 ;
        RECT 1516.1200 881.7400 1517.7200 881.9800 ;
        RECT 1279.6800 1085.3600 1285.0800 1086.9600 ;
        RECT 1283.3400 1084.0500 1291.1400 1085.6500 ;
        RECT 1279.6800 1107.4500 1285.0800 1109.0500 ;
        RECT 1283.3400 1107.1900 1291.1400 1108.7900 ;
        RECT 1295.9000 1111.3800 1297.5000 1111.6200 ;
        RECT 1499.7600 1084.0500 1505.1600 1085.6500 ;
        RECT 1503.5600 1084.0500 1511.3600 1085.6500 ;
        RECT 1499.7600 1107.1900 1505.1600 1108.7900 ;
        RECT 1503.5600 1107.1900 1511.3600 1108.7900 ;
        RECT 1516.1200 1111.3800 1517.7200 1111.6200 ;
        RECT 1723.7800 146.9100 1731.5800 148.5100 ;
        RECT 1719.9800 146.9100 1725.3800 148.5100 ;
        RECT 1719.9800 166.4400 1725.3800 168.0400 ;
        RECT 1723.7800 166.4400 1731.5800 168.0400 ;
        RECT 1723.7800 188.6300 1731.5800 190.2300 ;
        RECT 1736.3400 192.8200 1737.9400 193.0600 ;
        RECT 1944.0000 146.9100 1951.8000 148.5100 ;
        RECT 1944.0000 166.4400 1951.8000 168.0400 ;
        RECT 1940.2000 146.9100 1945.6000 148.5100 ;
        RECT 1940.2000 166.4400 1945.6000 168.0400 ;
        RECT 1944.0000 188.6300 1951.8000 190.2300 ;
        RECT 1956.5600 192.8200 1958.1600 193.0600 ;
        RECT 1736.3400 422.4600 1737.9400 422.7000 ;
        RECT 1719.9800 418.2700 1725.3800 419.8700 ;
        RECT 1723.7800 418.2700 1731.5800 419.8700 ;
        RECT 1719.9800 395.1300 1725.3800 396.7300 ;
        RECT 1723.7800 395.1300 1731.5800 396.7300 ;
        RECT 1940.2000 418.2700 1945.6000 419.8700 ;
        RECT 1940.2000 395.1300 1945.6000 396.7300 ;
        RECT 2164.2200 146.9100 2172.0200 148.5100 ;
        RECT 2160.4200 146.9100 2165.8200 148.5100 ;
        RECT 2160.4200 166.4400 2165.8200 168.0400 ;
        RECT 2164.2200 166.4400 2172.0200 168.0400 ;
        RECT 2160.4200 188.6300 2165.8200 190.2300 ;
        RECT 2164.2200 188.6300 2172.0200 190.2300 ;
        RECT 2176.7800 192.8200 2178.3800 193.0600 ;
        RECT 2380.6400 146.9100 2386.0400 148.5100 ;
        RECT 2380.6400 166.4400 2386.0400 168.0400 ;
        RECT 2384.4400 188.6300 2392.2400 190.2300 ;
        RECT 2440.7800 188.6300 2446.1800 190.2300 ;
        RECT 2164.2200 408.2400 2446.1800 409.8400 ;
        RECT 2164.2200 395.1300 2172.0200 396.7300 ;
        RECT 2176.7800 422.4600 2178.3800 422.7000 ;
        RECT 2164.2200 418.2700 2172.0200 419.8700 ;
        RECT 2384.4400 395.1300 2392.2400 396.7300 ;
        RECT 2380.6400 395.1300 2386.0400 396.7300 ;
        RECT 2384.4400 418.2700 2392.2400 419.8700 ;
        RECT 2380.6400 418.2700 2386.0400 419.8700 ;
        RECT 2440.7800 395.1300 2446.1800 396.7300 ;
        RECT 2440.7800 418.2700 2446.1800 419.8700 ;
        RECT 1736.3400 652.1000 1737.9400 652.3400 ;
        RECT 1723.7800 624.7700 1731.5800 626.3700 ;
        RECT 1723.7800 647.9100 1731.5800 649.5100 ;
        RECT 1719.9800 647.9100 1725.3800 649.5100 ;
        RECT 1719.9800 624.7700 1725.3800 626.3700 ;
        RECT 1944.0000 625.8200 1951.8000 627.4200 ;
        RECT 1944.0000 647.9100 1951.8000 649.5100 ;
        RECT 1940.2000 647.9100 1945.6000 649.5100 ;
        RECT 1940.2000 624.7700 1945.6000 626.3700 ;
        RECT 1956.5600 652.1000 1958.1600 652.3400 ;
        RECT 1940.2000 854.4100 1945.6000 856.0100 ;
        RECT 1723.7800 854.4100 1731.5800 856.0100 ;
        RECT 1719.9800 854.4100 1725.3800 856.0100 ;
        RECT 2160.4200 625.8200 2165.8200 627.4200 ;
        RECT 2164.2200 624.7700 2172.0200 626.3700 ;
        RECT 2160.4200 647.9100 2165.8200 649.5100 ;
        RECT 2164.2200 647.9100 2172.0200 649.5100 ;
        RECT 2176.7800 652.1000 2178.3800 652.3400 ;
        RECT 2384.4400 647.9100 2392.2400 649.5100 ;
        RECT 2380.6400 647.9100 2386.0400 649.5100 ;
        RECT 2384.4400 624.7700 2392.2400 626.3700 ;
        RECT 2380.6400 624.7700 2386.0400 626.3700 ;
        RECT 2440.7800 624.7700 2446.1800 626.3700 ;
        RECT 2440.7800 647.9100 2446.1800 649.5100 ;
        RECT 2164.2200 854.4100 2172.0200 856.0100 ;
        RECT 2440.7800 854.4100 2446.1800 856.0100 ;
        RECT 2384.4400 854.4100 2392.2400 856.0100 ;
        RECT 2380.6400 854.4100 2386.0400 856.0100 ;
        RECT 1719.9800 877.5500 1725.3800 879.1500 ;
        RECT 1723.7800 877.5500 1731.5800 879.1500 ;
        RECT 1736.3400 881.7400 1737.9400 881.9800 ;
        RECT 1940.2000 877.5500 1945.6000 879.1500 ;
        RECT 1736.3400 1111.3800 1737.9400 1111.6200 ;
        RECT 1723.7800 1107.1900 1731.5800 1108.7900 ;
        RECT 1719.9800 1107.1900 1725.3800 1108.7900 ;
        RECT 1723.7800 1084.0500 1731.5800 1085.6500 ;
        RECT 1719.9800 1084.0500 1725.3800 1085.6500 ;
        RECT 1944.0000 1085.1000 1951.8000 1086.7000 ;
        RECT 1944.0000 1107.1900 1951.8000 1108.7900 ;
        RECT 1940.2000 1107.1900 1945.6000 1108.7900 ;
        RECT 1940.2000 1084.0500 1945.6000 1085.6500 ;
        RECT 1956.5600 1111.3800 1958.1600 1111.6200 ;
        RECT 2164.2200 867.5200 2446.1800 869.1200 ;
        RECT 2164.2200 877.5500 2172.0200 879.1500 ;
        RECT 2176.7800 881.7400 2178.3800 881.9800 ;
        RECT 2380.6400 877.5500 2386.0400 879.1500 ;
        RECT 2384.4400 877.5500 2392.2400 879.1500 ;
        RECT 2440.7800 877.5500 2446.1800 879.1500 ;
        RECT 2160.4200 1085.1000 2165.8200 1086.7000 ;
        RECT 2164.2200 1084.0500 2172.0200 1085.6500 ;
        RECT 2160.4200 1107.1900 2165.8200 1108.7900 ;
        RECT 2176.7800 1111.3800 2178.3800 1111.6200 ;
        RECT 2164.2200 1107.1900 2172.0200 1108.7900 ;
        RECT 2380.6400 1107.1900 2386.0400 1108.7900 ;
        RECT 2384.4400 1107.1900 2392.2400 1108.7900 ;
        RECT 2384.4400 1084.0500 2392.2400 1085.6500 ;
        RECT 2380.6400 1084.0500 2386.0400 1085.6500 ;
        RECT 2440.7800 1107.1900 2446.1800 1108.7900 ;
        RECT 2440.7800 1084.0500 2446.1800 1085.6500 ;
        RECT 2.0000 2564.7200 3368.4200 2567.7200 ;
        RECT 1063.2600 2475.0000 2386.0400 2476.6000 ;
        RECT 1283.3400 2015.7200 2446.1800 2017.3200 ;
        RECT 1283.3400 1556.4400 2446.1800 1558.0400 ;
        RECT 1283.3400 2245.3600 1945.6000 2246.9600 ;
        RECT 1283.3400 1786.0800 1945.6000 1787.6800 ;
        RECT 1283.3400 1326.8000 1945.6000 1328.4000 ;
        RECT 2.0000 2015.9800 1285.0800 2017.5800 ;
        RECT 2.0000 1327.0600 167.1150 1328.6600 ;
        RECT 2.0000 1556.7000 167.1150 1558.3000 ;
        RECT 2.0000 1786.3400 167.1150 1787.9400 ;
        RECT 953.4450 1556.7000 1285.0800 1558.3000 ;
        RECT 953.4450 1327.0600 1064.8600 1328.6600 ;
        RECT 1005.5200 1314.0500 1010.9200 1315.6500 ;
        RECT 1005.5200 1336.9900 1010.9200 1338.5900 ;
        RECT 1059.4600 1314.0500 1064.8600 1315.6500 ;
        RECT 1059.4600 1336.9900 1064.8600 1338.5900 ;
        RECT 1005.5200 1543.6900 1010.9200 1545.2900 ;
        RECT 1005.5200 1566.6300 1010.9200 1568.2300 ;
        RECT 1059.4600 1543.6900 1064.8600 1545.2900 ;
        RECT 1063.2600 1544.6400 1071.0600 1546.2400 ;
        RECT 1075.8200 1570.9200 1077.4200 1571.1600 ;
        RECT 1063.2600 1566.7300 1071.0600 1568.3300 ;
        RECT 1059.4600 1566.6300 1064.8600 1568.2300 ;
        RECT 1295.9000 1341.0200 1297.5000 1341.2600 ;
        RECT 1283.3400 1336.8300 1291.1400 1338.4300 ;
        RECT 1283.3400 1313.6900 1291.1400 1315.2900 ;
        RECT 1503.5600 1336.8300 1511.3600 1338.4300 ;
        RECT 1499.7600 1336.8300 1505.1600 1338.4300 ;
        RECT 1499.7600 1313.6900 1505.1600 1315.2900 ;
        RECT 1503.5600 1313.6900 1511.3600 1315.2900 ;
        RECT 1516.1200 1341.0200 1517.7200 1341.2600 ;
        RECT 1279.6800 1544.6400 1285.0800 1546.2400 ;
        RECT 1283.3400 1543.3300 1291.1400 1544.9300 ;
        RECT 1279.6800 1566.7300 1285.0800 1568.3300 ;
        RECT 1283.3400 1566.4700 1291.1400 1568.0700 ;
        RECT 1295.9000 1570.6600 1297.5000 1570.9000 ;
        RECT 1499.7600 1543.3300 1505.1600 1544.9300 ;
        RECT 1503.5600 1543.3300 1511.3600 1544.9300 ;
        RECT 1499.7600 1566.4700 1505.1600 1568.0700 ;
        RECT 1503.5600 1566.4700 1511.3600 1568.0700 ;
        RECT 1516.1200 1570.6600 1517.7200 1570.9000 ;
        RECT 953.4450 1786.3400 1064.8600 1787.9400 ;
        RECT 1005.5200 1796.2700 1010.9200 1797.8700 ;
        RECT 1005.5200 1773.3300 1010.9200 1774.9300 ;
        RECT 1059.4600 1796.2700 1064.8600 1797.8700 ;
        RECT 1059.4600 1773.3300 1064.8600 1774.9300 ;
        RECT 1005.5200 2002.9700 1010.9200 2004.5700 ;
        RECT 1005.5200 2025.9100 1010.9200 2027.5100 ;
        RECT 1059.4600 2002.9700 1064.8600 2004.5700 ;
        RECT 1063.2600 2003.9200 1071.0600 2005.5200 ;
        RECT 1059.4600 2025.9100 1064.8600 2027.5100 ;
        RECT 1063.2600 2026.0100 1071.0600 2027.6100 ;
        RECT 1075.8200 2030.2000 1077.4200 2030.4400 ;
        RECT 1295.9000 1800.3000 1297.5000 1800.5400 ;
        RECT 1283.3400 1772.9700 1291.1400 1774.5700 ;
        RECT 1283.3400 1796.1100 1291.1400 1797.7100 ;
        RECT 1503.5600 1772.9700 1511.3600 1774.5700 ;
        RECT 1499.7600 1772.9700 1505.1600 1774.5700 ;
        RECT 1499.7600 1796.1100 1505.1600 1797.7100 ;
        RECT 1516.1200 1800.3000 1517.7200 1800.5400 ;
        RECT 1503.5600 1796.1100 1511.3600 1797.7100 ;
        RECT 1279.6800 2003.9200 1285.0800 2005.5200 ;
        RECT 1283.3400 2002.6100 1291.1400 2004.2100 ;
        RECT 1279.6800 2026.0100 1285.0800 2027.6100 ;
        RECT 1283.3400 2025.7500 1291.1400 2027.3500 ;
        RECT 1295.9000 2029.9400 1297.5000 2030.1800 ;
        RECT 1503.5600 2002.6100 1511.3600 2004.2100 ;
        RECT 1499.7600 2002.6100 1505.1600 2004.2100 ;
        RECT 1499.7600 2025.7500 1505.1600 2027.3500 ;
        RECT 1516.1200 2029.9400 1517.7200 2030.1800 ;
        RECT 1503.5600 2025.7500 1511.3600 2027.3500 ;
        RECT 2.0000 2245.6200 1064.8600 2247.2200 ;
        RECT 1005.5200 2232.6100 1010.9200 2234.2100 ;
        RECT 1005.5200 2255.5500 1010.9200 2257.1500 ;
        RECT 1059.4600 2255.5500 1064.8600 2257.1500 ;
        RECT 1059.4600 2232.6100 1064.8600 2234.2100 ;
        RECT 1005.5200 2462.2500 1010.9200 2463.8500 ;
        RECT 1063.2600 2463.2000 1071.0600 2464.8000 ;
        RECT 1059.4600 2462.2500 1064.8600 2463.8500 ;
        RECT 1063.2600 2483.5700 1070.9200 2485.1700 ;
        RECT 1063.2600 2503.1000 1070.9200 2504.7000 ;
        RECT 1295.9000 2259.5800 1297.5000 2259.8200 ;
        RECT 1283.3400 2255.3900 1291.1400 2256.9900 ;
        RECT 1283.3400 2232.2500 1291.1400 2233.8500 ;
        RECT 1499.7600 2232.2500 1505.1600 2233.8500 ;
        RECT 1503.5600 2232.2500 1511.3600 2233.8500 ;
        RECT 1503.5600 2255.3900 1511.3600 2256.9900 ;
        RECT 1516.1200 2259.5800 1517.7200 2259.8200 ;
        RECT 1499.7600 2255.3900 1505.1600 2256.9900 ;
        RECT 1279.6800 2463.2000 1285.0800 2464.8000 ;
        RECT 1283.3400 2461.8900 1291.1400 2463.4900 ;
        RECT 1283.3400 2483.5700 1291.1400 2485.1700 ;
        RECT 1279.5400 2483.5700 1285.0800 2485.1700 ;
        RECT 1279.5400 2503.1000 1285.0800 2504.7000 ;
        RECT 1283.3400 2503.1000 1291.1400 2504.7000 ;
        RECT 1503.5600 2461.8900 1511.3600 2463.4900 ;
        RECT 1499.7600 2461.8900 1505.1600 2463.4900 ;
        RECT 1503.5600 2483.5700 1511.3600 2485.1700 ;
        RECT 1499.7600 2483.5700 1505.1600 2485.1700 ;
        RECT 1499.7600 2503.1000 1505.1600 2504.7000 ;
        RECT 1503.5600 2503.1000 1511.3600 2504.7000 ;
        RECT 1719.9800 1336.8300 1725.3800 1338.4300 ;
        RECT 1723.7800 1336.8300 1731.5800 1338.4300 ;
        RECT 1719.9800 1313.6900 1725.3800 1315.2900 ;
        RECT 1723.7800 1313.6900 1731.5800 1315.2900 ;
        RECT 1736.3400 1341.0200 1737.9400 1341.2600 ;
        RECT 1940.2000 1336.8300 1945.6000 1338.4300 ;
        RECT 1940.2000 1313.6900 1945.6000 1315.2900 ;
        RECT 1719.9800 1543.3300 1725.3800 1544.9300 ;
        RECT 1723.7800 1543.3300 1731.5800 1544.9300 ;
        RECT 1723.7800 1566.4700 1731.5800 1568.0700 ;
        RECT 1736.3400 1570.6600 1737.9400 1570.9000 ;
        RECT 1719.9800 1566.4700 1725.3800 1568.0700 ;
        RECT 1944.0000 1544.3800 1951.8000 1545.9800 ;
        RECT 1940.2000 1543.3300 1945.6000 1544.9300 ;
        RECT 1944.0000 1566.4700 1951.8000 1568.0700 ;
        RECT 1940.2000 1566.4700 1945.6000 1568.0700 ;
        RECT 1956.5600 1570.6600 1958.1600 1570.9000 ;
        RECT 2164.2200 1326.8000 2446.1800 1328.4000 ;
        RECT 2176.7800 1341.0200 2178.3800 1341.2600 ;
        RECT 2164.2200 1313.6900 2172.0200 1315.2900 ;
        RECT 2164.2200 1336.8300 2172.0200 1338.4300 ;
        RECT 2384.4400 1336.8300 2392.2400 1338.4300 ;
        RECT 2384.4400 1313.6900 2392.2400 1315.2900 ;
        RECT 2380.6400 1336.8300 2386.0400 1338.4300 ;
        RECT 2380.6400 1313.6900 2386.0400 1315.2900 ;
        RECT 2440.7800 1336.8300 2446.1800 1338.4300 ;
        RECT 2440.7800 1313.6900 2446.1800 1315.2900 ;
        RECT 2160.4200 1544.3800 2165.8200 1545.9800 ;
        RECT 2164.2200 1543.3300 2172.0200 1544.9300 ;
        RECT 2160.4200 1566.4700 2165.8200 1568.0700 ;
        RECT 2164.2200 1566.4700 2172.0200 1568.0700 ;
        RECT 2176.7800 1570.6600 2178.3800 1570.9000 ;
        RECT 2384.4400 1566.4700 2392.2400 1568.0700 ;
        RECT 2380.6400 1566.4700 2386.0400 1568.0700 ;
        RECT 2380.6400 1543.3300 2386.0400 1544.9300 ;
        RECT 2384.4400 1543.3300 2392.2400 1544.9300 ;
        RECT 2440.7800 1566.4700 2446.1800 1568.0700 ;
        RECT 2440.7800 1543.3300 2446.1800 1544.9300 ;
        RECT 1736.3400 1800.3000 1737.9400 1800.5400 ;
        RECT 1719.9800 1796.1100 1725.3800 1797.7100 ;
        RECT 1719.9800 1772.9700 1725.3800 1774.5700 ;
        RECT 1723.7800 1772.9700 1731.5800 1774.5700 ;
        RECT 1723.7800 1796.1100 1731.5800 1797.7100 ;
        RECT 1940.2000 1796.1100 1945.6000 1797.7100 ;
        RECT 1940.2000 1772.9700 1945.6000 1774.5700 ;
        RECT 1723.7800 2002.6100 1731.5800 2004.2100 ;
        RECT 1719.9800 2002.6100 1725.3800 2004.2100 ;
        RECT 1719.9800 2025.7500 1725.3800 2027.3500 ;
        RECT 1736.3400 2029.9400 1737.9400 2030.1800 ;
        RECT 1723.7800 2025.7500 1731.5800 2027.3500 ;
        RECT 1944.0000 2003.6600 1951.8000 2005.2600 ;
        RECT 1940.2000 2002.6100 1945.6000 2004.2100 ;
        RECT 1944.0000 2025.7500 1951.8000 2027.3500 ;
        RECT 1956.5600 2029.9400 1958.1600 2030.1800 ;
        RECT 1940.2000 2025.7500 1945.6000 2027.3500 ;
        RECT 2164.2200 1786.0800 2446.1800 1787.6800 ;
        RECT 2176.7800 1800.3000 2178.3800 1800.5400 ;
        RECT 2164.2200 1772.9700 2172.0200 1774.5700 ;
        RECT 2164.2200 1796.1100 2172.0200 1797.7100 ;
        RECT 2384.4400 1772.9700 2392.2400 1774.5700 ;
        RECT 2380.6400 1772.9700 2386.0400 1774.5700 ;
        RECT 2380.6400 1796.1100 2386.0400 1797.7100 ;
        RECT 2384.4400 1796.1100 2392.2400 1797.7100 ;
        RECT 2440.7800 1772.9700 2446.1800 1774.5700 ;
        RECT 2440.7800 1796.1100 2446.1800 1797.7100 ;
        RECT 2160.4200 2003.6600 2165.8200 2005.2600 ;
        RECT 2164.2200 2002.6100 2172.0200 2004.2100 ;
        RECT 2160.4200 2025.7500 2165.8200 2027.3500 ;
        RECT 2164.2200 2025.7500 2172.0200 2027.3500 ;
        RECT 2176.7800 2029.9400 2178.3800 2030.1800 ;
        RECT 2380.6400 2002.6100 2386.0400 2004.2100 ;
        RECT 2384.4400 2002.6100 2392.2400 2004.2100 ;
        RECT 2440.7800 2002.6100 2446.1800 2004.2100 ;
        RECT 2384.4400 2025.7500 2392.2400 2027.3500 ;
        RECT 2380.6400 2025.7500 2386.0400 2027.3500 ;
        RECT 2440.7800 2025.7500 2446.1800 2027.3500 ;
        RECT 1719.9800 2232.2500 1725.3800 2233.8500 ;
        RECT 1723.7800 2232.2500 1731.5800 2233.8500 ;
        RECT 1736.3400 2259.5800 1737.9400 2259.8200 ;
        RECT 1719.9800 2255.3900 1725.3800 2256.9900 ;
        RECT 1723.7800 2255.3900 1731.5800 2256.9900 ;
        RECT 1940.2000 2232.2500 1945.6000 2233.8500 ;
        RECT 1940.2000 2255.3900 1945.6000 2256.9900 ;
        RECT 1723.7800 2461.8900 1731.5800 2463.4900 ;
        RECT 1719.9800 2461.8900 1725.3800 2463.4900 ;
        RECT 1723.7800 2483.5700 1731.5800 2485.1700 ;
        RECT 1719.9800 2483.5700 1725.3800 2485.1700 ;
        RECT 1723.7800 2503.1000 1731.5800 2504.7000 ;
        RECT 1719.9800 2503.1000 1725.3800 2504.7000 ;
        RECT 1944.0000 2483.5700 1951.8000 2485.1700 ;
        RECT 1944.0000 2462.9400 1951.8000 2464.5400 ;
        RECT 1940.2000 2461.8900 1945.6000 2463.4900 ;
        RECT 1940.2000 2483.5700 1945.6000 2485.1700 ;
        RECT 1944.0000 2503.1000 1951.8000 2504.7000 ;
        RECT 1940.2000 2503.1000 1945.6000 2504.7000 ;
        RECT 2164.2200 2245.3600 2446.1800 2246.9600 ;
        RECT 2176.7800 2259.5800 2178.3800 2259.8200 ;
        RECT 2164.2200 2255.3900 2172.0200 2256.9900 ;
        RECT 2164.2200 2232.2500 2172.0200 2233.8500 ;
        RECT 2440.7800 2232.2500 2446.1800 2233.8500 ;
        RECT 2384.4400 2232.2500 2392.2400 2233.8500 ;
        RECT 2380.6400 2232.2500 2386.0400 2233.8500 ;
        RECT 2384.4400 2255.3900 2392.2400 2256.9900 ;
        RECT 2380.6400 2255.3900 2386.0400 2256.9900 ;
        RECT 2440.7800 2255.3900 2446.1800 2256.9900 ;
        RECT 2160.4200 2462.9400 2165.8200 2464.5400 ;
        RECT 2164.2200 2461.8900 2172.0200 2463.4900 ;
        RECT 2164.2200 2483.5700 2172.0200 2485.1700 ;
        RECT 2160.4200 2483.5700 2165.8200 2485.1700 ;
        RECT 2160.4200 2503.1000 2165.8200 2504.7000 ;
        RECT 2164.2200 2503.1000 2172.0200 2504.7000 ;
        RECT 2384.4400 2461.8900 2392.2400 2463.4900 ;
        RECT 2380.6400 2461.8900 2386.0400 2463.4900 ;
        RECT 2380.6400 2483.5700 2386.0400 2485.1700 ;
        RECT 2380.6400 2503.1000 2386.0400 2504.7000 ;
        RECT 2440.7800 2461.8900 2446.1800 2463.4900 ;
        RECT 2.0000 20.5000 5.0000 20.9800 ;
        RECT 2.0000 9.6200 5.0000 10.1000 ;
        RECT 2.0000 15.0600 5.0000 15.5400 ;
        RECT 2.0000 25.9400 5.0000 26.4200 ;
        RECT 2.0000 31.3800 5.0000 31.8600 ;
        RECT 2.0000 36.8200 5.0000 37.3000 ;
        RECT 2.0000 42.2600 5.0000 42.7400 ;
        RECT 2.0000 47.7000 5.0000 48.1800 ;
        RECT 2.0000 53.1400 5.0000 53.6200 ;
        RECT 2.0000 58.5800 5.0000 59.0600 ;
        RECT 2.0000 64.0200 5.0000 64.5000 ;
        RECT 2.0000 69.4600 5.0000 69.9400 ;
        RECT 2.0000 74.9000 5.0000 75.3800 ;
        RECT 2.0000 80.3400 5.0000 80.8200 ;
        RECT 2.0000 85.7800 5.0000 86.2600 ;
        RECT 2.0000 91.2200 5.0000 91.7000 ;
        RECT 2.0000 96.6600 5.0000 97.1400 ;
        RECT 2.0000 112.9800 5.0000 113.4600 ;
        RECT 2.0000 102.1000 5.0000 102.5800 ;
        RECT 2.0000 107.5400 5.0000 108.0200 ;
        RECT 2.0000 118.4200 5.0000 118.9000 ;
        RECT 2.0000 123.8600 5.0000 124.3400 ;
        RECT 2.0000 178.4300 5.0000 180.4600 ;
        RECT 2.0000 129.3000 5.0000 129.7800 ;
        RECT 2.0000 134.7400 5.0000 135.2200 ;
        RECT 2.0000 140.1800 5.0000 140.6600 ;
        RECT 2.0000 145.6200 5.0000 146.1000 ;
        RECT 2.0000 151.0600 5.0000 151.5400 ;
        RECT 2.0000 156.5000 5.0000 156.9800 ;
        RECT 2.0000 161.9400 5.0000 162.4200 ;
        RECT 2.0000 167.3800 5.0000 167.8600 ;
        RECT 2.0000 172.8200 5.0000 173.3000 ;
        RECT 2.0000 183.7000 5.0000 184.1800 ;
        RECT 2.0000 189.1400 5.0000 189.6200 ;
        RECT 2.0000 194.5800 5.0000 195.0600 ;
        RECT 2.0000 200.0200 5.0000 200.5000 ;
        RECT 2.0000 205.4600 5.0000 205.9400 ;
        RECT 2.0000 210.9000 5.0000 211.3800 ;
        RECT 2.0000 216.3400 5.0000 216.8200 ;
        RECT 2.0000 221.7800 5.0000 222.2600 ;
        RECT 2.0000 227.2200 5.0000 227.7000 ;
        RECT 2.0000 232.6600 5.0000 233.1400 ;
        RECT 2.0000 238.1000 5.0000 238.5800 ;
        RECT 2.0000 243.5400 5.0000 244.0200 ;
        RECT 2.0000 248.9800 5.0000 249.4600 ;
        RECT 2.0000 254.4200 5.0000 254.9000 ;
        RECT 2.0000 270.7400 5.0000 271.2200 ;
        RECT 2.0000 259.8600 5.0000 260.3400 ;
        RECT 2.0000 265.3000 5.0000 265.7800 ;
        RECT 2.0000 276.1800 5.0000 276.6600 ;
        RECT 2.0000 281.6200 5.0000 282.1000 ;
        RECT 2.0000 287.0600 5.0000 287.5400 ;
        RECT 2.0000 292.5000 5.0000 292.9800 ;
        RECT 2.0000 297.9400 5.0000 298.4200 ;
        RECT 2.0000 303.3800 5.0000 303.8600 ;
        RECT 2.0000 308.8200 5.0000 309.3000 ;
        RECT 2.0000 314.2600 5.0000 314.7400 ;
        RECT 2.0000 319.7000 5.0000 320.1800 ;
        RECT 2.0000 325.1400 5.0000 325.6200 ;
        RECT 2.0000 330.5800 5.0000 331.0600 ;
        RECT 2.0000 336.0200 5.0000 336.5000 ;
        RECT 2.0000 363.2200 5.0000 363.7000 ;
        RECT 2.0000 341.4600 5.0000 341.9400 ;
        RECT 2.0000 346.9000 5.0000 347.3800 ;
        RECT 2.0000 352.3400 5.0000 352.8200 ;
        RECT 2.0000 357.7800 5.0000 358.2600 ;
        RECT 2.0000 368.6600 5.0000 369.1400 ;
        RECT 2.0000 374.1000 5.0000 374.5800 ;
        RECT 2.0000 379.5400 5.0000 380.0200 ;
        RECT 2.0000 384.9800 5.0000 385.4600 ;
        RECT 2.0000 390.4200 5.0000 390.9000 ;
        RECT 2.0000 395.8600 5.0000 396.3400 ;
        RECT 2.0000 401.3000 5.0000 401.7800 ;
        RECT 2.0000 406.7400 5.0000 407.2200 ;
        RECT 2.0000 412.1800 5.0000 412.6600 ;
        RECT 2.0000 417.6200 5.0000 418.1000 ;
        RECT 2.0000 423.0600 5.0000 423.5400 ;
        RECT 2.0000 428.5000 5.0000 428.9800 ;
        RECT 2.0000 433.9400 5.0000 434.4200 ;
        RECT 2.0000 439.3800 5.0000 439.8600 ;
        RECT 505.5200 183.7000 507.1200 184.1800 ;
        RECT 505.5200 189.1400 507.1200 189.6200 ;
        RECT 505.5200 194.5800 507.1200 195.0600 ;
        RECT 505.5200 200.0200 507.1200 200.5000 ;
        RECT 505.5200 205.4600 507.1200 205.9400 ;
        RECT 505.5200 210.9000 507.1200 211.3800 ;
        RECT 505.5200 216.3400 507.1200 216.8200 ;
        RECT 505.5200 221.7800 507.1200 222.2600 ;
        RECT 505.5200 227.2200 507.1200 227.7000 ;
        RECT 663.1200 183.7000 664.7200 184.1800 ;
        RECT 663.1200 189.1400 664.7200 189.6200 ;
        RECT 663.1200 194.5800 664.7200 195.0600 ;
        RECT 663.1200 200.0200 664.7200 200.5000 ;
        RECT 663.1200 205.4600 664.7200 205.9400 ;
        RECT 663.1200 210.9000 664.7200 211.3800 ;
        RECT 663.1200 216.3400 664.7200 216.8200 ;
        RECT 663.1200 221.7800 664.7200 222.2600 ;
        RECT 663.1200 227.2200 664.7200 227.7000 ;
        RECT 505.5200 232.6600 507.1200 233.1400 ;
        RECT 505.5200 238.1000 507.1200 238.5800 ;
        RECT 505.5200 243.5400 507.1200 244.0200 ;
        RECT 505.5200 248.9800 507.1200 249.4600 ;
        RECT 505.5200 254.4200 507.1200 254.9000 ;
        RECT 505.5200 270.7400 507.1200 271.2200 ;
        RECT 505.5200 259.8600 507.1200 260.3400 ;
        RECT 505.5200 265.3000 507.1200 265.7800 ;
        RECT 505.5200 276.1800 507.1200 276.6600 ;
        RECT 505.5200 281.6200 507.1200 282.1000 ;
        RECT 505.5200 287.0600 507.1200 287.5400 ;
        RECT 505.5200 292.5000 507.1200 292.9800 ;
        RECT 505.5200 297.9400 507.1200 298.4200 ;
        RECT 505.5200 303.3800 507.1200 303.8600 ;
        RECT 505.5200 308.8200 507.1200 309.3000 ;
        RECT 505.5200 314.2600 507.1200 314.7400 ;
        RECT 505.5200 319.7000 507.1200 320.1800 ;
        RECT 505.5200 325.1400 507.1200 325.6200 ;
        RECT 505.5200 330.5800 507.1200 331.0600 ;
        RECT 505.5200 336.0200 507.1200 336.5000 ;
        RECT 505.5200 363.2200 507.1200 363.7000 ;
        RECT 505.5200 341.4600 507.1200 341.9400 ;
        RECT 505.5200 346.9000 507.1200 347.3800 ;
        RECT 505.5200 352.3400 507.1200 352.8200 ;
        RECT 505.5200 357.7800 507.1200 358.2600 ;
        RECT 505.5200 368.6600 507.1200 369.1400 ;
        RECT 505.5200 374.1000 507.1200 374.5800 ;
        RECT 505.5200 379.5400 507.1200 380.0200 ;
        RECT 505.5200 384.9800 507.1200 385.4600 ;
        RECT 505.5200 390.4200 507.1200 390.9000 ;
        RECT 505.5200 395.8600 507.1200 396.3400 ;
        RECT 505.5200 401.3000 507.1200 401.7800 ;
        RECT 505.5200 408.1200 507.1200 410.1000 ;
        RECT 505.5200 412.1800 507.1200 412.6600 ;
        RECT 505.5200 417.6200 507.1200 418.1000 ;
        RECT 505.5200 423.0600 507.1200 423.5400 ;
        RECT 505.5200 428.5000 507.1200 428.9800 ;
        RECT 505.5200 433.9400 507.1200 434.4200 ;
        RECT 505.5200 439.3800 507.1200 439.8600 ;
        RECT 663.1200 232.6600 664.7200 233.1400 ;
        RECT 663.1200 238.1000 664.7200 238.5800 ;
        RECT 663.1200 243.5400 664.7200 244.0200 ;
        RECT 663.1200 248.9800 664.7200 249.4600 ;
        RECT 663.1200 254.4200 664.7200 254.9000 ;
        RECT 663.1200 270.7400 664.7200 271.2200 ;
        RECT 663.1200 259.8600 664.7200 260.3400 ;
        RECT 663.1200 265.3000 664.7200 265.7800 ;
        RECT 663.1200 276.1800 664.7200 276.6600 ;
        RECT 663.1200 281.6200 664.7200 282.1000 ;
        RECT 663.1200 287.0600 664.7200 287.5400 ;
        RECT 663.1200 292.5000 664.7200 292.9800 ;
        RECT 663.1200 297.9400 664.7200 298.4200 ;
        RECT 663.1200 303.3800 664.7200 303.8600 ;
        RECT 663.1200 308.8200 664.7200 309.3000 ;
        RECT 663.1200 314.2600 664.7200 314.7400 ;
        RECT 663.1200 319.7000 664.7200 320.1800 ;
        RECT 663.1200 325.1400 664.7200 325.6200 ;
        RECT 663.1200 330.5800 664.7200 331.0600 ;
        RECT 663.1200 336.0200 664.7200 336.5000 ;
        RECT 663.1200 363.2200 664.7200 363.7000 ;
        RECT 663.1200 341.4600 664.7200 341.9400 ;
        RECT 663.1200 346.9000 664.7200 347.3800 ;
        RECT 663.1200 352.3400 664.7200 352.8200 ;
        RECT 663.1200 357.7800 664.7200 358.2600 ;
        RECT 663.1200 368.6600 664.7200 369.1400 ;
        RECT 663.1200 374.1000 664.7200 374.5800 ;
        RECT 663.1200 379.5400 664.7200 380.0200 ;
        RECT 663.1200 384.9800 664.7200 385.4600 ;
        RECT 663.1200 390.4200 664.7200 390.9000 ;
        RECT 663.1200 395.8600 664.7200 396.3400 ;
        RECT 663.1200 401.3000 664.7200 401.7800 ;
        RECT 663.1200 408.1200 664.7200 410.1000 ;
        RECT 663.1200 412.1800 664.7200 412.6600 ;
        RECT 663.1200 417.6200 664.7200 418.1000 ;
        RECT 663.1200 423.0600 664.7200 423.5400 ;
        RECT 663.1200 428.5000 664.7200 428.9800 ;
        RECT 663.1200 433.9400 664.7200 434.4200 ;
        RECT 663.1200 439.3800 664.7200 439.8600 ;
        RECT 1063.2600 20.5000 1064.8600 20.9800 ;
        RECT 1283.3400 20.5000 1285.0800 20.9800 ;
        RECT 1503.5600 20.5000 1505.1600 20.9800 ;
        RECT 1063.2600 15.0600 1064.8600 15.5400 ;
        RECT 1283.3400 9.6200 1285.0800 10.1000 ;
        RECT 1283.3400 15.0600 1285.0800 15.5400 ;
        RECT 1503.5600 9.6200 1505.1600 10.1000 ;
        RECT 1503.5600 15.0600 1505.1600 15.5400 ;
        RECT 1005.5200 183.7000 1007.1200 184.1800 ;
        RECT 1005.5200 194.5800 1007.1200 195.0600 ;
        RECT 1005.5200 200.0200 1007.1200 200.5000 ;
        RECT 1015.5800 193.0800 1017.1800 193.5600 ;
        RECT 1005.5200 205.4600 1007.1200 205.9400 ;
        RECT 1005.5200 210.9000 1007.1200 211.3800 ;
        RECT 1005.5200 216.3400 1007.1200 216.8200 ;
        RECT 1005.5200 221.7800 1007.1200 222.2600 ;
        RECT 1005.5200 227.2200 1007.1200 227.7000 ;
        RECT 1063.2600 25.9400 1064.8600 26.4200 ;
        RECT 1063.2600 31.3800 1064.8600 31.8600 ;
        RECT 1063.2600 36.8200 1064.8600 37.3000 ;
        RECT 1063.2600 42.2600 1064.8600 42.7400 ;
        RECT 1063.2600 47.7000 1064.8600 48.1800 ;
        RECT 1063.2600 53.1400 1064.8600 53.6200 ;
        RECT 1063.2600 58.5800 1064.8600 59.0600 ;
        RECT 1063.2600 64.0200 1064.8600 64.5000 ;
        RECT 1063.2600 69.4600 1064.8600 69.9400 ;
        RECT 1063.2600 74.9000 1064.8600 75.3800 ;
        RECT 1063.2600 80.3400 1064.8600 80.8200 ;
        RECT 1063.2600 85.7800 1064.8600 86.2600 ;
        RECT 1063.2600 91.2200 1064.8600 91.7000 ;
        RECT 1063.2600 96.6600 1064.8600 97.1400 ;
        RECT 1063.2600 112.9800 1064.8600 113.4600 ;
        RECT 1063.2600 102.1000 1064.8600 102.5800 ;
        RECT 1063.2600 107.5400 1064.8600 108.0200 ;
        RECT 1063.2600 118.4200 1064.8600 118.9000 ;
        RECT 1063.2600 123.8600 1064.8600 124.3400 ;
        RECT 1063.2600 138.6000 1064.8600 140.6600 ;
        RECT 1063.2600 129.3000 1064.8600 129.7800 ;
        RECT 1063.2600 134.7400 1064.8600 135.2200 ;
        RECT 1063.2600 145.6200 1064.8600 146.1000 ;
        RECT 1063.2600 151.0600 1064.8600 151.5400 ;
        RECT 1063.2600 156.5000 1064.8600 156.9800 ;
        RECT 1063.2600 161.9400 1064.8600 162.4200 ;
        RECT 1063.2600 172.8200 1064.8600 173.3000 ;
        RECT 1063.2600 188.7900 1064.8600 190.4900 ;
        RECT 1075.8200 193.0800 1077.4200 193.5600 ;
        RECT 1005.5200 232.6600 1007.1200 233.1400 ;
        RECT 1005.5200 238.1000 1007.1200 238.5800 ;
        RECT 1005.5200 243.5400 1007.1200 244.0200 ;
        RECT 1005.5200 248.9800 1007.1200 249.4600 ;
        RECT 1005.5200 254.4200 1007.1200 254.9000 ;
        RECT 1005.5200 270.7400 1007.1200 271.2200 ;
        RECT 1005.5200 259.8600 1007.1200 260.3400 ;
        RECT 1005.5200 265.3000 1007.1200 265.7800 ;
        RECT 1005.5200 276.1800 1007.1200 276.6600 ;
        RECT 1005.5200 281.6200 1007.1200 282.1000 ;
        RECT 1005.5200 287.0600 1007.1200 287.5400 ;
        RECT 1005.5200 292.5000 1007.1200 292.9800 ;
        RECT 1005.5200 297.9400 1007.1200 298.4200 ;
        RECT 1005.5200 303.3800 1007.1200 303.8600 ;
        RECT 1005.5200 308.8200 1007.1200 309.3000 ;
        RECT 1005.5200 314.2600 1007.1200 314.7400 ;
        RECT 1005.5200 319.7000 1007.1200 320.1800 ;
        RECT 1005.5200 325.1400 1007.1200 325.6200 ;
        RECT 1005.5200 330.5800 1007.1200 331.0600 ;
        RECT 1005.5200 336.0200 1007.1200 336.5000 ;
        RECT 1005.5200 363.2200 1007.1200 363.7000 ;
        RECT 1005.5200 341.4600 1007.1200 341.9400 ;
        RECT 1005.5200 346.9000 1007.1200 347.3800 ;
        RECT 1005.5200 352.3400 1007.1200 352.8200 ;
        RECT 1005.5200 357.7800 1007.1200 358.2600 ;
        RECT 1005.5200 368.6600 1007.1200 369.1400 ;
        RECT 1005.5200 374.1000 1007.1200 374.5800 ;
        RECT 1005.5200 379.5400 1007.1200 380.0200 ;
        RECT 1005.5200 384.9800 1007.1200 385.4600 ;
        RECT 1005.5200 390.4200 1007.1200 390.9000 ;
        RECT 1005.5200 401.3000 1007.1200 401.7800 ;
        RECT 1005.5200 408.1200 1007.1200 410.1000 ;
        RECT 1005.5200 412.1800 1007.1200 412.6600 ;
        RECT 1005.5200 418.1300 1007.1200 420.0300 ;
        RECT 1005.5200 423.0600 1007.1200 423.5400 ;
        RECT 1005.5200 428.5000 1007.1200 428.9800 ;
        RECT 1015.5800 422.7200 1017.1800 423.2000 ;
        RECT 1005.5200 433.9400 1007.1200 434.4200 ;
        RECT 1005.5200 439.3800 1007.1200 439.8600 ;
        RECT 1283.3400 25.9400 1285.0800 26.4200 ;
        RECT 1283.3400 31.3800 1285.0800 31.8600 ;
        RECT 1283.3400 36.8200 1285.0800 37.3000 ;
        RECT 1283.3400 42.2600 1285.0800 42.7400 ;
        RECT 1283.3400 47.7000 1285.0800 48.1800 ;
        RECT 1283.3400 53.1400 1285.0800 53.6200 ;
        RECT 1283.3400 58.5800 1285.0800 59.0600 ;
        RECT 1283.3400 64.0200 1285.0800 64.5000 ;
        RECT 1283.3400 69.4600 1285.0800 69.9400 ;
        RECT 1283.3400 74.9000 1285.0800 75.3800 ;
        RECT 1283.3400 80.3400 1285.0800 80.8200 ;
        RECT 1283.3400 85.7800 1285.0800 86.2600 ;
        RECT 1283.3400 91.2200 1285.0800 91.7000 ;
        RECT 1283.3400 96.6600 1285.0800 97.1400 ;
        RECT 1283.3400 112.9800 1285.0800 113.4600 ;
        RECT 1283.3400 102.1000 1285.0800 102.5800 ;
        RECT 1283.3400 107.5400 1285.0800 108.0200 ;
        RECT 1283.3400 118.4200 1285.0800 118.9000 ;
        RECT 1283.3400 123.8600 1285.0800 124.3400 ;
        RECT 1283.3400 178.6000 1285.0800 180.4600 ;
        RECT 1283.3400 138.3400 1285.0800 140.2000 ;
        RECT 1273.4200 150.1000 1275.0200 150.5800 ;
        RECT 1283.3400 129.3000 1285.0800 129.7800 ;
        RECT 1283.3400 146.9100 1285.0800 148.7700 ;
        RECT 1283.3400 166.4400 1285.0800 168.3000 ;
        RECT 1283.3400 188.6300 1285.0800 190.4900 ;
        RECT 1295.9000 192.8200 1297.5000 193.3000 ;
        RECT 1503.5600 25.9400 1505.1600 26.4200 ;
        RECT 1503.5600 31.3800 1505.1600 31.8600 ;
        RECT 1503.5600 36.8200 1505.1600 37.3000 ;
        RECT 1503.5600 42.2600 1505.1600 42.7400 ;
        RECT 1503.5600 47.7000 1505.1600 48.1800 ;
        RECT 1503.5600 53.1400 1505.1600 53.6200 ;
        RECT 1503.5600 58.5800 1505.1600 59.0600 ;
        RECT 1503.5600 64.0200 1505.1600 64.5000 ;
        RECT 1503.5600 69.4600 1505.1600 69.9400 ;
        RECT 1503.5600 74.9000 1505.1600 75.3800 ;
        RECT 1503.5600 80.3400 1505.1600 80.8200 ;
        RECT 1503.5600 85.7800 1505.1600 86.2600 ;
        RECT 1503.5600 91.2200 1505.1600 91.7000 ;
        RECT 1503.5600 96.6600 1505.1600 97.1400 ;
        RECT 1503.5600 112.9800 1505.1600 113.4600 ;
        RECT 1503.5600 102.1000 1505.1600 102.5800 ;
        RECT 1503.5600 107.5400 1505.1600 108.0200 ;
        RECT 1503.5600 118.4200 1505.1600 118.9000 ;
        RECT 1503.5600 123.8600 1505.1600 124.3400 ;
        RECT 1493.5000 149.8400 1495.1000 150.3200 ;
        RECT 1503.5600 129.3000 1505.1600 129.7800 ;
        RECT 1516.1200 192.8200 1517.7200 193.3000 ;
        RECT 1295.9000 422.4600 1297.5000 422.9400 ;
        RECT 1516.1200 422.4600 1517.7200 422.9400 ;
        RECT 2.0000 444.8200 5.0000 445.3000 ;
        RECT 2.0000 450.2600 5.0000 450.7400 ;
        RECT 2.0000 455.7000 5.0000 456.1800 ;
        RECT 2.0000 461.1400 5.0000 461.6200 ;
        RECT 2.0000 466.5800 5.0000 467.0600 ;
        RECT 2.0000 472.0200 5.0000 472.5000 ;
        RECT 2.0000 477.4600 5.0000 477.9400 ;
        RECT 2.0000 482.9000 5.0000 483.3800 ;
        RECT 2.0000 488.3400 5.0000 488.8200 ;
        RECT 2.0000 493.7800 5.0000 494.2600 ;
        RECT 2.0000 520.9800 5.0000 521.4600 ;
        RECT 2.0000 499.2200 5.0000 499.7000 ;
        RECT 2.0000 504.6600 5.0000 505.1400 ;
        RECT 2.0000 510.1000 5.0000 510.5800 ;
        RECT 2.0000 515.5400 5.0000 516.0200 ;
        RECT 2.0000 526.4200 5.0000 526.9000 ;
        RECT 2.0000 531.8600 5.0000 532.3400 ;
        RECT 2.0000 537.3000 5.0000 537.7800 ;
        RECT 2.0000 542.7400 5.0000 543.2200 ;
        RECT 2.0000 548.1800 5.0000 548.6600 ;
        RECT 2.0000 553.6200 5.0000 554.1000 ;
        RECT 2.0000 559.0600 5.0000 559.5400 ;
        RECT 2.0000 564.5000 5.0000 564.9800 ;
        RECT 2.0000 569.9400 5.0000 570.4200 ;
        RECT 2.0000 575.3800 5.0000 575.8600 ;
        RECT 2.0000 580.8200 5.0000 581.3000 ;
        RECT 2.0000 586.2600 5.0000 586.7400 ;
        RECT 2.0000 591.7000 5.0000 592.1800 ;
        RECT 2.0000 597.1400 5.0000 597.6200 ;
        RECT 2.0000 602.5800 5.0000 603.0600 ;
        RECT 2.0000 608.0200 5.0000 608.5000 ;
        RECT 2.0000 613.4600 5.0000 613.9400 ;
        RECT 2.0000 618.9000 5.0000 619.3800 ;
        RECT 2.0000 624.3400 5.0000 624.8200 ;
        RECT 2.0000 629.7800 5.0000 630.2600 ;
        RECT 2.0000 635.2200 5.0000 635.7000 ;
        RECT 2.0000 640.6600 5.0000 641.1400 ;
        RECT 2.0000 646.1000 5.0000 646.5800 ;
        RECT 2.0000 651.5400 5.0000 652.0200 ;
        RECT 155.5200 640.6600 157.1200 641.1400 ;
        RECT 155.5200 646.1000 157.1200 646.5800 ;
        RECT 155.5200 651.5400 157.1200 652.0200 ;
        RECT 2.0000 656.9800 5.0000 657.4600 ;
        RECT 2.0000 662.4200 5.0000 662.9000 ;
        RECT 2.0000 667.8600 5.0000 668.3400 ;
        RECT 2.0000 673.3000 5.0000 673.7800 ;
        RECT 2.0000 678.7400 5.0000 679.2200 ;
        RECT 2.0000 684.1800 5.0000 684.6600 ;
        RECT 2.0000 689.6200 5.0000 690.1000 ;
        RECT 2.0000 695.0600 5.0000 695.5400 ;
        RECT 2.0000 700.5000 5.0000 700.9800 ;
        RECT 2.0000 705.9400 5.0000 706.4200 ;
        RECT 2.0000 711.3800 5.0000 711.8600 ;
        RECT 2.0000 716.8200 5.0000 717.3000 ;
        RECT 2.0000 722.2600 5.0000 722.7400 ;
        RECT 2.0000 727.7000 5.0000 728.1800 ;
        RECT 2.0000 733.1400 5.0000 733.6200 ;
        RECT 2.0000 738.5800 5.0000 739.0600 ;
        RECT 2.0000 744.0200 5.0000 744.5000 ;
        RECT 2.0000 749.4600 5.0000 749.9400 ;
        RECT 2.0000 754.9000 5.0000 755.3800 ;
        RECT 155.5200 656.9800 157.1200 657.4600 ;
        RECT 155.5200 662.4200 157.1200 662.9000 ;
        RECT 155.5200 667.8600 157.1200 668.3400 ;
        RECT 155.5200 673.3000 157.1200 673.7800 ;
        RECT 155.5200 678.7400 157.1200 679.2200 ;
        RECT 155.5200 684.1800 157.1200 684.6600 ;
        RECT 155.5200 689.6200 157.1200 690.1000 ;
        RECT 155.5200 695.0600 157.1200 695.5400 ;
        RECT 155.5200 700.5000 157.1200 700.9800 ;
        RECT 155.5200 705.9400 157.1200 706.4200 ;
        RECT 155.5200 711.3800 157.1200 711.8600 ;
        RECT 155.5200 716.8200 157.1200 717.3000 ;
        RECT 155.5200 722.2600 157.1200 722.7400 ;
        RECT 155.5200 727.7000 157.1200 728.1800 ;
        RECT 155.5200 733.1400 157.1200 733.6200 ;
        RECT 155.5200 738.5800 157.1200 739.0600 ;
        RECT 155.5200 744.0200 157.1200 744.5000 ;
        RECT 155.5200 749.4600 157.1200 749.9400 ;
        RECT 155.5200 754.9000 157.1200 755.3800 ;
        RECT 2.0000 771.2200 5.0000 771.7000 ;
        RECT 2.0000 760.3400 5.0000 760.8200 ;
        RECT 2.0000 765.7800 5.0000 766.2600 ;
        RECT 2.0000 776.6600 5.0000 777.1400 ;
        RECT 2.0000 782.1000 5.0000 782.5800 ;
        RECT 2.0000 787.5400 5.0000 788.0200 ;
        RECT 2.0000 792.9800 5.0000 793.4600 ;
        RECT 2.0000 798.4200 5.0000 798.9000 ;
        RECT 2.0000 803.8600 5.0000 804.3400 ;
        RECT 2.0000 809.3000 5.0000 809.7800 ;
        RECT 2.0000 814.7400 5.0000 815.2200 ;
        RECT 2.0000 820.1800 5.0000 820.6600 ;
        RECT 2.0000 825.6200 5.0000 826.1000 ;
        RECT 2.0000 831.0600 5.0000 831.5400 ;
        RECT 2.0000 836.5000 5.0000 836.9800 ;
        RECT 2.0000 841.9400 5.0000 842.4200 ;
        RECT 2.0000 847.3800 5.0000 847.8600 ;
        RECT 2.0000 852.8200 5.0000 853.3000 ;
        RECT 2.0000 858.2600 5.0000 858.7400 ;
        RECT 155.5200 771.2200 157.1200 771.7000 ;
        RECT 155.5200 760.3400 157.1200 760.8200 ;
        RECT 155.5200 765.7800 157.1200 766.2600 ;
        RECT 155.5200 776.6600 157.1200 777.1400 ;
        RECT 155.5200 782.1000 157.1200 782.5800 ;
        RECT 155.5200 787.5400 157.1200 788.0200 ;
        RECT 155.5200 792.9800 157.1200 793.4600 ;
        RECT 155.5200 798.4200 157.1200 798.9000 ;
        RECT 155.5200 803.8600 157.1200 804.3400 ;
        RECT 155.5200 809.3000 157.1200 809.7800 ;
        RECT 155.5200 814.7400 157.1200 815.2200 ;
        RECT 155.5200 820.1800 157.1200 820.6600 ;
        RECT 155.5200 825.6200 157.1200 826.1000 ;
        RECT 155.5200 831.0600 157.1200 831.5400 ;
        RECT 155.5200 836.5000 157.1200 836.9800 ;
        RECT 155.5200 841.9400 157.1200 842.4200 ;
        RECT 155.5200 847.3800 157.1200 847.8600 ;
        RECT 155.5200 852.8200 157.1200 853.3000 ;
        RECT 155.5200 858.2600 157.1200 858.7400 ;
        RECT 505.5200 444.8200 507.1200 445.3000 ;
        RECT 505.5200 450.2600 507.1200 450.7400 ;
        RECT 505.5200 455.7000 507.1200 456.1800 ;
        RECT 505.5200 461.1400 507.1200 461.6200 ;
        RECT 505.5200 466.5800 507.1200 467.0600 ;
        RECT 505.5200 472.0200 507.1200 472.5000 ;
        RECT 505.5200 477.4600 507.1200 477.9400 ;
        RECT 505.5200 482.9000 507.1200 483.3800 ;
        RECT 505.5200 488.3400 507.1200 488.8200 ;
        RECT 505.5200 493.7800 507.1200 494.2600 ;
        RECT 505.5200 520.9800 507.1200 521.4600 ;
        RECT 505.5200 499.2200 507.1200 499.7000 ;
        RECT 505.5200 504.6600 507.1200 505.1400 ;
        RECT 505.5200 510.1000 507.1200 510.5800 ;
        RECT 505.5200 515.5400 507.1200 516.0200 ;
        RECT 505.5200 526.4200 507.1200 526.9000 ;
        RECT 505.5200 531.8600 507.1200 532.3400 ;
        RECT 505.5200 537.3000 507.1200 537.7800 ;
        RECT 505.5200 542.7400 507.1200 543.2200 ;
        RECT 505.5200 548.1800 507.1200 548.6600 ;
        RECT 505.5200 553.6200 507.1200 554.1000 ;
        RECT 505.5200 559.0600 507.1200 559.5400 ;
        RECT 505.5200 564.5000 507.1200 564.9800 ;
        RECT 505.5200 569.9400 507.1200 570.4200 ;
        RECT 505.5200 575.3800 507.1200 575.8600 ;
        RECT 505.5200 580.8200 507.1200 581.3000 ;
        RECT 505.5200 586.2600 507.1200 586.7400 ;
        RECT 505.5200 591.7000 507.1200 592.1800 ;
        RECT 505.5200 597.1400 507.1200 597.6200 ;
        RECT 505.5200 602.5800 507.1200 603.0600 ;
        RECT 505.5200 608.0200 507.1200 608.5000 ;
        RECT 505.5200 613.4600 507.1200 613.9400 ;
        RECT 505.5200 618.9000 507.1200 619.3800 ;
        RECT 505.5200 624.3400 507.1200 624.8200 ;
        RECT 505.5200 629.7800 507.1200 630.2600 ;
        RECT 663.1200 444.8200 664.7200 445.3000 ;
        RECT 663.1200 450.2600 664.7200 450.7400 ;
        RECT 663.1200 466.5800 664.7200 467.0600 ;
        RECT 663.1200 461.1400 664.7200 461.6200 ;
        RECT 663.1200 455.7000 664.7200 456.1800 ;
        RECT 663.1200 472.0200 664.7200 472.5000 ;
        RECT 663.1200 477.4600 664.7200 477.9400 ;
        RECT 663.1200 482.9000 664.7200 483.3800 ;
        RECT 663.1200 488.3400 664.7200 488.8200 ;
        RECT 663.1200 493.7800 664.7200 494.2600 ;
        RECT 663.1200 520.9800 664.7200 521.4600 ;
        RECT 663.1200 504.6600 664.7200 505.1400 ;
        RECT 663.1200 499.2200 664.7200 499.7000 ;
        RECT 663.1200 510.1000 664.7200 510.5800 ;
        RECT 663.1200 515.5400 664.7200 516.0200 ;
        RECT 663.1200 526.4200 664.7200 526.9000 ;
        RECT 663.1200 531.8600 664.7200 532.3400 ;
        RECT 663.1200 537.3000 664.7200 537.7800 ;
        RECT 663.1200 542.7400 664.7200 543.2200 ;
        RECT 663.1200 548.1800 664.7200 548.6600 ;
        RECT 663.1200 553.6200 664.7200 554.1000 ;
        RECT 663.1200 559.0600 664.7200 559.5400 ;
        RECT 663.1200 564.5000 664.7200 564.9800 ;
        RECT 663.1200 569.9400 664.7200 570.4200 ;
        RECT 663.1200 575.3800 664.7200 575.8600 ;
        RECT 663.1200 580.8200 664.7200 581.3000 ;
        RECT 663.1200 586.2600 664.7200 586.7400 ;
        RECT 663.1200 591.7000 664.7200 592.1800 ;
        RECT 663.1200 597.1400 664.7200 597.6200 ;
        RECT 663.1200 602.5800 664.7200 603.0600 ;
        RECT 663.1200 608.0200 664.7200 608.5000 ;
        RECT 663.1200 613.4600 664.7200 613.9400 ;
        RECT 663.1200 618.9000 664.7200 619.3800 ;
        RECT 663.1200 624.3400 664.7200 624.8200 ;
        RECT 663.1200 629.7800 664.7200 630.2600 ;
        RECT 2.0000 874.5800 5.0000 875.0600 ;
        RECT 2.0000 867.7800 5.0000 869.6200 ;
        RECT 2.0000 863.7000 5.0000 864.1800 ;
        RECT 2.0000 880.0200 5.0000 880.5000 ;
        RECT 2.0000 885.4600 5.0000 885.9400 ;
        RECT 2.0000 890.9000 5.0000 891.3800 ;
        RECT 2.0000 896.3400 5.0000 896.8200 ;
        RECT 2.0000 901.7800 5.0000 902.2600 ;
        RECT 2.0000 907.2200 5.0000 907.7000 ;
        RECT 2.0000 912.6600 5.0000 913.1400 ;
        RECT 2.0000 928.9800 5.0000 929.4600 ;
        RECT 2.0000 918.1000 5.0000 918.5800 ;
        RECT 2.0000 923.5400 5.0000 924.0200 ;
        RECT 2.0000 934.4200 5.0000 934.9000 ;
        RECT 2.0000 939.8600 5.0000 940.3400 ;
        RECT 2.0000 945.3000 5.0000 945.7800 ;
        RECT 2.0000 950.7400 5.0000 951.2200 ;
        RECT 2.0000 956.1800 5.0000 956.6600 ;
        RECT 2.0000 961.6200 5.0000 962.1000 ;
        RECT 2.0000 967.0600 5.0000 967.5400 ;
        RECT 155.5200 874.5800 157.1200 875.0600 ;
        RECT 155.5200 867.7800 157.1200 869.6200 ;
        RECT 155.5200 863.7000 157.1200 864.1800 ;
        RECT 155.5200 880.0200 157.1200 880.5000 ;
        RECT 155.5200 885.4600 157.1200 885.9400 ;
        RECT 155.5200 890.9000 157.1200 891.3800 ;
        RECT 155.5200 896.3400 157.1200 896.8200 ;
        RECT 155.5200 901.7800 157.1200 902.2600 ;
        RECT 155.5200 907.2200 157.1200 907.7000 ;
        RECT 155.5200 912.6600 157.1200 913.1400 ;
        RECT 155.5200 928.9800 157.1200 929.4600 ;
        RECT 155.5200 918.1000 157.1200 918.5800 ;
        RECT 155.5200 923.5400 157.1200 924.0200 ;
        RECT 155.5200 934.4200 157.1200 934.9000 ;
        RECT 155.5200 939.8600 157.1200 940.3400 ;
        RECT 155.5200 945.3000 157.1200 945.7800 ;
        RECT 155.5200 950.7400 157.1200 951.2200 ;
        RECT 155.5200 956.1800 157.1200 956.6600 ;
        RECT 155.5200 961.6200 157.1200 962.1000 ;
        RECT 155.5200 967.0600 157.1200 967.5400 ;
        RECT 2.0000 1021.4600 5.0000 1021.9400 ;
        RECT 2.0000 972.5000 5.0000 972.9800 ;
        RECT 2.0000 977.9400 5.0000 978.4200 ;
        RECT 2.0000 983.3800 5.0000 983.8600 ;
        RECT 2.0000 988.8200 5.0000 989.3000 ;
        RECT 2.0000 994.2600 5.0000 994.7400 ;
        RECT 2.0000 999.7000 5.0000 1000.1800 ;
        RECT 2.0000 1005.1400 5.0000 1005.6200 ;
        RECT 2.0000 1010.5800 5.0000 1011.0600 ;
        RECT 2.0000 1016.0200 5.0000 1016.5000 ;
        RECT 2.0000 1026.9000 5.0000 1027.3800 ;
        RECT 2.0000 1032.3400 5.0000 1032.8200 ;
        RECT 2.0000 1037.7800 5.0000 1038.2600 ;
        RECT 2.0000 1043.2200 5.0000 1043.7000 ;
        RECT 2.0000 1048.6600 5.0000 1049.1400 ;
        RECT 2.0000 1054.1000 5.0000 1054.5800 ;
        RECT 2.0000 1059.5400 5.0000 1060.0200 ;
        RECT 2.0000 1064.9800 5.0000 1065.4600 ;
        RECT 2.0000 1070.4200 5.0000 1070.9000 ;
        RECT 155.5200 1021.4600 157.1200 1021.9400 ;
        RECT 155.5200 972.5000 157.1200 972.9800 ;
        RECT 155.5200 977.9400 157.1200 978.4200 ;
        RECT 155.5200 983.3800 157.1200 983.8600 ;
        RECT 155.5200 988.8200 157.1200 989.3000 ;
        RECT 155.5200 994.2600 157.1200 994.7400 ;
        RECT 155.5200 999.7000 157.1200 1000.1800 ;
        RECT 155.5200 1005.1400 157.1200 1005.6200 ;
        RECT 155.5200 1010.5800 157.1200 1011.0600 ;
        RECT 155.5200 1016.0200 157.1200 1016.5000 ;
        RECT 155.5200 1026.9000 157.1200 1027.3800 ;
        RECT 155.5200 1032.3400 157.1200 1032.8200 ;
        RECT 155.5200 1037.7800 157.1200 1038.2600 ;
        RECT 155.5200 1043.2200 157.1200 1043.7000 ;
        RECT 155.5200 1048.6600 157.1200 1049.1400 ;
        RECT 155.5200 1054.1000 157.1200 1054.5800 ;
        RECT 155.5200 1059.5400 157.1200 1060.0200 ;
        RECT 155.5200 1064.9800 157.1200 1065.4600 ;
        RECT 155.5200 1070.4200 157.1200 1070.9000 ;
        RECT 2.0000 1179.2200 5.0000 1179.7000 ;
        RECT 155.5200 1179.2200 157.1200 1179.7000 ;
        RECT 2.0000 1075.8600 5.0000 1076.3400 ;
        RECT 2.0000 1081.3000 5.0000 1081.7800 ;
        RECT 2.0000 1086.7400 5.0000 1087.2200 ;
        RECT 2.0000 1092.1800 5.0000 1092.6600 ;
        RECT 2.0000 1103.0600 5.0000 1103.5400 ;
        RECT 2.0000 1108.5000 5.0000 1108.9800 ;
        RECT 2.0000 1113.9400 5.0000 1114.4200 ;
        RECT 2.0000 1119.3800 5.0000 1119.8600 ;
        RECT 2.0000 1124.8200 5.0000 1125.3000 ;
        RECT 2.0000 1130.2600 5.0000 1130.7400 ;
        RECT 2.0000 1135.7000 5.0000 1136.1800 ;
        RECT 2.0000 1141.1400 5.0000 1141.6200 ;
        RECT 2.0000 1146.5800 5.0000 1147.0600 ;
        RECT 2.0000 1152.0200 5.0000 1152.5000 ;
        RECT 2.0000 1157.4600 5.0000 1157.9400 ;
        RECT 2.0000 1162.9000 5.0000 1163.3800 ;
        RECT 2.0000 1168.3400 5.0000 1168.8200 ;
        RECT 2.0000 1173.7800 5.0000 1174.2600 ;
        RECT 155.5200 1075.8600 157.1200 1076.3400 ;
        RECT 155.5200 1081.3000 157.1200 1081.7800 ;
        RECT 155.5200 1086.7400 157.1200 1087.2200 ;
        RECT 155.5200 1092.1800 157.1200 1092.6600 ;
        RECT 155.5200 1103.0600 157.1200 1103.5400 ;
        RECT 155.5200 1108.5000 157.1200 1108.9800 ;
        RECT 155.5200 1113.9400 157.1200 1114.4200 ;
        RECT 155.5200 1119.3800 157.1200 1119.8600 ;
        RECT 155.5200 1124.8200 157.1200 1125.3000 ;
        RECT 155.5200 1130.2600 157.1200 1130.7400 ;
        RECT 155.5200 1135.7000 157.1200 1136.1800 ;
        RECT 155.5200 1141.1400 157.1200 1141.6200 ;
        RECT 155.5200 1146.5800 157.1200 1147.0600 ;
        RECT 155.5200 1152.0200 157.1200 1152.5000 ;
        RECT 155.5200 1157.4600 157.1200 1157.9400 ;
        RECT 155.5200 1162.9000 157.1200 1163.3800 ;
        RECT 155.5200 1168.3400 157.1200 1168.8200 ;
        RECT 155.5200 1173.7800 157.1200 1174.2600 ;
        RECT 2.0000 1184.6600 5.0000 1185.1400 ;
        RECT 2.0000 1190.1000 5.0000 1190.5800 ;
        RECT 2.0000 1195.5400 5.0000 1196.0200 ;
        RECT 2.0000 1200.9800 5.0000 1201.4600 ;
        RECT 2.0000 1206.4200 5.0000 1206.9000 ;
        RECT 2.0000 1211.8600 5.0000 1212.3400 ;
        RECT 2.0000 1217.3000 5.0000 1217.7800 ;
        RECT 2.0000 1222.7400 5.0000 1223.2200 ;
        RECT 2.0000 1228.1800 5.0000 1228.6600 ;
        RECT 2.0000 1233.6200 5.0000 1234.1000 ;
        RECT 2.0000 1239.0600 5.0000 1239.5400 ;
        RECT 2.0000 1244.5000 5.0000 1244.9800 ;
        RECT 2.0000 1249.9400 5.0000 1250.4200 ;
        RECT 2.0000 1255.3800 5.0000 1255.8600 ;
        RECT 2.0000 1260.8200 5.0000 1261.3000 ;
        RECT 2.0000 1266.2600 5.0000 1266.7400 ;
        RECT 2.0000 1271.7000 5.0000 1272.1800 ;
        RECT 2.0000 1277.1400 5.0000 1277.6200 ;
        RECT 2.0000 1282.5800 5.0000 1283.0600 ;
        RECT 155.5200 1184.6600 157.1200 1185.1400 ;
        RECT 155.5200 1190.1000 157.1200 1190.5800 ;
        RECT 155.5200 1195.5400 157.1200 1196.0200 ;
        RECT 155.5200 1200.9800 157.1200 1201.4600 ;
        RECT 155.5200 1206.4200 157.1200 1206.9000 ;
        RECT 155.5200 1211.8600 157.1200 1212.3400 ;
        RECT 155.5200 1217.3000 157.1200 1217.7800 ;
        RECT 155.5200 1222.7400 157.1200 1223.2200 ;
        RECT 155.5200 1228.1800 157.1200 1228.6600 ;
        RECT 155.5200 1233.6200 157.1200 1234.1000 ;
        RECT 155.5200 1239.0600 157.1200 1239.5400 ;
        RECT 155.5200 1244.5000 157.1200 1244.9800 ;
        RECT 155.5200 1249.9400 157.1200 1250.4200 ;
        RECT 155.5200 1255.3800 157.1200 1255.8600 ;
        RECT 155.5200 1260.8200 157.1200 1261.3000 ;
        RECT 155.5200 1266.2600 157.1200 1266.7400 ;
        RECT 155.5200 1271.7000 157.1200 1272.1800 ;
        RECT 155.5200 1277.1400 157.1200 1277.6200 ;
        RECT 155.5200 1282.5800 157.1200 1283.0600 ;
        RECT 1005.5200 444.8200 1007.1200 445.3000 ;
        RECT 1005.5200 450.2600 1007.1200 450.7400 ;
        RECT 1005.5200 455.7000 1007.1200 456.1800 ;
        RECT 1005.5200 461.1400 1007.1200 461.6200 ;
        RECT 1005.5200 466.5800 1007.1200 467.0600 ;
        RECT 1005.5200 472.0200 1007.1200 472.5000 ;
        RECT 1005.5200 477.4600 1007.1200 477.9400 ;
        RECT 1005.5200 482.9000 1007.1200 483.3800 ;
        RECT 1005.5200 488.3400 1007.1200 488.8200 ;
        RECT 1005.5200 493.7800 1007.1200 494.2600 ;
        RECT 1005.5200 520.9800 1007.1200 521.4600 ;
        RECT 1005.5200 499.2200 1007.1200 499.7000 ;
        RECT 1005.5200 504.6600 1007.1200 505.1400 ;
        RECT 1005.5200 510.1000 1007.1200 510.5800 ;
        RECT 1005.5200 515.5400 1007.1200 516.0200 ;
        RECT 1005.5200 526.4200 1007.1200 526.9000 ;
        RECT 1005.5200 531.8600 1007.1200 532.3400 ;
        RECT 1005.5200 537.3000 1007.1200 537.7800 ;
        RECT 1005.5200 542.7400 1007.1200 543.2200 ;
        RECT 1005.5200 548.1800 1007.1200 548.6600 ;
        RECT 1005.5200 553.6200 1007.1200 554.1000 ;
        RECT 1005.5200 559.0600 1007.1200 559.5400 ;
        RECT 1005.5200 564.5000 1007.1200 564.9800 ;
        RECT 1005.5200 569.9400 1007.1200 570.4200 ;
        RECT 1005.5200 575.3800 1007.1200 575.8600 ;
        RECT 1005.5200 580.8200 1007.1200 581.3000 ;
        RECT 1005.5200 586.2600 1007.1200 586.7400 ;
        RECT 1005.5200 591.7000 1007.1200 592.1800 ;
        RECT 1005.5200 597.1400 1007.1200 597.6200 ;
        RECT 963.1200 640.6600 964.7200 641.1400 ;
        RECT 963.1200 646.1000 964.7200 646.5800 ;
        RECT 963.1200 651.5400 964.7200 652.0200 ;
        RECT 1005.5200 602.5800 1007.1200 603.0600 ;
        RECT 1005.5200 608.0200 1007.1200 608.5000 ;
        RECT 1005.5200 613.4600 1007.1200 613.9400 ;
        RECT 1005.5200 618.9000 1007.1200 619.3800 ;
        RECT 1005.5200 624.3400 1007.1200 624.8200 ;
        RECT 1005.5200 629.7800 1007.1200 630.2600 ;
        RECT 1005.5200 634.7100 1007.1200 635.1900 ;
        RECT 1005.5200 640.6600 1007.1200 641.1400 ;
        RECT 1005.5200 644.8000 1007.1200 645.2800 ;
        RECT 1005.5200 651.5400 1007.1200 652.0200 ;
        RECT 1015.5800 652.3600 1017.1800 652.8400 ;
        RECT 1063.2600 625.1300 1064.8600 627.6800 ;
        RECT 1063.2600 648.0700 1064.8600 649.7700 ;
        RECT 1075.8200 652.3600 1077.4200 652.8400 ;
        RECT 963.1200 656.9800 964.7200 657.4600 ;
        RECT 963.1200 662.4200 964.7200 662.9000 ;
        RECT 963.1200 667.8600 964.7200 668.3400 ;
        RECT 963.1200 673.3000 964.7200 673.7800 ;
        RECT 963.1200 678.7400 964.7200 679.2200 ;
        RECT 963.1200 684.1800 964.7200 684.6600 ;
        RECT 963.1200 689.6200 964.7200 690.1000 ;
        RECT 963.1200 695.0600 964.7200 695.5400 ;
        RECT 963.1200 700.5000 964.7200 700.9800 ;
        RECT 1005.5200 656.9800 1007.1200 657.4600 ;
        RECT 1005.5200 662.4200 1007.1200 662.9000 ;
        RECT 1005.5200 667.8600 1007.1200 668.3400 ;
        RECT 1005.5200 673.3000 1007.1200 673.7800 ;
        RECT 1005.5200 678.7400 1007.1200 679.2200 ;
        RECT 1005.5200 684.1800 1007.1200 684.6600 ;
        RECT 1005.5200 689.6200 1007.1200 690.1000 ;
        RECT 1005.5200 695.0600 1007.1200 695.5400 ;
        RECT 1005.5200 700.5000 1007.1200 700.9800 ;
        RECT 963.1200 705.9400 964.7200 706.4200 ;
        RECT 963.1200 711.3800 964.7200 711.8600 ;
        RECT 963.1200 716.8200 964.7200 717.3000 ;
        RECT 963.1200 722.2600 964.7200 722.7400 ;
        RECT 963.1200 727.7000 964.7200 728.1800 ;
        RECT 963.1200 744.0200 964.7200 744.5000 ;
        RECT 963.1200 738.5800 964.7200 739.0600 ;
        RECT 963.1200 733.1400 964.7200 733.6200 ;
        RECT 963.1200 749.4600 964.7200 749.9400 ;
        RECT 1005.5200 705.9400 1007.1200 706.4200 ;
        RECT 1005.5200 711.3800 1007.1200 711.8600 ;
        RECT 1005.5200 716.8200 1007.1200 717.3000 ;
        RECT 1005.5200 722.2600 1007.1200 722.7400 ;
        RECT 1005.5200 727.7000 1007.1200 728.1800 ;
        RECT 1005.5200 744.0200 1007.1200 744.5000 ;
        RECT 1005.5200 738.5800 1007.1200 739.0600 ;
        RECT 1005.5200 733.1400 1007.1200 733.6200 ;
        RECT 1005.5200 749.4600 1007.1200 749.9400 ;
        RECT 1283.3400 624.7700 1285.0800 627.6800 ;
        RECT 1283.3400 637.8800 1285.0800 639.7400 ;
        RECT 1283.3400 647.9100 1285.0800 649.7700 ;
        RECT 1295.9000 652.1000 1297.5000 652.5800 ;
        RECT 1516.1200 652.1000 1517.7200 652.5800 ;
        RECT 1015.5800 882.0000 1017.1800 882.4800 ;
        RECT 1015.5800 1111.6400 1017.1800 1112.1200 ;
        RECT 1063.2600 1084.4100 1064.8600 1086.9600 ;
        RECT 1063.2600 1107.3500 1064.8600 1109.0500 ;
        RECT 1075.8200 1111.6400 1077.4200 1112.1200 ;
        RECT 1295.9000 881.7400 1297.5000 882.2200 ;
        RECT 1516.1200 881.7400 1517.7200 882.2200 ;
        RECT 1283.3400 1097.1600 1285.0800 1099.0200 ;
        RECT 1283.3400 1084.0500 1285.0800 1086.9600 ;
        RECT 1283.3400 1107.1900 1285.0800 1109.0500 ;
        RECT 1295.9000 1111.3800 1297.5000 1111.8600 ;
        RECT 1516.1200 1111.3800 1517.7200 1111.8600 ;
        RECT 1944.0000 20.5000 1945.6000 20.9800 ;
        RECT 1723.7800 20.5000 1725.3800 20.9800 ;
        RECT 2384.4400 20.5000 2386.0400 20.9800 ;
        RECT 2164.2200 20.5000 2165.8200 20.9800 ;
        RECT 2444.5800 20.5000 2446.1800 20.9800 ;
        RECT 2495.5200 20.5000 2497.1200 20.9800 ;
        RECT 1723.7800 9.6200 1725.3800 10.1000 ;
        RECT 1723.7800 15.0600 1725.3800 15.5400 ;
        RECT 1944.0000 9.6200 1945.6000 10.1000 ;
        RECT 1944.0000 15.0600 1945.6000 15.5400 ;
        RECT 2164.2200 9.6200 2165.8200 10.1000 ;
        RECT 2164.2200 15.0600 2165.8200 15.5400 ;
        RECT 2384.4400 9.6200 2386.0400 10.1000 ;
        RECT 2384.4400 15.0600 2386.0400 15.5400 ;
        RECT 2444.5800 9.6200 2446.1800 10.1000 ;
        RECT 2444.5800 15.0600 2446.1800 15.5400 ;
        RECT 2495.5200 9.6200 2497.1200 10.1000 ;
        RECT 2495.5200 15.0600 2497.1200 15.5400 ;
        RECT 1723.7800 25.9400 1725.3800 26.4200 ;
        RECT 1723.7800 31.3800 1725.3800 31.8600 ;
        RECT 1723.7800 36.8200 1725.3800 37.3000 ;
        RECT 1723.7800 42.2600 1725.3800 42.7400 ;
        RECT 1723.7800 47.7000 1725.3800 48.1800 ;
        RECT 1723.7800 53.1400 1725.3800 53.6200 ;
        RECT 1723.7800 58.5800 1725.3800 59.0600 ;
        RECT 1723.7800 64.0200 1725.3800 64.5000 ;
        RECT 1723.7800 69.4600 1725.3800 69.9400 ;
        RECT 1723.7800 74.9000 1725.3800 75.3800 ;
        RECT 1723.7800 80.3400 1725.3800 80.8200 ;
        RECT 1723.7800 85.7800 1725.3800 86.2600 ;
        RECT 1723.7800 91.2200 1725.3800 91.7000 ;
        RECT 1723.7800 96.6600 1725.3800 97.1400 ;
        RECT 1723.7800 112.9800 1725.3800 113.4600 ;
        RECT 1723.7800 102.1000 1725.3800 102.5800 ;
        RECT 1723.7800 107.5400 1725.3800 108.0200 ;
        RECT 1723.7800 118.4200 1725.3800 118.9000 ;
        RECT 1723.7800 123.8600 1725.3800 124.3400 ;
        RECT 1723.7800 129.3000 1725.3800 129.7800 ;
        RECT 1713.7200 149.8400 1715.3200 150.3200 ;
        RECT 1736.3400 192.8200 1737.9400 193.3000 ;
        RECT 1944.0000 25.9400 1945.6000 26.4200 ;
        RECT 1944.0000 31.3800 1945.6000 31.8600 ;
        RECT 1944.0000 36.8200 1945.6000 37.3000 ;
        RECT 1944.0000 42.2600 1945.6000 42.7400 ;
        RECT 1944.0000 47.7000 1945.6000 48.1800 ;
        RECT 1944.0000 53.1400 1945.6000 53.6200 ;
        RECT 1944.0000 58.5800 1945.6000 59.0600 ;
        RECT 1944.0000 64.0200 1945.6000 64.5000 ;
        RECT 1944.0000 69.4600 1945.6000 69.9400 ;
        RECT 1944.0000 74.9000 1945.6000 75.3800 ;
        RECT 1944.0000 80.3400 1945.6000 80.8200 ;
        RECT 1944.0000 85.7800 1945.6000 86.2600 ;
        RECT 1944.0000 91.2200 1945.6000 91.7000 ;
        RECT 1944.0000 96.6600 1945.6000 97.1400 ;
        RECT 1944.0000 112.9800 1945.6000 113.4600 ;
        RECT 1944.0000 102.1000 1945.6000 102.5800 ;
        RECT 1944.0000 107.5400 1945.6000 108.0200 ;
        RECT 1944.0000 118.4200 1945.6000 118.9000 ;
        RECT 1944.0000 123.8600 1945.6000 124.3400 ;
        RECT 1933.9400 149.8400 1935.5400 150.3200 ;
        RECT 1944.0000 129.3000 1945.6000 129.7800 ;
        RECT 1956.5600 192.8200 1958.1600 193.3000 ;
        RECT 1736.3400 422.4600 1737.9400 422.9400 ;
        RECT 2164.2200 25.9400 2165.8200 26.4200 ;
        RECT 2164.2200 31.3800 2165.8200 31.8600 ;
        RECT 2164.2200 36.8200 2165.8200 37.3000 ;
        RECT 2164.2200 42.2600 2165.8200 42.7400 ;
        RECT 2164.2200 47.7000 2165.8200 48.1800 ;
        RECT 2164.2200 53.1400 2165.8200 53.6200 ;
        RECT 2164.2200 58.5800 2165.8200 59.0600 ;
        RECT 2164.2200 64.0200 2165.8200 64.5000 ;
        RECT 2164.2200 69.4600 2165.8200 69.9400 ;
        RECT 2164.2200 74.9000 2165.8200 75.3800 ;
        RECT 2164.2200 80.3400 2165.8200 80.8200 ;
        RECT 2164.2200 85.7800 2165.8200 86.2600 ;
        RECT 2164.2200 91.2200 2165.8200 91.7000 ;
        RECT 2164.2200 96.6600 2165.8200 97.1400 ;
        RECT 2164.2200 112.9800 2165.8200 113.4600 ;
        RECT 2164.2200 102.1000 2165.8200 102.5800 ;
        RECT 2164.2200 107.5400 2165.8200 108.0200 ;
        RECT 2164.2200 118.4200 2165.8200 118.9000 ;
        RECT 2164.2200 123.8600 2165.8200 124.3400 ;
        RECT 2154.1600 149.8400 2155.7600 150.3200 ;
        RECT 2164.2200 129.3000 2165.8200 129.7800 ;
        RECT 2176.7800 192.8200 2178.3800 193.3000 ;
        RECT 2384.4400 25.9400 2386.0400 26.4200 ;
        RECT 2384.4400 31.3800 2386.0400 31.8600 ;
        RECT 2384.4400 36.8200 2386.0400 37.3000 ;
        RECT 2384.4400 42.2600 2386.0400 42.7400 ;
        RECT 2384.4400 47.7000 2386.0400 48.1800 ;
        RECT 2384.4400 53.1400 2386.0400 53.6200 ;
        RECT 2384.4400 58.5800 2386.0400 59.0600 ;
        RECT 2384.4400 64.0200 2386.0400 64.5000 ;
        RECT 2384.4400 69.4600 2386.0400 69.9400 ;
        RECT 2384.4400 74.9000 2386.0400 75.3800 ;
        RECT 2384.4400 80.3400 2386.0400 80.8200 ;
        RECT 2384.4400 85.7800 2386.0400 86.2600 ;
        RECT 2384.4400 91.2200 2386.0400 91.7000 ;
        RECT 2384.4400 96.6600 2386.0400 97.1400 ;
        RECT 2384.4400 112.9800 2386.0400 113.4600 ;
        RECT 2384.4400 102.1000 2386.0400 102.5800 ;
        RECT 2384.4400 107.5400 2386.0400 108.0200 ;
        RECT 2384.4400 118.4200 2386.0400 118.9000 ;
        RECT 2384.4400 123.8600 2386.0400 124.3400 ;
        RECT 2444.5800 25.9400 2446.1800 26.4200 ;
        RECT 2444.5800 31.3800 2446.1800 31.8600 ;
        RECT 2444.5800 36.8200 2446.1800 37.3000 ;
        RECT 2444.5800 42.2600 2446.1800 42.7400 ;
        RECT 2444.5800 47.7000 2446.1800 48.1800 ;
        RECT 2444.5800 53.1400 2446.1800 53.6200 ;
        RECT 2444.5800 58.5800 2446.1800 59.0600 ;
        RECT 2444.5800 64.0200 2446.1800 64.5000 ;
        RECT 2444.5800 69.4600 2446.1800 69.9400 ;
        RECT 2495.5200 25.9400 2497.1200 26.4200 ;
        RECT 2495.5200 31.3800 2497.1200 31.8600 ;
        RECT 2495.5200 36.8200 2497.1200 37.3000 ;
        RECT 2495.5200 42.2600 2497.1200 42.7400 ;
        RECT 2495.5200 47.7000 2497.1200 48.1800 ;
        RECT 2495.5200 53.1400 2497.1200 53.6200 ;
        RECT 2495.5200 58.5800 2497.1200 59.0600 ;
        RECT 2495.5200 64.0200 2497.1200 64.5000 ;
        RECT 2495.5200 69.4600 2497.1200 69.9400 ;
        RECT 2444.5800 74.9000 2446.1800 75.3800 ;
        RECT 2444.5800 80.3400 2446.1800 80.8200 ;
        RECT 2444.5800 85.7800 2446.1800 86.2600 ;
        RECT 2444.5800 91.2200 2446.1800 91.7000 ;
        RECT 2444.5800 96.6600 2446.1800 97.1400 ;
        RECT 2444.5800 112.9800 2446.1800 113.4600 ;
        RECT 2444.5800 102.1000 2446.1800 102.5800 ;
        RECT 2444.5800 107.5400 2446.1800 108.0200 ;
        RECT 2444.5800 118.4200 2446.1800 118.9000 ;
        RECT 2444.5800 123.8600 2446.1800 124.3400 ;
        RECT 2495.5200 74.9000 2497.1200 75.3800 ;
        RECT 2495.5200 80.3400 2497.1200 80.8200 ;
        RECT 2495.5200 85.7800 2497.1200 86.2600 ;
        RECT 2495.5200 91.2200 2497.1200 91.7000 ;
        RECT 2495.5200 96.6600 2497.1200 97.1400 ;
        RECT 2495.5200 112.9800 2497.1200 113.4600 ;
        RECT 2495.5200 102.1000 2497.1200 102.5800 ;
        RECT 2495.5200 107.5400 2497.1200 108.0200 ;
        RECT 2495.5200 118.4200 2497.1200 118.9000 ;
        RECT 2495.5200 123.8600 2497.1200 124.3400 ;
        RECT 2384.4400 129.3000 2386.0400 129.7800 ;
        RECT 2384.4400 134.7400 2386.0400 135.2200 ;
        RECT 2374.3800 149.8400 2375.9800 150.3200 ;
        RECT 2384.4400 145.6200 2386.0400 146.1000 ;
        RECT 2384.4400 140.3300 2386.0400 140.8100 ;
        RECT 2384.4400 151.0600 2386.0400 151.5400 ;
        RECT 2384.4400 156.5000 2386.0400 156.9800 ;
        RECT 2384.4400 161.9400 2386.0400 162.4200 ;
        RECT 2384.4400 172.8200 2386.0400 173.3000 ;
        RECT 2444.5800 178.2600 2446.1800 180.2000 ;
        RECT 2444.5800 129.3000 2446.1800 129.7800 ;
        RECT 2444.5800 134.7400 2446.1800 135.2200 ;
        RECT 2444.5800 140.1800 2446.1800 140.6600 ;
        RECT 2444.5800 145.6200 2446.1800 146.1000 ;
        RECT 2444.5800 151.0600 2446.1800 151.5400 ;
        RECT 2444.5800 156.5000 2446.1800 156.9800 ;
        RECT 2444.5800 161.9400 2446.1800 162.4200 ;
        RECT 2444.5800 167.3800 2446.1800 167.8600 ;
        RECT 2444.5800 172.8200 2446.1800 173.3000 ;
        RECT 2495.5200 129.3000 2497.1200 129.7800 ;
        RECT 2495.5200 134.7400 2497.1200 135.2200 ;
        RECT 2495.5200 140.1800 2497.1200 140.6600 ;
        RECT 2495.5200 145.6200 2497.1200 146.1000 ;
        RECT 2495.5200 151.0600 2497.1200 151.5400 ;
        RECT 2495.5200 156.5000 2497.1200 156.9800 ;
        RECT 2495.5200 161.9400 2497.1200 162.4200 ;
        RECT 2495.5200 167.3800 2497.1200 167.8600 ;
        RECT 2495.5200 172.8200 2497.1200 173.3000 ;
        RECT 2495.5200 178.2600 2497.1200 178.7400 ;
        RECT 2444.5800 183.7000 2446.1800 184.1800 ;
        RECT 2434.4200 192.8200 2436.0200 193.3000 ;
        RECT 2444.5800 194.5800 2446.1800 195.0600 ;
        RECT 2444.5800 200.0200 2446.1800 200.5000 ;
        RECT 2444.5800 205.4600 2446.1800 205.9400 ;
        RECT 2444.5800 210.9000 2446.1800 211.3800 ;
        RECT 2444.5800 216.3400 2446.1800 216.8200 ;
        RECT 2444.5800 221.7800 2446.1800 222.2600 ;
        RECT 2444.5800 227.2200 2446.1800 227.7000 ;
        RECT 2495.5200 183.7000 2497.1200 184.1800 ;
        RECT 2495.5200 189.1400 2497.1200 189.6200 ;
        RECT 2495.5200 194.5800 2497.1200 195.0600 ;
        RECT 2495.5200 200.0200 2497.1200 200.5000 ;
        RECT 2495.5200 205.4600 2497.1200 205.9400 ;
        RECT 2495.5200 210.9000 2497.1200 211.3800 ;
        RECT 2495.5200 216.3400 2497.1200 216.8200 ;
        RECT 2495.5200 221.7800 2497.1200 222.2600 ;
        RECT 2495.5200 227.2200 2497.1200 227.7000 ;
        RECT 2176.7800 422.4600 2178.3800 422.9400 ;
        RECT 2444.5800 232.6600 2446.1800 233.1400 ;
        RECT 2444.5800 238.1000 2446.1800 238.5800 ;
        RECT 2444.5800 243.5400 2446.1800 244.0200 ;
        RECT 2444.5800 248.9800 2446.1800 249.4600 ;
        RECT 2444.5800 254.4200 2446.1800 254.9000 ;
        RECT 2444.5800 270.7400 2446.1800 271.2200 ;
        RECT 2444.5800 259.8600 2446.1800 260.3400 ;
        RECT 2444.5800 265.3000 2446.1800 265.7800 ;
        RECT 2444.5800 276.1800 2446.1800 276.6600 ;
        RECT 2444.5800 281.6200 2446.1800 282.1000 ;
        RECT 2495.5200 232.6600 2497.1200 233.1400 ;
        RECT 2495.5200 238.1000 2497.1200 238.5800 ;
        RECT 2495.5200 243.5400 2497.1200 244.0200 ;
        RECT 2495.5200 248.9800 2497.1200 249.4600 ;
        RECT 2495.5200 254.4200 2497.1200 254.9000 ;
        RECT 2495.5200 270.7400 2497.1200 271.2200 ;
        RECT 2495.5200 259.8600 2497.1200 260.3400 ;
        RECT 2495.5200 265.3000 2497.1200 265.7800 ;
        RECT 2495.5200 276.1800 2497.1200 276.6600 ;
        RECT 2495.5200 281.6200 2497.1200 282.1000 ;
        RECT 2444.5800 287.0600 2446.1800 287.5400 ;
        RECT 2444.5800 292.5000 2446.1800 292.9800 ;
        RECT 2444.5800 297.9400 2446.1800 298.4200 ;
        RECT 2444.5800 303.3800 2446.1800 303.8600 ;
        RECT 2444.5800 308.8200 2446.1800 309.3000 ;
        RECT 2444.5800 314.2600 2446.1800 314.7400 ;
        RECT 2444.5800 319.7000 2446.1800 320.1800 ;
        RECT 2444.5800 325.1400 2446.1800 325.6200 ;
        RECT 2444.5800 330.5800 2446.1800 331.0600 ;
        RECT 2444.5800 336.0200 2446.1800 336.5000 ;
        RECT 2495.5200 287.0600 2497.1200 287.5400 ;
        RECT 2495.5200 292.5000 2497.1200 292.9800 ;
        RECT 2495.5200 297.9400 2497.1200 298.4200 ;
        RECT 2495.5200 303.3800 2497.1200 303.8600 ;
        RECT 2495.5200 308.8200 2497.1200 309.3000 ;
        RECT 2495.5200 314.2600 2497.1200 314.7400 ;
        RECT 2495.5200 319.7000 2497.1200 320.1800 ;
        RECT 2495.5200 325.1400 2497.1200 325.6200 ;
        RECT 2495.5200 330.5800 2497.1200 331.0600 ;
        RECT 2495.5200 336.0200 2497.1200 336.5000 ;
        RECT 2444.5800 363.2200 2446.1800 363.7000 ;
        RECT 2444.5800 341.4600 2446.1800 341.9400 ;
        RECT 2444.5800 346.9000 2446.1800 347.3800 ;
        RECT 2444.5800 352.3400 2446.1800 352.8200 ;
        RECT 2444.5800 357.7800 2446.1800 358.2600 ;
        RECT 2444.5800 368.6600 2446.1800 369.1400 ;
        RECT 2444.5800 374.1000 2446.1800 374.5800 ;
        RECT 2444.5800 379.5400 2446.1800 380.0200 ;
        RECT 2444.5800 384.9800 2446.1800 385.4600 ;
        RECT 2495.5200 363.2200 2497.1200 363.7000 ;
        RECT 2495.5200 341.4600 2497.1200 341.9400 ;
        RECT 2495.5200 346.9000 2497.1200 347.3800 ;
        RECT 2495.5200 352.3400 2497.1200 352.8200 ;
        RECT 2495.5200 357.7800 2497.1200 358.2600 ;
        RECT 2495.5200 368.6600 2497.1200 369.1400 ;
        RECT 2495.5200 374.1000 2497.1200 374.5800 ;
        RECT 2495.5200 379.5400 2497.1200 380.0200 ;
        RECT 2495.5200 384.9800 2497.1200 385.4600 ;
        RECT 2444.5800 390.4200 2446.1800 390.9000 ;
        RECT 2444.5800 401.3000 2446.1800 401.7800 ;
        RECT 2444.5800 407.9300 2446.1800 409.8400 ;
        RECT 2444.5800 412.1800 2446.1800 412.6600 ;
        RECT 2434.4200 422.4600 2436.0200 422.9400 ;
        RECT 2444.5800 428.5000 2446.1800 428.9800 ;
        RECT 2444.5800 423.0600 2446.1800 423.5400 ;
        RECT 2444.5800 417.7900 2446.1800 419.8700 ;
        RECT 2444.5800 433.9400 2446.1800 434.4200 ;
        RECT 2444.5800 439.3800 2446.1800 439.8600 ;
        RECT 2495.5200 390.4200 2497.1200 390.9000 ;
        RECT 2495.5200 395.8600 2497.1200 396.3400 ;
        RECT 2495.5200 401.3000 2497.1200 401.7800 ;
        RECT 2495.5200 406.7400 2497.1200 407.2200 ;
        RECT 2495.5200 412.1800 2497.1200 412.6600 ;
        RECT 2495.5200 417.6200 2497.1200 418.1000 ;
        RECT 2495.5200 423.0600 2497.1200 423.5400 ;
        RECT 2495.5200 428.5000 2497.1200 428.9800 ;
        RECT 2495.5200 433.9400 2497.1200 434.4200 ;
        RECT 2495.5200 439.3800 2497.1200 439.8600 ;
        RECT 3365.4200 20.5000 3368.4200 20.9800 ;
        RECT 3303.1200 20.5000 3304.7200 20.9800 ;
        RECT 3303.1200 9.6200 3304.7200 10.1000 ;
        RECT 3303.1200 15.0600 3304.7200 15.5400 ;
        RECT 3365.4200 9.6200 3368.4200 10.1000 ;
        RECT 3365.4200 15.0600 3368.4200 15.5400 ;
        RECT 3303.1200 25.9400 3304.7200 26.4200 ;
        RECT 3303.1200 31.3800 3304.7200 31.8600 ;
        RECT 3303.1200 36.8200 3304.7200 37.3000 ;
        RECT 3303.1200 42.2600 3304.7200 42.7400 ;
        RECT 3303.1200 47.7000 3304.7200 48.1800 ;
        RECT 3303.1200 53.1400 3304.7200 53.6200 ;
        RECT 3303.1200 58.5800 3304.7200 59.0600 ;
        RECT 3303.1200 64.0200 3304.7200 64.5000 ;
        RECT 3303.1200 69.4600 3304.7200 69.9400 ;
        RECT 3365.4200 25.9400 3368.4200 26.4200 ;
        RECT 3365.4200 31.3800 3368.4200 31.8600 ;
        RECT 3365.4200 36.8200 3368.4200 37.3000 ;
        RECT 3365.4200 42.2600 3368.4200 42.7400 ;
        RECT 3365.4200 47.7000 3368.4200 48.1800 ;
        RECT 3365.4200 53.1400 3368.4200 53.6200 ;
        RECT 3365.4200 58.5800 3368.4200 59.0600 ;
        RECT 3365.4200 64.0200 3368.4200 64.5000 ;
        RECT 3365.4200 69.4600 3368.4200 69.9400 ;
        RECT 3303.1200 74.9000 3304.7200 75.3800 ;
        RECT 3303.1200 80.3400 3304.7200 80.8200 ;
        RECT 3303.1200 85.7800 3304.7200 86.2600 ;
        RECT 3303.1200 91.2200 3304.7200 91.7000 ;
        RECT 3303.1200 96.6600 3304.7200 97.1400 ;
        RECT 3303.1200 112.9800 3304.7200 113.4600 ;
        RECT 3303.1200 102.1000 3304.7200 102.5800 ;
        RECT 3303.1200 107.5400 3304.7200 108.0200 ;
        RECT 3303.1200 118.4200 3304.7200 118.9000 ;
        RECT 3303.1200 123.8600 3304.7200 124.3400 ;
        RECT 3365.4200 74.9000 3368.4200 75.3800 ;
        RECT 3365.4200 80.3400 3368.4200 80.8200 ;
        RECT 3365.4200 85.7800 3368.4200 86.2600 ;
        RECT 3365.4200 91.2200 3368.4200 91.7000 ;
        RECT 3365.4200 96.6600 3368.4200 97.1400 ;
        RECT 3365.4200 112.9800 3368.4200 113.4600 ;
        RECT 3365.4200 102.1000 3368.4200 102.5800 ;
        RECT 3365.4200 107.5400 3368.4200 108.0200 ;
        RECT 3365.4200 118.4200 3368.4200 118.9000 ;
        RECT 3365.4200 123.8600 3368.4200 124.3400 ;
        RECT 3303.1200 129.3000 3304.7200 129.7800 ;
        RECT 3303.1200 134.7400 3304.7200 135.2200 ;
        RECT 3303.1200 140.1800 3304.7200 140.6600 ;
        RECT 3303.1200 145.6200 3304.7200 146.1000 ;
        RECT 3303.1200 151.0600 3304.7200 151.5400 ;
        RECT 3303.1200 156.5000 3304.7200 156.9800 ;
        RECT 3303.1200 161.9400 3304.7200 162.4200 ;
        RECT 3303.1200 167.3800 3304.7200 167.8600 ;
        RECT 3303.1200 172.8200 3304.7200 173.3000 ;
        RECT 3303.1200 178.2600 3304.7200 178.7400 ;
        RECT 3365.4200 129.3000 3368.4200 129.7800 ;
        RECT 3365.4200 134.7400 3368.4200 135.2200 ;
        RECT 3365.4200 140.1800 3368.4200 140.6600 ;
        RECT 3365.4200 145.6200 3368.4200 146.1000 ;
        RECT 3365.4200 151.0600 3368.4200 151.5400 ;
        RECT 3365.4200 156.5000 3368.4200 156.9800 ;
        RECT 3365.4200 161.9400 3368.4200 162.4200 ;
        RECT 3365.4200 167.3800 3368.4200 167.8600 ;
        RECT 3365.4200 172.8200 3368.4200 173.3000 ;
        RECT 3365.4200 178.2600 3368.4200 178.7400 ;
        RECT 3303.1200 183.7000 3304.7200 184.1800 ;
        RECT 3303.1200 189.1400 3304.7200 189.6200 ;
        RECT 3303.1200 194.5800 3304.7200 195.0600 ;
        RECT 3303.1200 200.0200 3304.7200 200.5000 ;
        RECT 3303.1200 205.4600 3304.7200 205.9400 ;
        RECT 3303.1200 210.9000 3304.7200 211.3800 ;
        RECT 3303.1200 216.3400 3304.7200 216.8200 ;
        RECT 3303.1200 221.7800 3304.7200 222.2600 ;
        RECT 3303.1200 227.2200 3304.7200 227.7000 ;
        RECT 3365.4200 183.7000 3368.4200 184.1800 ;
        RECT 3365.4200 189.1400 3368.4200 189.6200 ;
        RECT 3365.4200 194.5800 3368.4200 195.0600 ;
        RECT 3365.4200 200.0200 3368.4200 200.5000 ;
        RECT 3365.4200 205.4600 3368.4200 205.9400 ;
        RECT 3365.4200 210.9000 3368.4200 211.3800 ;
        RECT 3365.4200 216.3400 3368.4200 216.8200 ;
        RECT 3365.4200 221.7800 3368.4200 222.2600 ;
        RECT 3365.4200 227.2200 3368.4200 227.7000 ;
        RECT 3303.1200 232.6600 3304.7200 233.1400 ;
        RECT 3303.1200 238.1000 3304.7200 238.5800 ;
        RECT 3303.1200 243.5400 3304.7200 244.0200 ;
        RECT 3303.1200 248.9800 3304.7200 249.4600 ;
        RECT 3303.1200 254.4200 3304.7200 254.9000 ;
        RECT 3303.1200 270.7400 3304.7200 271.2200 ;
        RECT 3303.1200 259.8600 3304.7200 260.3400 ;
        RECT 3303.1200 265.3000 3304.7200 265.7800 ;
        RECT 3303.1200 276.1800 3304.7200 276.6600 ;
        RECT 3303.1200 281.6200 3304.7200 282.1000 ;
        RECT 3365.4200 232.6600 3368.4200 233.1400 ;
        RECT 3365.4200 238.1000 3368.4200 238.5800 ;
        RECT 3365.4200 243.5400 3368.4200 244.0200 ;
        RECT 3365.4200 248.9800 3368.4200 249.4600 ;
        RECT 3365.4200 254.4200 3368.4200 254.9000 ;
        RECT 3365.4200 270.7400 3368.4200 271.2200 ;
        RECT 3365.4200 259.8600 3368.4200 260.3400 ;
        RECT 3365.4200 265.3000 3368.4200 265.7800 ;
        RECT 3365.4200 276.1800 3368.4200 276.6600 ;
        RECT 3365.4200 281.6200 3368.4200 282.1000 ;
        RECT 3303.1200 287.0600 3304.7200 287.5400 ;
        RECT 3303.1200 292.5000 3304.7200 292.9800 ;
        RECT 3303.1200 297.9400 3304.7200 298.4200 ;
        RECT 3303.1200 303.3800 3304.7200 303.8600 ;
        RECT 3303.1200 308.8200 3304.7200 309.3000 ;
        RECT 3303.1200 314.2600 3304.7200 314.7400 ;
        RECT 3303.1200 319.7000 3304.7200 320.1800 ;
        RECT 3303.1200 325.1400 3304.7200 325.6200 ;
        RECT 3303.1200 330.5800 3304.7200 331.0600 ;
        RECT 3303.1200 336.0200 3304.7200 336.5000 ;
        RECT 3365.4200 287.0600 3368.4200 287.5400 ;
        RECT 3365.4200 292.5000 3368.4200 292.9800 ;
        RECT 3365.4200 297.9400 3368.4200 298.4200 ;
        RECT 3365.4200 303.3800 3368.4200 303.8600 ;
        RECT 3365.4200 308.8200 3368.4200 309.3000 ;
        RECT 3365.4200 314.2600 3368.4200 314.7400 ;
        RECT 3365.4200 319.7000 3368.4200 320.1800 ;
        RECT 3365.4200 325.1400 3368.4200 325.6200 ;
        RECT 3365.4200 330.5800 3368.4200 331.0600 ;
        RECT 3365.4200 336.0200 3368.4200 336.5000 ;
        RECT 3303.1200 363.2200 3304.7200 363.7000 ;
        RECT 3303.1200 341.4600 3304.7200 341.9400 ;
        RECT 3303.1200 346.9000 3304.7200 347.3800 ;
        RECT 3303.1200 352.3400 3304.7200 352.8200 ;
        RECT 3303.1200 357.7800 3304.7200 358.2600 ;
        RECT 3303.1200 368.6600 3304.7200 369.1400 ;
        RECT 3303.1200 374.1000 3304.7200 374.5800 ;
        RECT 3303.1200 379.5400 3304.7200 380.0200 ;
        RECT 3303.1200 384.9800 3304.7200 385.4600 ;
        RECT 3365.4200 363.2200 3368.4200 363.7000 ;
        RECT 3365.4200 341.4600 3368.4200 341.9400 ;
        RECT 3365.4200 346.9000 3368.4200 347.3800 ;
        RECT 3365.4200 352.3400 3368.4200 352.8200 ;
        RECT 3365.4200 357.7800 3368.4200 358.2600 ;
        RECT 3365.4200 368.6600 3368.4200 369.1400 ;
        RECT 3365.4200 374.1000 3368.4200 374.5800 ;
        RECT 3365.4200 379.5400 3368.4200 380.0200 ;
        RECT 3365.4200 384.9800 3368.4200 385.4600 ;
        RECT 3303.1200 390.4200 3304.7200 390.9000 ;
        RECT 3303.1200 395.8600 3304.7200 396.3400 ;
        RECT 3303.1200 401.3000 3304.7200 401.7800 ;
        RECT 3303.1200 406.7400 3304.7200 407.2200 ;
        RECT 3303.1200 412.1800 3304.7200 412.6600 ;
        RECT 3303.1200 417.6200 3304.7200 418.1000 ;
        RECT 3303.1200 423.0600 3304.7200 423.5400 ;
        RECT 3303.1200 428.5000 3304.7200 428.9800 ;
        RECT 3303.1200 433.9400 3304.7200 434.4200 ;
        RECT 3303.1200 439.3800 3304.7200 439.8600 ;
        RECT 3365.4200 390.4200 3368.4200 390.9000 ;
        RECT 3365.4200 395.8600 3368.4200 396.3400 ;
        RECT 3365.4200 401.3000 3368.4200 401.7800 ;
        RECT 3365.4200 406.7400 3368.4200 407.2200 ;
        RECT 3365.4200 412.1800 3368.4200 412.6600 ;
        RECT 3365.4200 417.6200 3368.4200 418.1000 ;
        RECT 3365.4200 423.0600 3368.4200 423.5400 ;
        RECT 3365.4200 428.5000 3368.4200 428.9800 ;
        RECT 3365.4200 433.9400 3368.4200 434.4200 ;
        RECT 3365.4200 439.3800 3368.4200 439.8600 ;
        RECT 1736.3400 652.1000 1737.9400 652.5800 ;
        RECT 1944.0000 624.7700 1945.6000 627.4200 ;
        RECT 1956.5600 652.1000 1958.1600 652.5800 ;
        RECT 2164.2200 624.7700 2165.8200 627.4200 ;
        RECT 2176.7800 652.1000 2178.3800 652.5800 ;
        RECT 2444.5800 444.8200 2446.1800 445.3000 ;
        RECT 2444.5800 450.2600 2446.1800 450.7400 ;
        RECT 2444.5800 455.7000 2446.1800 456.1800 ;
        RECT 2444.5800 461.1400 2446.1800 461.6200 ;
        RECT 2444.5800 466.5800 2446.1800 467.0600 ;
        RECT 2444.5800 472.0200 2446.1800 472.5000 ;
        RECT 2444.5800 477.4600 2446.1800 477.9400 ;
        RECT 2444.5800 482.9000 2446.1800 483.3800 ;
        RECT 2444.5800 488.3400 2446.1800 488.8200 ;
        RECT 2444.5800 493.7800 2446.1800 494.2600 ;
        RECT 2495.5200 444.8200 2497.1200 445.3000 ;
        RECT 2495.5200 450.2600 2497.1200 450.7400 ;
        RECT 2495.5200 455.7000 2497.1200 456.1800 ;
        RECT 2495.5200 461.1400 2497.1200 461.6200 ;
        RECT 2495.5200 466.5800 2497.1200 467.0600 ;
        RECT 2495.5200 472.0200 2497.1200 472.5000 ;
        RECT 2495.5200 477.4600 2497.1200 477.9400 ;
        RECT 2495.5200 482.9000 2497.1200 483.3800 ;
        RECT 2495.5200 488.3400 2497.1200 488.8200 ;
        RECT 2495.5200 493.7800 2497.1200 494.2600 ;
        RECT 2444.5800 520.9800 2446.1800 521.4600 ;
        RECT 2444.5800 499.2200 2446.1800 499.7000 ;
        RECT 2444.5800 504.6600 2446.1800 505.1400 ;
        RECT 2444.5800 510.1000 2446.1800 510.5800 ;
        RECT 2444.5800 515.5400 2446.1800 516.0200 ;
        RECT 2444.5800 526.4200 2446.1800 526.9000 ;
        RECT 2444.5800 531.8600 2446.1800 532.3400 ;
        RECT 2444.5800 537.3000 2446.1800 537.7800 ;
        RECT 2444.5800 542.7400 2446.1800 543.2200 ;
        RECT 2495.5200 520.9800 2497.1200 521.4600 ;
        RECT 2495.5200 499.2200 2497.1200 499.7000 ;
        RECT 2495.5200 504.6600 2497.1200 505.1400 ;
        RECT 2495.5200 510.1000 2497.1200 510.5800 ;
        RECT 2495.5200 515.5400 2497.1200 516.0200 ;
        RECT 2495.5200 526.4200 2497.1200 526.9000 ;
        RECT 2495.5200 531.8600 2497.1200 532.3400 ;
        RECT 2495.5200 537.3000 2497.1200 537.7800 ;
        RECT 2495.5200 542.7400 2497.1200 543.2200 ;
        RECT 2444.5800 548.1800 2446.1800 548.6600 ;
        RECT 2444.5800 553.6200 2446.1800 554.1000 ;
        RECT 2444.5800 559.0600 2446.1800 559.5400 ;
        RECT 2444.5800 564.5000 2446.1800 564.9800 ;
        RECT 2444.5800 569.9400 2446.1800 570.4200 ;
        RECT 2444.5800 575.3800 2446.1800 575.8600 ;
        RECT 2444.5800 580.8200 2446.1800 581.3000 ;
        RECT 2444.5800 586.2600 2446.1800 586.7400 ;
        RECT 2444.5800 591.7000 2446.1800 592.1800 ;
        RECT 2444.5800 597.1400 2446.1800 597.6200 ;
        RECT 2495.5200 548.1800 2497.1200 548.6600 ;
        RECT 2495.5200 553.6200 2497.1200 554.1000 ;
        RECT 2495.5200 559.0600 2497.1200 559.5400 ;
        RECT 2495.5200 564.5000 2497.1200 564.9800 ;
        RECT 2495.5200 569.9400 2497.1200 570.4200 ;
        RECT 2495.5200 575.3800 2497.1200 575.8600 ;
        RECT 2495.5200 580.8200 2497.1200 581.3000 ;
        RECT 2495.5200 586.2600 2497.1200 586.7400 ;
        RECT 2495.5200 591.7000 2497.1200 592.1800 ;
        RECT 2495.5200 597.1400 2497.1200 597.6200 ;
        RECT 2444.5800 602.5800 2446.1800 603.0600 ;
        RECT 2444.5800 608.0200 2446.1800 608.5000 ;
        RECT 2444.5800 613.4600 2446.1800 613.9400 ;
        RECT 2444.5800 618.9000 2446.1800 619.3800 ;
        RECT 2444.5800 624.3400 2446.1800 626.3700 ;
        RECT 2444.5800 629.7800 2446.1800 630.2600 ;
        RECT 2444.5800 634.4300 2446.1800 634.9100 ;
        RECT 2434.4200 652.1000 2436.0200 652.5800 ;
        RECT 2444.5800 640.6600 2446.1800 641.1400 ;
        RECT 2444.5800 647.6300 2446.1800 649.5100 ;
        RECT 2444.5800 651.5400 2446.1800 652.0200 ;
        RECT 2495.5200 602.5800 2497.1200 603.0600 ;
        RECT 2495.5200 608.0200 2497.1200 608.5000 ;
        RECT 2495.5200 613.4600 2497.1200 613.9400 ;
        RECT 2495.5200 618.9000 2497.1200 619.3800 ;
        RECT 2495.5200 624.3400 2497.1200 624.8200 ;
        RECT 2495.5200 629.7800 2497.1200 630.2600 ;
        RECT 2495.5200 635.2200 2497.1200 635.7000 ;
        RECT 2495.5200 640.6600 2497.1200 641.1400 ;
        RECT 2495.5200 646.1000 2497.1200 646.5800 ;
        RECT 2495.5200 651.5400 2497.1200 652.0200 ;
        RECT 2444.5800 656.9800 2446.1800 657.4600 ;
        RECT 2444.5800 662.4200 2446.1800 662.9000 ;
        RECT 2444.5800 667.8600 2446.1800 668.3400 ;
        RECT 2444.5800 673.3000 2446.1800 673.7800 ;
        RECT 2444.5800 678.7400 2446.1800 679.2200 ;
        RECT 2444.5800 684.1800 2446.1800 684.6600 ;
        RECT 2444.5800 689.6200 2446.1800 690.1000 ;
        RECT 2444.5800 695.0600 2446.1800 695.5400 ;
        RECT 2444.5800 700.5000 2446.1800 700.9800 ;
        RECT 2495.5200 656.9800 2497.1200 657.4600 ;
        RECT 2495.5200 662.4200 2497.1200 662.9000 ;
        RECT 2495.5200 667.8600 2497.1200 668.3400 ;
        RECT 2495.5200 673.3000 2497.1200 673.7800 ;
        RECT 2495.5200 678.7400 2497.1200 679.2200 ;
        RECT 2495.5200 684.1800 2497.1200 684.6600 ;
        RECT 2495.5200 689.6200 2497.1200 690.1000 ;
        RECT 2495.5200 695.0600 2497.1200 695.5400 ;
        RECT 2495.5200 700.5000 2497.1200 700.9800 ;
        RECT 2444.5800 705.9400 2446.1800 706.4200 ;
        RECT 2444.5800 711.3800 2446.1800 711.8600 ;
        RECT 2444.5800 716.8200 2446.1800 717.3000 ;
        RECT 2444.5800 722.2600 2446.1800 722.7400 ;
        RECT 2444.5800 727.7000 2446.1800 728.1800 ;
        RECT 2444.5800 733.1400 2446.1800 733.6200 ;
        RECT 2444.5800 738.5800 2446.1800 739.0600 ;
        RECT 2444.5800 744.0200 2446.1800 744.5000 ;
        RECT 2444.5800 749.4600 2446.1800 749.9400 ;
        RECT 2495.5200 705.9400 2497.1200 706.4200 ;
        RECT 2495.5200 711.3800 2497.1200 711.8600 ;
        RECT 2495.5200 716.8200 2497.1200 717.3000 ;
        RECT 2495.5200 722.2600 2497.1200 722.7400 ;
        RECT 2495.5200 727.7000 2497.1200 728.1800 ;
        RECT 2495.5200 744.0200 2497.1200 744.5000 ;
        RECT 2495.5200 738.5800 2497.1200 739.0600 ;
        RECT 2495.5200 733.1400 2497.1200 733.6200 ;
        RECT 2495.5200 749.4600 2497.1200 749.9400 ;
        RECT 1736.3400 881.7400 1737.9400 882.2200 ;
        RECT 1736.3400 1111.3800 1737.9400 1111.8600 ;
        RECT 1944.0000 1084.0500 1945.6000 1086.7000 ;
        RECT 1956.5600 1111.3800 1958.1600 1111.8600 ;
        RECT 2176.7800 881.7400 2178.3800 882.2200 ;
        RECT 2434.4200 881.7400 2436.0200 882.2200 ;
        RECT 2164.2200 1084.0500 2165.8200 1086.7000 ;
        RECT 2176.7800 1111.3800 2178.3800 1111.8600 ;
        RECT 2434.4200 1111.3800 2436.0200 1111.8600 ;
        RECT 3303.1200 444.8200 3304.7200 445.3000 ;
        RECT 3303.1200 450.2600 3304.7200 450.7400 ;
        RECT 3303.1200 455.7000 3304.7200 456.1800 ;
        RECT 3303.1200 461.1400 3304.7200 461.6200 ;
        RECT 3303.1200 466.5800 3304.7200 467.0600 ;
        RECT 3303.1200 472.0200 3304.7200 472.5000 ;
        RECT 3303.1200 477.4600 3304.7200 477.9400 ;
        RECT 3303.1200 482.9000 3304.7200 483.3800 ;
        RECT 3303.1200 488.3400 3304.7200 488.8200 ;
        RECT 3303.1200 493.7800 3304.7200 494.2600 ;
        RECT 3365.4200 444.8200 3368.4200 445.3000 ;
        RECT 3365.4200 450.2600 3368.4200 450.7400 ;
        RECT 3365.4200 455.7000 3368.4200 456.1800 ;
        RECT 3365.4200 461.1400 3368.4200 461.6200 ;
        RECT 3365.4200 466.5800 3368.4200 467.0600 ;
        RECT 3365.4200 472.0200 3368.4200 472.5000 ;
        RECT 3365.4200 477.4600 3368.4200 477.9400 ;
        RECT 3365.4200 482.9000 3368.4200 483.3800 ;
        RECT 3365.4200 488.3400 3368.4200 488.8200 ;
        RECT 3365.4200 493.7800 3368.4200 494.2600 ;
        RECT 3303.1200 520.9800 3304.7200 521.4600 ;
        RECT 3303.1200 499.2200 3304.7200 499.7000 ;
        RECT 3303.1200 504.6600 3304.7200 505.1400 ;
        RECT 3303.1200 510.1000 3304.7200 510.5800 ;
        RECT 3303.1200 515.5400 3304.7200 516.0200 ;
        RECT 3303.1200 526.4200 3304.7200 526.9000 ;
        RECT 3303.1200 531.8600 3304.7200 532.3400 ;
        RECT 3303.1200 537.3000 3304.7200 537.7800 ;
        RECT 3303.1200 542.7400 3304.7200 543.2200 ;
        RECT 3365.4200 520.9800 3368.4200 521.4600 ;
        RECT 3365.4200 499.2200 3368.4200 499.7000 ;
        RECT 3365.4200 504.6600 3368.4200 505.1400 ;
        RECT 3365.4200 510.1000 3368.4200 510.5800 ;
        RECT 3365.4200 515.5400 3368.4200 516.0200 ;
        RECT 3365.4200 526.4200 3368.4200 526.9000 ;
        RECT 3365.4200 531.8600 3368.4200 532.3400 ;
        RECT 3365.4200 537.3000 3368.4200 537.7800 ;
        RECT 3365.4200 542.7400 3368.4200 543.2200 ;
        RECT 3303.1200 548.1800 3304.7200 548.6600 ;
        RECT 3303.1200 553.6200 3304.7200 554.1000 ;
        RECT 3303.1200 559.0600 3304.7200 559.5400 ;
        RECT 3303.1200 564.5000 3304.7200 564.9800 ;
        RECT 3303.1200 569.9400 3304.7200 570.4200 ;
        RECT 3303.1200 575.3800 3304.7200 575.8600 ;
        RECT 3303.1200 580.8200 3304.7200 581.3000 ;
        RECT 3303.1200 586.2600 3304.7200 586.7400 ;
        RECT 3303.1200 591.7000 3304.7200 592.1800 ;
        RECT 3303.1200 597.1400 3304.7200 597.6200 ;
        RECT 3365.4200 548.1800 3368.4200 548.6600 ;
        RECT 3365.4200 553.6200 3368.4200 554.1000 ;
        RECT 3365.4200 559.0600 3368.4200 559.5400 ;
        RECT 3365.4200 564.5000 3368.4200 564.9800 ;
        RECT 3365.4200 569.9400 3368.4200 570.4200 ;
        RECT 3365.4200 575.3800 3368.4200 575.8600 ;
        RECT 3365.4200 580.8200 3368.4200 581.3000 ;
        RECT 3365.4200 586.2600 3368.4200 586.7400 ;
        RECT 3365.4200 591.7000 3368.4200 592.1800 ;
        RECT 3365.4200 597.1400 3368.4200 597.6200 ;
        RECT 3303.1200 602.5800 3304.7200 603.0600 ;
        RECT 3303.1200 608.0200 3304.7200 608.5000 ;
        RECT 3303.1200 613.4600 3304.7200 613.9400 ;
        RECT 3303.1200 618.9000 3304.7200 619.3800 ;
        RECT 3303.1200 624.3400 3304.7200 624.8200 ;
        RECT 3303.1200 629.7800 3304.7200 630.2600 ;
        RECT 3303.1200 635.2200 3304.7200 635.7000 ;
        RECT 3303.1200 640.6600 3304.7200 641.1400 ;
        RECT 3303.1200 646.1000 3304.7200 646.5800 ;
        RECT 3303.1200 651.5400 3304.7200 652.0200 ;
        RECT 3365.4200 602.5800 3368.4200 603.0600 ;
        RECT 3365.4200 608.0200 3368.4200 608.5000 ;
        RECT 3365.4200 613.4600 3368.4200 613.9400 ;
        RECT 3365.4200 618.9000 3368.4200 619.3800 ;
        RECT 3365.4200 624.3400 3368.4200 624.8200 ;
        RECT 3365.4200 629.7800 3368.4200 630.2600 ;
        RECT 3365.4200 635.2200 3368.4200 635.7000 ;
        RECT 3365.4200 640.6600 3368.4200 641.1400 ;
        RECT 3365.4200 646.1000 3368.4200 646.5800 ;
        RECT 3365.4200 651.5400 3368.4200 652.0200 ;
        RECT 3303.1200 656.9800 3304.7200 657.4600 ;
        RECT 3303.1200 662.4200 3304.7200 662.9000 ;
        RECT 3303.1200 667.8600 3304.7200 668.3400 ;
        RECT 3303.1200 673.3000 3304.7200 673.7800 ;
        RECT 3303.1200 678.7400 3304.7200 679.2200 ;
        RECT 3303.1200 684.1800 3304.7200 684.6600 ;
        RECT 3303.1200 689.6200 3304.7200 690.1000 ;
        RECT 3303.1200 695.0600 3304.7200 695.5400 ;
        RECT 3303.1200 700.5000 3304.7200 700.9800 ;
        RECT 3365.4200 656.9800 3368.4200 657.4600 ;
        RECT 3365.4200 662.4200 3368.4200 662.9000 ;
        RECT 3365.4200 667.8600 3368.4200 668.3400 ;
        RECT 3365.4200 673.3000 3368.4200 673.7800 ;
        RECT 3365.4200 678.7400 3368.4200 679.2200 ;
        RECT 3365.4200 684.1800 3368.4200 684.6600 ;
        RECT 3365.4200 689.6200 3368.4200 690.1000 ;
        RECT 3365.4200 695.0600 3368.4200 695.5400 ;
        RECT 3365.4200 700.5000 3368.4200 700.9800 ;
        RECT 3303.1200 705.9400 3304.7200 706.4200 ;
        RECT 3303.1200 711.3800 3304.7200 711.8600 ;
        RECT 3303.1200 716.8200 3304.7200 717.3000 ;
        RECT 3303.1200 722.2600 3304.7200 722.7400 ;
        RECT 3303.1200 727.7000 3304.7200 728.1800 ;
        RECT 3303.1200 733.1400 3304.7200 733.6200 ;
        RECT 3303.1200 738.5800 3304.7200 739.0600 ;
        RECT 3303.1200 744.0200 3304.7200 744.5000 ;
        RECT 3303.1200 749.4600 3304.7200 749.9400 ;
        RECT 3303.1200 754.9000 3304.7200 755.3800 ;
        RECT 3365.4200 705.9400 3368.4200 706.4200 ;
        RECT 3365.4200 711.3800 3368.4200 711.8600 ;
        RECT 3365.4200 716.8200 3368.4200 717.3000 ;
        RECT 3365.4200 722.2600 3368.4200 722.7400 ;
        RECT 3365.4200 727.7000 3368.4200 728.1800 ;
        RECT 3365.4200 733.1400 3368.4200 733.6200 ;
        RECT 3365.4200 738.5800 3368.4200 739.0600 ;
        RECT 3365.4200 744.0200 3368.4200 744.5000 ;
        RECT 3365.4200 749.4600 3368.4200 749.9400 ;
        RECT 3365.4200 754.9000 3368.4200 755.3800 ;
        RECT 3303.1200 771.2200 3304.7200 771.7000 ;
        RECT 3303.1200 760.3400 3304.7200 760.8200 ;
        RECT 3303.1200 765.7800 3304.7200 766.2600 ;
        RECT 3303.1200 776.6600 3304.7200 777.1400 ;
        RECT 3303.1200 782.1000 3304.7200 782.5800 ;
        RECT 3303.1200 787.5400 3304.7200 788.0200 ;
        RECT 3303.1200 792.9800 3304.7200 793.4600 ;
        RECT 3303.1200 798.4200 3304.7200 798.9000 ;
        RECT 3303.1200 803.8600 3304.7200 804.3400 ;
        RECT 3303.1200 809.3000 3304.7200 809.7800 ;
        RECT 3365.4200 771.2200 3368.4200 771.7000 ;
        RECT 3365.4200 760.3400 3368.4200 760.8200 ;
        RECT 3365.4200 765.7800 3368.4200 766.2600 ;
        RECT 3365.4200 776.6600 3368.4200 777.1400 ;
        RECT 3365.4200 782.1000 3368.4200 782.5800 ;
        RECT 3365.4200 787.5400 3368.4200 788.0200 ;
        RECT 3365.4200 792.9800 3368.4200 793.4600 ;
        RECT 3365.4200 798.4200 3368.4200 798.9000 ;
        RECT 3365.4200 803.8600 3368.4200 804.3400 ;
        RECT 3365.4200 809.3000 3368.4200 809.7800 ;
        RECT 3303.1200 814.7400 3304.7200 815.2200 ;
        RECT 3303.1200 820.1800 3304.7200 820.6600 ;
        RECT 3303.1200 825.6200 3304.7200 826.1000 ;
        RECT 3303.1200 831.0600 3304.7200 831.5400 ;
        RECT 3303.1200 836.5000 3304.7200 836.9800 ;
        RECT 3303.1200 841.9400 3304.7200 842.4200 ;
        RECT 3303.1200 847.3800 3304.7200 847.8600 ;
        RECT 3303.1200 852.8200 3304.7200 853.3000 ;
        RECT 3303.1200 858.2600 3304.7200 858.7400 ;
        RECT 3365.4200 814.7400 3368.4200 815.2200 ;
        RECT 3365.4200 820.1800 3368.4200 820.6600 ;
        RECT 3365.4200 825.6200 3368.4200 826.1000 ;
        RECT 3365.4200 831.0600 3368.4200 831.5400 ;
        RECT 3365.4200 836.5000 3368.4200 836.9800 ;
        RECT 3365.4200 841.9400 3368.4200 842.4200 ;
        RECT 3365.4200 847.3800 3368.4200 847.8600 ;
        RECT 3365.4200 852.8200 3368.4200 853.3000 ;
        RECT 3365.4200 858.2600 3368.4200 858.7400 ;
        RECT 3303.1200 863.7000 3304.7200 864.1800 ;
        RECT 3303.1200 869.1400 3304.7200 869.6200 ;
        RECT 3303.1200 874.5800 3304.7200 875.0600 ;
        RECT 3303.1200 880.0200 3304.7200 880.5000 ;
        RECT 3303.1200 885.4600 3304.7200 885.9400 ;
        RECT 3303.1200 890.9000 3304.7200 891.3800 ;
        RECT 3303.1200 896.3400 3304.7200 896.8200 ;
        RECT 3303.1200 901.7800 3304.7200 902.2600 ;
        RECT 3303.1200 907.2200 3304.7200 907.7000 ;
        RECT 3303.1200 912.6600 3304.7200 913.1400 ;
        RECT 3365.4200 863.7000 3368.4200 864.1800 ;
        RECT 3365.4200 869.1400 3368.4200 869.6200 ;
        RECT 3365.4200 874.5800 3368.4200 875.0600 ;
        RECT 3365.4200 880.0200 3368.4200 880.5000 ;
        RECT 3365.4200 885.4600 3368.4200 885.9400 ;
        RECT 3365.4200 890.9000 3368.4200 891.3800 ;
        RECT 3365.4200 896.3400 3368.4200 896.8200 ;
        RECT 3365.4200 901.7800 3368.4200 902.2600 ;
        RECT 3365.4200 907.2200 3368.4200 907.7000 ;
        RECT 3365.4200 912.6600 3368.4200 913.1400 ;
        RECT 3303.1200 928.9800 3304.7200 929.4600 ;
        RECT 3303.1200 918.1000 3304.7200 918.5800 ;
        RECT 3303.1200 923.5400 3304.7200 924.0200 ;
        RECT 3303.1200 934.4200 3304.7200 934.9000 ;
        RECT 3303.1200 939.8600 3304.7200 940.3400 ;
        RECT 3303.1200 945.3000 3304.7200 945.7800 ;
        RECT 3303.1200 950.7400 3304.7200 951.2200 ;
        RECT 3303.1200 956.1800 3304.7200 956.6600 ;
        RECT 3303.1200 961.6200 3304.7200 962.1000 ;
        RECT 3303.1200 967.0600 3304.7200 967.5400 ;
        RECT 3365.4200 928.9800 3368.4200 929.4600 ;
        RECT 3365.4200 918.1000 3368.4200 918.5800 ;
        RECT 3365.4200 923.5400 3368.4200 924.0200 ;
        RECT 3365.4200 934.4200 3368.4200 934.9000 ;
        RECT 3365.4200 939.8600 3368.4200 940.3400 ;
        RECT 3365.4200 945.3000 3368.4200 945.7800 ;
        RECT 3365.4200 950.7400 3368.4200 951.2200 ;
        RECT 3365.4200 956.1800 3368.4200 956.6600 ;
        RECT 3365.4200 961.6200 3368.4200 962.1000 ;
        RECT 3365.4200 967.0600 3368.4200 967.5400 ;
        RECT 3365.4200 1021.4600 3368.4200 1021.9400 ;
        RECT 3303.1200 1021.4600 3304.7200 1021.9400 ;
        RECT 3303.1200 972.5000 3304.7200 972.9800 ;
        RECT 3303.1200 977.9400 3304.7200 978.4200 ;
        RECT 3303.1200 983.3800 3304.7200 983.8600 ;
        RECT 3303.1200 988.8200 3304.7200 989.3000 ;
        RECT 3303.1200 994.2600 3304.7200 994.7400 ;
        RECT 3303.1200 999.7000 3304.7200 1000.1800 ;
        RECT 3303.1200 1005.1400 3304.7200 1005.6200 ;
        RECT 3303.1200 1010.5800 3304.7200 1011.0600 ;
        RECT 3303.1200 1016.0200 3304.7200 1016.5000 ;
        RECT 3365.4200 972.5000 3368.4200 972.9800 ;
        RECT 3365.4200 977.9400 3368.4200 978.4200 ;
        RECT 3365.4200 983.3800 3368.4200 983.8600 ;
        RECT 3365.4200 988.8200 3368.4200 989.3000 ;
        RECT 3365.4200 994.2600 3368.4200 994.7400 ;
        RECT 3365.4200 999.7000 3368.4200 1000.1800 ;
        RECT 3365.4200 1005.1400 3368.4200 1005.6200 ;
        RECT 3365.4200 1010.5800 3368.4200 1011.0600 ;
        RECT 3365.4200 1016.0200 3368.4200 1016.5000 ;
        RECT 3303.1200 1026.9000 3304.7200 1027.3800 ;
        RECT 3303.1200 1032.3400 3304.7200 1032.8200 ;
        RECT 3303.1200 1037.7800 3304.7200 1038.2600 ;
        RECT 3303.1200 1043.2200 3304.7200 1043.7000 ;
        RECT 3303.1200 1048.6600 3304.7200 1049.1400 ;
        RECT 3303.1200 1054.1000 3304.7200 1054.5800 ;
        RECT 3303.1200 1059.5400 3304.7200 1060.0200 ;
        RECT 3303.1200 1064.9800 3304.7200 1065.4600 ;
        RECT 3303.1200 1070.4200 3304.7200 1070.9000 ;
        RECT 3365.4200 1026.9000 3368.4200 1027.3800 ;
        RECT 3365.4200 1032.3400 3368.4200 1032.8200 ;
        RECT 3365.4200 1037.7800 3368.4200 1038.2600 ;
        RECT 3365.4200 1043.2200 3368.4200 1043.7000 ;
        RECT 3365.4200 1048.6600 3368.4200 1049.1400 ;
        RECT 3365.4200 1054.1000 3368.4200 1054.5800 ;
        RECT 3365.4200 1059.5400 3368.4200 1060.0200 ;
        RECT 3365.4200 1064.9800 3368.4200 1065.4600 ;
        RECT 3365.4200 1070.4200 3368.4200 1070.9000 ;
        RECT 3365.4200 1179.2200 3368.4200 1179.7000 ;
        RECT 3303.1200 1179.2200 3304.7200 1179.7000 ;
        RECT 3303.1200 1075.8600 3304.7200 1076.3400 ;
        RECT 3303.1200 1081.3000 3304.7200 1081.7800 ;
        RECT 3303.1200 1086.7400 3304.7200 1087.2200 ;
        RECT 3303.1200 1092.1800 3304.7200 1092.6600 ;
        RECT 3303.1200 1097.6200 3304.7200 1098.1000 ;
        RECT 3303.1200 1103.0600 3304.7200 1103.5400 ;
        RECT 3303.1200 1108.5000 3304.7200 1108.9800 ;
        RECT 3303.1200 1113.9400 3304.7200 1114.4200 ;
        RECT 3303.1200 1119.3800 3304.7200 1119.8600 ;
        RECT 3303.1200 1124.8200 3304.7200 1125.3000 ;
        RECT 3365.4200 1075.8600 3368.4200 1076.3400 ;
        RECT 3365.4200 1081.3000 3368.4200 1081.7800 ;
        RECT 3365.4200 1086.7400 3368.4200 1087.2200 ;
        RECT 3365.4200 1092.1800 3368.4200 1092.6600 ;
        RECT 3365.4200 1097.6200 3368.4200 1098.1000 ;
        RECT 3365.4200 1103.0600 3368.4200 1103.5400 ;
        RECT 3365.4200 1108.5000 3368.4200 1108.9800 ;
        RECT 3365.4200 1113.9400 3368.4200 1114.4200 ;
        RECT 3365.4200 1119.3800 3368.4200 1119.8600 ;
        RECT 3365.4200 1124.8200 3368.4200 1125.3000 ;
        RECT 3303.1200 1130.2600 3304.7200 1130.7400 ;
        RECT 3303.1200 1135.7000 3304.7200 1136.1800 ;
        RECT 3303.1200 1141.1400 3304.7200 1141.6200 ;
        RECT 3303.1200 1146.5800 3304.7200 1147.0600 ;
        RECT 3303.1200 1152.0200 3304.7200 1152.5000 ;
        RECT 3303.1200 1157.4600 3304.7200 1157.9400 ;
        RECT 3303.1200 1162.9000 3304.7200 1163.3800 ;
        RECT 3303.1200 1168.3400 3304.7200 1168.8200 ;
        RECT 3303.1200 1173.7800 3304.7200 1174.2600 ;
        RECT 3365.4200 1130.2600 3368.4200 1130.7400 ;
        RECT 3365.4200 1135.7000 3368.4200 1136.1800 ;
        RECT 3365.4200 1141.1400 3368.4200 1141.6200 ;
        RECT 3365.4200 1146.5800 3368.4200 1147.0600 ;
        RECT 3365.4200 1152.0200 3368.4200 1152.5000 ;
        RECT 3365.4200 1157.4600 3368.4200 1157.9400 ;
        RECT 3365.4200 1162.9000 3368.4200 1163.3800 ;
        RECT 3365.4200 1168.3400 3368.4200 1168.8200 ;
        RECT 3365.4200 1173.7800 3368.4200 1174.2600 ;
        RECT 3303.1200 1184.6600 3304.7200 1185.1400 ;
        RECT 3303.1200 1190.1000 3304.7200 1190.5800 ;
        RECT 3303.1200 1195.5400 3304.7200 1196.0200 ;
        RECT 3303.1200 1200.9800 3304.7200 1201.4600 ;
        RECT 3303.1200 1206.4200 3304.7200 1206.9000 ;
        RECT 3303.1200 1211.8600 3304.7200 1212.3400 ;
        RECT 3303.1200 1217.3000 3304.7200 1217.7800 ;
        RECT 3303.1200 1222.7400 3304.7200 1223.2200 ;
        RECT 3303.1200 1228.1800 3304.7200 1228.6600 ;
        RECT 3365.4200 1184.6600 3368.4200 1185.1400 ;
        RECT 3365.4200 1190.1000 3368.4200 1190.5800 ;
        RECT 3365.4200 1195.5400 3368.4200 1196.0200 ;
        RECT 3365.4200 1200.9800 3368.4200 1201.4600 ;
        RECT 3365.4200 1206.4200 3368.4200 1206.9000 ;
        RECT 3365.4200 1211.8600 3368.4200 1212.3400 ;
        RECT 3365.4200 1217.3000 3368.4200 1217.7800 ;
        RECT 3365.4200 1222.7400 3368.4200 1223.2200 ;
        RECT 3365.4200 1228.1800 3368.4200 1228.6600 ;
        RECT 3303.1200 1233.6200 3304.7200 1234.1000 ;
        RECT 3303.1200 1239.0600 3304.7200 1239.5400 ;
        RECT 3303.1200 1244.5000 3304.7200 1244.9800 ;
        RECT 3303.1200 1249.9400 3304.7200 1250.4200 ;
        RECT 3303.1200 1255.3800 3304.7200 1255.8600 ;
        RECT 3303.1200 1260.8200 3304.7200 1261.3000 ;
        RECT 3303.1200 1266.2600 3304.7200 1266.7400 ;
        RECT 3303.1200 1271.7000 3304.7200 1272.1800 ;
        RECT 3303.1200 1277.1400 3304.7200 1277.6200 ;
        RECT 3303.1200 1282.5800 3304.7200 1283.0600 ;
        RECT 3365.4200 1233.6200 3368.4200 1234.1000 ;
        RECT 3365.4200 1239.0600 3368.4200 1239.5400 ;
        RECT 3365.4200 1244.5000 3368.4200 1244.9800 ;
        RECT 3365.4200 1249.9400 3368.4200 1250.4200 ;
        RECT 3365.4200 1255.3800 3368.4200 1255.8600 ;
        RECT 3365.4200 1260.8200 3368.4200 1261.3000 ;
        RECT 3365.4200 1266.2600 3368.4200 1266.7400 ;
        RECT 3365.4200 1271.7000 3368.4200 1272.1800 ;
        RECT 3365.4200 1277.1400 3368.4200 1277.6200 ;
        RECT 3365.4200 1282.5800 3368.4200 1283.0600 ;
        RECT 2.0000 1288.0200 5.0000 1288.5000 ;
        RECT 2.0000 1293.4600 5.0000 1293.9400 ;
        RECT 2.0000 1298.9000 5.0000 1299.3800 ;
        RECT 2.0000 1304.3400 5.0000 1304.8200 ;
        RECT 2.0000 1309.7800 5.0000 1310.2600 ;
        RECT 2.0000 1315.2200 5.0000 1315.7000 ;
        RECT 2.0000 1320.6600 5.0000 1321.1400 ;
        RECT 2.0000 1326.1000 5.0000 1326.5800 ;
        RECT 2.0000 1331.5400 5.0000 1332.0200 ;
        RECT 2.0000 1336.9800 5.0000 1337.4600 ;
        RECT 2.0000 1342.4200 5.0000 1342.9000 ;
        RECT 2.0000 1347.8600 5.0000 1348.3400 ;
        RECT 2.0000 1353.3000 5.0000 1353.7800 ;
        RECT 2.0000 1358.7400 5.0000 1359.2200 ;
        RECT 2.0000 1364.1800 5.0000 1364.6600 ;
        RECT 2.0000 1369.6200 5.0000 1370.1000 ;
        RECT 2.0000 1375.0600 5.0000 1375.5400 ;
        RECT 2.0000 1380.5000 5.0000 1380.9800 ;
        RECT 2.0000 1385.9400 5.0000 1386.4200 ;
        RECT 155.5200 1288.0200 157.1200 1288.5000 ;
        RECT 155.5200 1293.4600 157.1200 1293.9400 ;
        RECT 155.5200 1298.9000 157.1200 1299.3800 ;
        RECT 155.5200 1304.3400 157.1200 1304.8200 ;
        RECT 155.5200 1309.7800 157.1200 1310.2600 ;
        RECT 155.5200 1315.2200 157.1200 1315.7000 ;
        RECT 155.5200 1320.6600 157.1200 1321.1400 ;
        RECT 155.5200 1326.6100 157.1200 1328.6600 ;
        RECT 155.5200 1331.5400 157.1200 1332.0200 ;
        RECT 155.5200 1336.9800 157.1200 1337.4600 ;
        RECT 155.5200 1342.4200 157.1200 1342.9000 ;
        RECT 155.5200 1347.8600 157.1200 1348.3400 ;
        RECT 155.5200 1353.3000 157.1200 1353.7800 ;
        RECT 155.5200 1358.7400 157.1200 1359.2200 ;
        RECT 155.5200 1364.1800 157.1200 1364.6600 ;
        RECT 155.5200 1369.6200 157.1200 1370.1000 ;
        RECT 155.5200 1375.0600 157.1200 1375.5400 ;
        RECT 155.5200 1380.5000 157.1200 1380.9800 ;
        RECT 155.5200 1385.9400 157.1200 1386.4200 ;
        RECT 2.0000 1391.3800 5.0000 1391.8600 ;
        RECT 2.0000 1396.8200 5.0000 1397.3000 ;
        RECT 2.0000 1402.2600 5.0000 1402.7400 ;
        RECT 2.0000 1407.7000 5.0000 1408.1800 ;
        RECT 2.0000 1413.1400 5.0000 1413.6200 ;
        RECT 2.0000 1429.4600 5.0000 1429.9400 ;
        RECT 2.0000 1418.5800 5.0000 1419.0600 ;
        RECT 2.0000 1424.0200 5.0000 1424.5000 ;
        RECT 2.0000 1434.9000 5.0000 1435.3800 ;
        RECT 2.0000 1440.3400 5.0000 1440.8200 ;
        RECT 2.0000 1445.7800 5.0000 1446.2600 ;
        RECT 2.0000 1451.2200 5.0000 1451.7000 ;
        RECT 2.0000 1456.6600 5.0000 1457.1400 ;
        RECT 2.0000 1462.1000 5.0000 1462.5800 ;
        RECT 2.0000 1467.5400 5.0000 1468.0200 ;
        RECT 2.0000 1472.9800 5.0000 1473.4600 ;
        RECT 2.0000 1478.4200 5.0000 1478.9000 ;
        RECT 2.0000 1483.8600 5.0000 1484.3400 ;
        RECT 2.0000 1489.3000 5.0000 1489.7800 ;
        RECT 2.0000 1494.7400 5.0000 1495.2200 ;
        RECT 155.5200 1391.3800 157.1200 1391.8600 ;
        RECT 155.5200 1396.8200 157.1200 1397.3000 ;
        RECT 155.5200 1402.2600 157.1200 1402.7400 ;
        RECT 155.5200 1407.7000 157.1200 1408.1800 ;
        RECT 155.5200 1413.1400 157.1200 1413.6200 ;
        RECT 155.5200 1429.4600 157.1200 1429.9400 ;
        RECT 155.5200 1418.5800 157.1200 1419.0600 ;
        RECT 155.5200 1424.0200 157.1200 1424.5000 ;
        RECT 155.5200 1434.9000 157.1200 1435.3800 ;
        RECT 155.5200 1440.3400 157.1200 1440.8200 ;
        RECT 155.5200 1445.7800 157.1200 1446.2600 ;
        RECT 155.5200 1451.2200 157.1200 1451.7000 ;
        RECT 155.5200 1456.6600 157.1200 1457.1400 ;
        RECT 155.5200 1462.1000 157.1200 1462.5800 ;
        RECT 155.5200 1467.5400 157.1200 1468.0200 ;
        RECT 155.5200 1472.9800 157.1200 1473.4600 ;
        RECT 155.5200 1478.4200 157.1200 1478.9000 ;
        RECT 155.5200 1483.8600 157.1200 1484.3400 ;
        RECT 155.5200 1489.3000 157.1200 1489.7800 ;
        RECT 155.5200 1494.7400 157.1200 1495.2200 ;
        RECT 2.0000 1500.1800 5.0000 1500.6600 ;
        RECT 2.0000 1505.6200 5.0000 1506.1000 ;
        RECT 2.0000 1511.0600 5.0000 1511.5400 ;
        RECT 2.0000 1516.5000 5.0000 1516.9800 ;
        RECT 2.0000 1521.9400 5.0000 1522.4200 ;
        RECT 2.0000 1527.3800 5.0000 1527.8600 ;
        RECT 2.0000 1532.8200 5.0000 1533.3000 ;
        RECT 2.0000 1538.2600 5.0000 1538.7400 ;
        RECT 2.0000 1543.7000 5.0000 1544.1800 ;
        RECT 2.0000 1554.5800 5.0000 1555.0600 ;
        RECT 2.0000 1549.1400 5.0000 1549.6200 ;
        RECT 2.0000 1560.0200 5.0000 1560.5000 ;
        RECT 2.0000 1565.4600 5.0000 1565.9400 ;
        RECT 2.0000 1570.9000 5.0000 1571.3800 ;
        RECT 2.0000 1587.2200 5.0000 1587.7000 ;
        RECT 2.0000 1576.3400 5.0000 1576.8200 ;
        RECT 2.0000 1581.7800 5.0000 1582.2600 ;
        RECT 2.0000 1592.6600 5.0000 1593.1400 ;
        RECT 2.0000 1598.1000 5.0000 1598.5800 ;
        RECT 155.5200 1500.1800 157.1200 1500.6600 ;
        RECT 155.5200 1505.6200 157.1200 1506.1000 ;
        RECT 155.5200 1511.0600 157.1200 1511.5400 ;
        RECT 155.5200 1516.5000 157.1200 1516.9800 ;
        RECT 155.5200 1521.9400 157.1200 1522.4200 ;
        RECT 155.5200 1527.3800 157.1200 1527.8600 ;
        RECT 155.5200 1532.8200 157.1200 1533.3000 ;
        RECT 155.5200 1538.2600 157.1200 1538.7400 ;
        RECT 155.5200 1543.7000 157.1200 1544.1800 ;
        RECT 155.5200 1549.1400 157.1200 1549.6200 ;
        RECT 155.5200 1553.0900 157.1200 1553.5700 ;
        RECT 155.5200 1560.0200 157.1200 1560.5000 ;
        RECT 155.5200 1565.4600 157.1200 1565.9400 ;
        RECT 155.5200 1570.9000 157.1200 1571.3800 ;
        RECT 155.5200 1587.2200 157.1200 1587.7000 ;
        RECT 155.5200 1576.3400 157.1200 1576.8200 ;
        RECT 155.5200 1581.7800 157.1200 1582.2600 ;
        RECT 155.5200 1592.6600 157.1200 1593.1400 ;
        RECT 155.5200 1598.1000 157.1200 1598.5800 ;
        RECT 2.0000 1603.5400 5.0000 1604.0200 ;
        RECT 2.0000 1608.9800 5.0000 1609.4600 ;
        RECT 2.0000 1614.4200 5.0000 1614.9000 ;
        RECT 2.0000 1619.8600 5.0000 1620.3400 ;
        RECT 2.0000 1625.3000 5.0000 1625.7800 ;
        RECT 2.0000 1630.7400 5.0000 1631.2200 ;
        RECT 2.0000 1636.1800 5.0000 1636.6600 ;
        RECT 2.0000 1641.6200 5.0000 1642.1000 ;
        RECT 2.0000 1647.0600 5.0000 1647.5400 ;
        RECT 2.0000 1652.5000 5.0000 1652.9800 ;
        RECT 2.0000 1679.7000 5.0000 1680.1800 ;
        RECT 2.0000 1657.9400 5.0000 1658.4200 ;
        RECT 2.0000 1663.3800 5.0000 1663.8600 ;
        RECT 2.0000 1668.8200 5.0000 1669.3000 ;
        RECT 2.0000 1674.2600 5.0000 1674.7400 ;
        RECT 2.0000 1685.1400 5.0000 1685.6200 ;
        RECT 2.0000 1690.5800 5.0000 1691.0600 ;
        RECT 2.0000 1696.0200 5.0000 1696.5000 ;
        RECT 2.0000 1701.4600 5.0000 1701.9400 ;
        RECT 155.5200 1603.5400 157.1200 1604.0200 ;
        RECT 155.5200 1608.9800 157.1200 1609.4600 ;
        RECT 155.5200 1614.4200 157.1200 1614.9000 ;
        RECT 155.5200 1619.8600 157.1200 1620.3400 ;
        RECT 155.5200 1625.3000 157.1200 1625.7800 ;
        RECT 155.5200 1630.7400 157.1200 1631.2200 ;
        RECT 155.5200 1636.1800 157.1200 1636.6600 ;
        RECT 155.5200 1641.6200 157.1200 1642.1000 ;
        RECT 155.5200 1647.0600 157.1200 1647.5400 ;
        RECT 155.5200 1652.5000 157.1200 1652.9800 ;
        RECT 155.5200 1679.7000 157.1200 1680.1800 ;
        RECT 155.5200 1657.9400 157.1200 1658.4200 ;
        RECT 155.5200 1663.3800 157.1200 1663.8600 ;
        RECT 155.5200 1668.8200 157.1200 1669.3000 ;
        RECT 155.5200 1674.2600 157.1200 1674.7400 ;
        RECT 155.5200 1685.1400 157.1200 1685.6200 ;
        RECT 155.5200 1690.5800 157.1200 1691.0600 ;
        RECT 155.5200 1696.0200 157.1200 1696.5000 ;
        RECT 155.5200 1701.4600 157.1200 1701.9400 ;
        RECT 2.0000 1706.9000 5.0000 1707.3800 ;
        RECT 2.0000 1712.3400 5.0000 1712.8200 ;
        RECT 2.0000 1717.7800 5.0000 1718.2600 ;
        RECT 2.0000 1723.2200 5.0000 1723.7000 ;
        RECT 2.0000 1728.6600 5.0000 1729.1400 ;
        RECT 2.0000 1734.1000 5.0000 1734.5800 ;
        RECT 2.0000 1739.5400 5.0000 1740.0200 ;
        RECT 2.0000 1744.9800 5.0000 1745.4600 ;
        RECT 2.0000 1750.4200 5.0000 1750.9000 ;
        RECT 2.0000 1755.8600 5.0000 1756.3400 ;
        RECT 2.0000 1761.3000 5.0000 1761.7800 ;
        RECT 2.0000 1766.7400 5.0000 1767.2200 ;
        RECT 2.0000 1772.1800 5.0000 1772.6600 ;
        RECT 2.0000 1777.6200 5.0000 1778.1000 ;
        RECT 2.0000 1783.0600 5.0000 1783.5400 ;
        RECT 2.0000 1788.5000 5.0000 1788.9800 ;
        RECT 2.0000 1793.9400 5.0000 1794.4200 ;
        RECT 2.0000 1799.3800 5.0000 1799.8600 ;
        RECT 2.0000 1804.8200 5.0000 1805.3000 ;
        RECT 2.0000 1810.2600 5.0000 1810.7400 ;
        RECT 155.5200 1706.9000 157.1200 1707.3800 ;
        RECT 155.5200 1712.3400 157.1200 1712.8200 ;
        RECT 155.5200 1717.7800 157.1200 1718.2600 ;
        RECT 155.5200 1723.2200 157.1200 1723.7000 ;
        RECT 155.5200 1728.6600 157.1200 1729.1400 ;
        RECT 155.5200 1734.1000 157.1200 1734.5800 ;
        RECT 155.5200 1739.5400 157.1200 1740.0200 ;
        RECT 155.5200 1744.9800 157.1200 1745.4600 ;
        RECT 155.5200 1750.4200 157.1200 1750.9000 ;
        RECT 155.5200 1755.8600 157.1200 1756.3400 ;
        RECT 155.5200 1761.3000 157.1200 1761.7800 ;
        RECT 155.5200 1766.7400 157.1200 1767.2200 ;
        RECT 155.5200 1772.1800 157.1200 1772.6600 ;
        RECT 155.5200 1777.6200 157.1200 1778.1000 ;
        RECT 155.5200 1782.8900 157.1200 1783.3700 ;
        RECT 155.5200 1788.5000 157.1200 1788.9800 ;
        RECT 155.5200 1793.9400 157.1200 1794.4200 ;
        RECT 155.5200 1799.3800 157.1200 1799.8600 ;
        RECT 155.5200 1804.8200 157.1200 1805.3000 ;
        RECT 155.5200 1810.2600 157.1200 1810.7400 ;
        RECT 2.0000 1837.4600 5.0000 1837.9400 ;
        RECT 2.0000 1815.7000 5.0000 1816.1800 ;
        RECT 2.0000 1821.1400 5.0000 1821.6200 ;
        RECT 2.0000 1826.5800 5.0000 1827.0600 ;
        RECT 2.0000 1832.0200 5.0000 1832.5000 ;
        RECT 2.0000 1842.9000 5.0000 1843.3800 ;
        RECT 2.0000 1848.3400 5.0000 1848.8200 ;
        RECT 2.0000 1853.7800 5.0000 1854.2600 ;
        RECT 2.0000 1859.2200 5.0000 1859.7000 ;
        RECT 2.0000 1864.6600 5.0000 1865.1400 ;
        RECT 2.0000 1870.1000 5.0000 1870.5800 ;
        RECT 2.0000 1875.5400 5.0000 1876.0200 ;
        RECT 2.0000 1880.9800 5.0000 1881.4600 ;
        RECT 2.0000 1886.4200 5.0000 1886.9000 ;
        RECT 2.0000 1891.8600 5.0000 1892.3400 ;
        RECT 2.0000 1897.3000 5.0000 1897.7800 ;
        RECT 2.0000 1902.7400 5.0000 1903.2200 ;
        RECT 2.0000 1908.1800 5.0000 1908.6600 ;
        RECT 2.0000 1913.6200 5.0000 1914.1000 ;
        RECT 155.5200 1837.4600 157.1200 1837.9400 ;
        RECT 155.5200 1815.7000 157.1200 1816.1800 ;
        RECT 155.5200 1821.1400 157.1200 1821.6200 ;
        RECT 155.5200 1826.5800 157.1200 1827.0600 ;
        RECT 155.5200 1832.0200 157.1200 1832.5000 ;
        RECT 155.5200 1842.9000 157.1200 1843.3800 ;
        RECT 155.5200 1848.3400 157.1200 1848.8200 ;
        RECT 155.5200 1853.7800 157.1200 1854.2600 ;
        RECT 155.5200 1859.2200 157.1200 1859.7000 ;
        RECT 155.5200 1864.6600 157.1200 1865.1400 ;
        RECT 155.5200 1870.1000 157.1200 1870.5800 ;
        RECT 155.5200 1875.5400 157.1200 1876.0200 ;
        RECT 155.5200 1880.9800 157.1200 1881.4600 ;
        RECT 155.5200 1886.4200 157.1200 1886.9000 ;
        RECT 155.5200 1891.8600 157.1200 1892.3400 ;
        RECT 155.5200 1897.3000 157.1200 1897.7800 ;
        RECT 155.5200 1902.7400 157.1200 1903.2200 ;
        RECT 155.5200 1908.1800 157.1200 1908.6600 ;
        RECT 155.5200 1913.6200 157.1200 1914.1000 ;
        RECT 2.0000 1929.9400 5.0000 1930.4200 ;
        RECT 2.0000 1919.0600 5.0000 1919.5400 ;
        RECT 2.0000 1924.5000 5.0000 1924.9800 ;
        RECT 2.0000 1935.3800 5.0000 1935.8600 ;
        RECT 2.0000 1940.8200 5.0000 1941.3000 ;
        RECT 2.0000 1946.2600 5.0000 1946.7400 ;
        RECT 2.0000 1951.7000 5.0000 1952.1800 ;
        RECT 2.0000 1957.1400 5.0000 1957.6200 ;
        RECT 2.0000 1962.5800 5.0000 1963.0600 ;
        RECT 2.0000 1968.0200 5.0000 1968.5000 ;
        RECT 2.0000 1973.4600 5.0000 1973.9400 ;
        RECT 2.0000 1978.9000 5.0000 1979.3800 ;
        RECT 2.0000 1984.3400 5.0000 1984.8200 ;
        RECT 2.0000 1989.7800 5.0000 1990.2600 ;
        RECT 2.0000 1995.2200 5.0000 1995.7000 ;
        RECT 2.0000 2000.6600 5.0000 2001.1400 ;
        RECT 2.0000 2006.1000 5.0000 2006.5800 ;
        RECT 2.0000 2011.5400 5.0000 2012.0200 ;
        RECT 155.5200 1929.9400 157.1200 1930.4200 ;
        RECT 155.5200 1919.0600 157.1200 1919.5400 ;
        RECT 155.5200 1924.5000 157.1200 1924.9800 ;
        RECT 155.5200 1935.3800 157.1200 1935.8600 ;
        RECT 155.5200 1940.8200 157.1200 1941.3000 ;
        RECT 155.5200 1946.2600 157.1200 1946.7400 ;
        RECT 155.5200 1951.7000 157.1200 1952.1800 ;
        RECT 155.5200 1957.1400 157.1200 1957.6200 ;
        RECT 155.5200 1962.5800 157.1200 1963.0600 ;
        RECT 155.5200 1968.0200 157.1200 1968.5000 ;
        RECT 155.5200 1973.4600 157.1200 1973.9400 ;
        RECT 155.5200 1978.9000 157.1200 1979.3800 ;
        RECT 155.5200 1984.3400 157.1200 1984.8200 ;
        RECT 155.5200 1989.7800 157.1200 1990.2600 ;
        RECT 155.5200 1995.2200 157.1200 1995.7000 ;
        RECT 155.5200 2000.6600 157.1200 2001.1400 ;
        RECT 155.5200 2006.1000 157.1200 2006.5800 ;
        RECT 155.5200 2011.5400 157.1200 2012.0200 ;
        RECT 2.0000 2022.4200 5.0000 2022.9000 ;
        RECT 2.0000 2027.8600 5.0000 2028.3400 ;
        RECT 2.0000 2033.3000 5.0000 2033.7800 ;
        RECT 2.0000 2038.7400 5.0000 2039.2200 ;
        RECT 2.0000 2044.1800 5.0000 2044.6600 ;
        RECT 2.0000 2049.6200 5.0000 2050.1000 ;
        RECT 2.0000 2055.0600 5.0000 2055.5400 ;
        RECT 2.0000 2060.5000 5.0000 2060.9800 ;
        RECT 2.0000 2065.9400 5.0000 2066.4200 ;
        RECT 2.0000 2071.3800 5.0000 2071.8600 ;
        RECT 2.0000 2087.7000 5.0000 2088.1800 ;
        RECT 2.0000 2076.8200 5.0000 2077.3000 ;
        RECT 2.0000 2082.2600 5.0000 2082.7400 ;
        RECT 2.0000 2093.1400 5.0000 2093.6200 ;
        RECT 2.0000 2098.5800 5.0000 2099.0600 ;
        RECT 2.0000 2104.0200 5.0000 2104.5000 ;
        RECT 2.0000 2109.4600 5.0000 2109.9400 ;
        RECT 2.0000 2114.9000 5.0000 2115.3800 ;
        RECT 2.0000 2120.3400 5.0000 2120.8200 ;
        RECT 2.0000 2125.7800 5.0000 2126.2600 ;
        RECT 1015.5800 1341.2800 1017.1800 1341.7600 ;
        RECT 1015.5800 1570.9200 1017.1800 1571.4000 ;
        RECT 1063.2600 1543.6900 1064.8600 1546.2400 ;
        RECT 1075.8200 1570.9200 1077.4200 1571.4000 ;
        RECT 1063.2600 1566.6300 1064.8600 1568.3300 ;
        RECT 1295.9000 1341.0200 1297.5000 1341.5000 ;
        RECT 1516.1200 1341.0200 1517.7200 1341.5000 ;
        RECT 1283.3400 1543.3300 1285.0800 1546.2400 ;
        RECT 1295.9000 1570.6600 1297.5000 1571.1400 ;
        RECT 1283.3400 1556.4400 1285.0800 1558.3000 ;
        RECT 1283.3400 1566.4700 1285.0800 1568.3300 ;
        RECT 1516.1200 1570.6600 1517.7200 1571.1400 ;
        RECT 1015.5800 1800.5600 1017.1800 1801.0400 ;
        RECT 963.1200 1973.4600 964.7200 1973.9400 ;
        RECT 963.1200 1978.9000 964.7200 1979.3800 ;
        RECT 963.1200 1984.3400 964.7200 1984.8200 ;
        RECT 963.1200 1989.7800 964.7200 1990.2600 ;
        RECT 963.1200 1995.2200 964.7200 1995.7000 ;
        RECT 963.1200 2000.6600 964.7200 2001.1400 ;
        RECT 963.1200 2006.1000 964.7200 2006.5800 ;
        RECT 963.1200 2011.5400 964.7200 2012.0200 ;
        RECT 1005.5200 1973.4600 1007.1200 1973.9400 ;
        RECT 1005.5200 1978.9000 1007.1200 1979.3800 ;
        RECT 1005.5200 1984.3400 1007.1200 1984.8200 ;
        RECT 1005.5200 1989.7800 1007.1200 1990.2600 ;
        RECT 1005.5200 1995.2200 1007.1200 1995.7000 ;
        RECT 1005.5200 2000.6600 1007.1200 2001.1400 ;
        RECT 1005.5200 2007.2900 1007.1200 2007.7700 ;
        RECT 1005.5200 2011.5400 1007.1200 2012.0200 ;
        RECT 1005.5200 2033.3000 1007.1200 2033.7800 ;
        RECT 1005.5200 2027.8600 1007.1200 2028.3400 ;
        RECT 1005.5200 2022.4200 1007.1200 2022.9000 ;
        RECT 1015.5800 2030.2000 1017.1800 2030.6800 ;
        RECT 1005.5200 2038.7400 1007.1200 2039.2200 ;
        RECT 1005.5200 2044.1800 1007.1200 2044.6600 ;
        RECT 1005.5200 2049.6200 1007.1200 2050.1000 ;
        RECT 1005.5200 2055.0600 1007.1200 2055.5400 ;
        RECT 1005.5200 2060.5000 1007.1200 2060.9800 ;
        RECT 1005.5200 2065.9400 1007.1200 2066.4200 ;
        RECT 1005.5200 2071.3800 1007.1200 2071.8600 ;
        RECT 1005.5200 2087.7000 1007.1200 2088.1800 ;
        RECT 1005.5200 2076.8200 1007.1200 2077.3000 ;
        RECT 1005.5200 2082.2600 1007.1200 2082.7400 ;
        RECT 1005.5200 2093.1400 1007.1200 2093.6200 ;
        RECT 1005.5200 2098.5800 1007.1200 2099.0600 ;
        RECT 1005.5200 2104.0200 1007.1200 2104.5000 ;
        RECT 1005.5200 2109.4600 1007.1200 2109.9400 ;
        RECT 1005.5200 2114.9000 1007.1200 2115.3800 ;
        RECT 1005.5200 2120.3400 1007.1200 2120.8200 ;
        RECT 1005.5200 2125.7800 1007.1200 2126.2600 ;
        RECT 1063.2600 2002.9700 1064.8600 2005.5200 ;
        RECT 1063.2600 2025.9100 1064.8600 2027.6100 ;
        RECT 1075.8200 2030.2000 1077.4200 2030.6800 ;
        RECT 1295.9000 1800.3000 1297.5000 1800.7800 ;
        RECT 1516.1200 1800.3000 1517.7200 1800.7800 ;
        RECT 1283.3400 2015.7200 1285.0800 2017.5800 ;
        RECT 1283.3400 2002.6100 1285.0800 2005.5200 ;
        RECT 1283.3400 2025.7500 1285.0800 2027.6100 ;
        RECT 1295.9000 2029.9400 1297.5000 2030.4200 ;
        RECT 1516.1200 2029.9400 1517.7200 2030.4200 ;
        RECT 2.0000 2337.9400 5.0000 2338.4200 ;
        RECT 2.0000 2131.2200 5.0000 2131.7000 ;
        RECT 2.0000 2136.6600 5.0000 2137.1400 ;
        RECT 2.0000 2142.1000 5.0000 2142.5800 ;
        RECT 2.0000 2147.5400 5.0000 2148.0200 ;
        RECT 2.0000 2152.9800 5.0000 2153.4600 ;
        RECT 2.0000 2158.4200 5.0000 2158.9000 ;
        RECT 2.0000 2163.8600 5.0000 2164.3400 ;
        RECT 2.0000 2169.3000 5.0000 2169.7800 ;
        RECT 2.0000 2174.7400 5.0000 2175.2200 ;
        RECT 2.0000 2180.1800 5.0000 2180.6600 ;
        RECT 2.0000 2185.6200 5.0000 2186.1000 ;
        RECT 2.0000 2191.0600 5.0000 2191.5400 ;
        RECT 2.0000 2196.5000 5.0000 2196.9800 ;
        RECT 2.0000 2201.9400 5.0000 2202.4200 ;
        RECT 2.0000 2207.3800 5.0000 2207.8600 ;
        RECT 2.0000 2212.8200 5.0000 2213.3000 ;
        RECT 2.0000 2218.2600 5.0000 2218.7400 ;
        RECT 2.0000 2223.7000 5.0000 2224.1800 ;
        RECT 2.0000 2229.1400 5.0000 2229.6200 ;
        RECT 2.0000 2245.4600 5.0000 2247.2200 ;
        RECT 2.0000 2234.5800 5.0000 2235.0600 ;
        RECT 2.0000 2240.0200 5.0000 2240.5000 ;
        RECT 2.0000 2250.9000 5.0000 2251.3800 ;
        RECT 2.0000 2256.3400 5.0000 2256.8200 ;
        RECT 2.0000 2261.7800 5.0000 2262.2600 ;
        RECT 2.0000 2267.2200 5.0000 2267.7000 ;
        RECT 2.0000 2272.6600 5.0000 2273.1400 ;
        RECT 2.0000 2278.1000 5.0000 2278.5800 ;
        RECT 2.0000 2283.5400 5.0000 2284.0200 ;
        RECT 2.0000 2288.9800 5.0000 2289.4600 ;
        RECT 2.0000 2294.4200 5.0000 2294.9000 ;
        RECT 2.0000 2299.8600 5.0000 2300.3400 ;
        RECT 2.0000 2305.3000 5.0000 2305.7800 ;
        RECT 2.0000 2310.7400 5.0000 2311.2200 ;
        RECT 2.0000 2316.1800 5.0000 2316.6600 ;
        RECT 2.0000 2321.6200 5.0000 2322.1000 ;
        RECT 2.0000 2327.0600 5.0000 2327.5400 ;
        RECT 2.0000 2332.5000 5.0000 2332.9800 ;
        RECT 2.0000 2343.3800 5.0000 2343.8600 ;
        RECT 2.0000 2348.8200 5.0000 2349.3000 ;
        RECT 2.0000 2354.2600 5.0000 2354.7400 ;
        RECT 2.0000 2359.7000 5.0000 2360.1800 ;
        RECT 2.0000 2365.1400 5.0000 2365.6200 ;
        RECT 2.0000 2370.5800 5.0000 2371.0600 ;
        RECT 2.0000 2376.0200 5.0000 2376.5000 ;
        RECT 2.0000 2381.4600 5.0000 2381.9400 ;
        RECT 2.0000 2386.9000 5.0000 2387.3800 ;
        RECT 2.0000 2392.3400 5.0000 2392.8200 ;
        RECT 2.0000 2397.7800 5.0000 2398.2600 ;
        RECT 2.0000 2403.2200 5.0000 2403.7000 ;
        RECT 2.0000 2408.6600 5.0000 2409.1400 ;
        RECT 2.0000 2414.1000 5.0000 2414.5800 ;
        RECT 2.0000 2419.5400 5.0000 2420.0200 ;
        RECT 2.0000 2424.9800 5.0000 2425.4600 ;
        RECT 2.0000 2430.4200 5.0000 2430.9000 ;
        RECT 2.0000 2435.8600 5.0000 2436.3400 ;
        RECT 2.0000 2441.3000 5.0000 2441.7800 ;
        RECT 2.0000 2495.7000 5.0000 2496.1800 ;
        RECT 2.0000 2446.7400 5.0000 2447.2200 ;
        RECT 2.0000 2452.1800 5.0000 2452.6600 ;
        RECT 2.0000 2457.6200 5.0000 2458.1000 ;
        RECT 2.0000 2463.0600 5.0000 2463.5400 ;
        RECT 2.0000 2468.5000 5.0000 2468.9800 ;
        RECT 2.0000 2473.9400 5.0000 2474.4200 ;
        RECT 2.0000 2479.3800 5.0000 2479.8600 ;
        RECT 2.0000 2484.8200 5.0000 2485.3000 ;
        RECT 2.0000 2490.2600 5.0000 2490.7400 ;
        RECT 2.0000 2501.1400 5.0000 2501.6200 ;
        RECT 2.0000 2506.5800 5.0000 2507.0600 ;
        RECT 2.0000 2512.0200 5.0000 2512.5000 ;
        RECT 2.0000 2517.4600 5.0000 2517.9400 ;
        RECT 2.0000 2522.9000 5.0000 2523.3800 ;
        RECT 2.0000 2528.3400 5.0000 2528.8200 ;
        RECT 2.0000 2533.7800 5.0000 2534.2600 ;
        RECT 2.0000 2539.2200 5.0000 2539.7000 ;
        RECT 2.0000 2544.6600 5.0000 2545.1400 ;
        RECT 2.0000 2550.1000 5.0000 2550.5800 ;
        RECT 2.0000 2555.5400 5.0000 2556.0200 ;
        RECT 1005.5200 2337.9400 1007.1200 2338.4200 ;
        RECT 1005.5200 2232.6100 1007.1200 2234.5500 ;
        RECT 1005.5200 2131.2200 1007.1200 2131.7000 ;
        RECT 1005.5200 2136.6600 1007.1200 2137.1400 ;
        RECT 1005.5200 2142.1000 1007.1200 2142.5800 ;
        RECT 1005.5200 2147.5400 1007.1200 2148.0200 ;
        RECT 1005.5200 2152.9800 1007.1200 2153.4600 ;
        RECT 1005.5200 2158.4200 1007.1200 2158.9000 ;
        RECT 1005.5200 2163.8600 1007.1200 2164.3400 ;
        RECT 1005.5200 2169.3000 1007.1200 2169.7800 ;
        RECT 1005.5200 2174.7400 1007.1200 2175.2200 ;
        RECT 1005.5200 2180.1800 1007.1200 2180.6600 ;
        RECT 1005.5200 2185.6200 1007.1200 2186.1000 ;
        RECT 1005.5200 2191.0600 1007.1200 2191.5400 ;
        RECT 1005.5200 2196.5000 1007.1200 2196.9800 ;
        RECT 1005.5200 2201.9400 1007.1200 2202.4200 ;
        RECT 1005.5200 2207.3800 1007.1200 2207.8600 ;
        RECT 1005.5200 2212.8200 1007.1200 2213.3000 ;
        RECT 1005.5200 2218.2600 1007.1200 2218.7400 ;
        RECT 1005.5200 2223.7000 1007.1200 2224.1800 ;
        RECT 1005.5200 2229.1400 1007.1200 2229.6200 ;
        RECT 1005.5200 2245.4600 1007.1200 2247.2200 ;
        RECT 1005.5200 2240.0200 1007.1200 2240.5000 ;
        RECT 1005.5200 2250.9000 1007.1200 2251.3800 ;
        RECT 1005.5200 2261.7800 1007.1200 2262.2600 ;
        RECT 1005.5200 2267.2200 1007.1200 2267.7000 ;
        RECT 1015.5800 2259.8400 1017.1800 2260.3200 ;
        RECT 1005.5200 2272.6600 1007.1200 2273.1400 ;
        RECT 1005.5200 2278.1000 1007.1200 2278.5800 ;
        RECT 1005.5200 2283.5400 1007.1200 2284.0200 ;
        RECT 1005.5200 2288.9800 1007.1200 2289.4600 ;
        RECT 1005.5200 2294.4200 1007.1200 2294.9000 ;
        RECT 1005.5200 2299.8600 1007.1200 2300.3400 ;
        RECT 1005.5200 2305.3000 1007.1200 2305.7800 ;
        RECT 1005.5200 2310.7400 1007.1200 2311.2200 ;
        RECT 1005.5200 2316.1800 1007.1200 2316.6600 ;
        RECT 1005.5200 2321.6200 1007.1200 2322.1000 ;
        RECT 1005.5200 2327.0600 1007.1200 2327.5400 ;
        RECT 1005.5200 2332.5000 1007.1200 2332.9800 ;
        RECT 1053.2000 2495.7000 1054.8000 2496.1800 ;
        RECT 1053.2000 2484.8200 1054.8000 2485.3000 ;
        RECT 1053.2000 2490.2600 1054.8000 2490.7400 ;
        RECT 1053.2000 2501.1400 1054.8000 2501.6200 ;
        RECT 1053.2000 2506.5800 1054.8000 2507.0600 ;
        RECT 1053.2000 2512.0200 1054.8000 2512.5000 ;
        RECT 1053.2000 2517.4600 1054.8000 2517.9400 ;
        RECT 1053.2000 2533.7800 1054.8000 2534.2600 ;
        RECT 1053.2000 2528.3400 1054.8000 2528.8200 ;
        RECT 1053.2000 2522.9000 1054.8000 2523.3800 ;
        RECT 1053.2000 2544.6600 1054.8000 2545.1400 ;
        RECT 1053.2000 2539.2200 1054.8000 2539.7000 ;
        RECT 1005.5200 2343.3800 1007.1200 2343.8600 ;
        RECT 1005.5200 2348.8200 1007.1200 2349.3000 ;
        RECT 1005.5200 2354.2600 1007.1200 2354.7400 ;
        RECT 1005.5200 2359.7000 1007.1200 2360.1800 ;
        RECT 1005.5200 2365.1400 1007.1200 2365.6200 ;
        RECT 1005.5200 2370.5800 1007.1200 2371.0600 ;
        RECT 1005.5200 2376.0200 1007.1200 2376.5000 ;
        RECT 1005.5200 2381.4600 1007.1200 2381.9400 ;
        RECT 1005.5200 2386.9000 1007.1200 2387.3800 ;
        RECT 1005.5200 2392.3400 1007.1200 2392.8200 ;
        RECT 1005.5200 2397.7800 1007.1200 2398.2600 ;
        RECT 1005.5200 2403.2200 1007.1200 2403.7000 ;
        RECT 1005.5200 2408.6600 1007.1200 2409.1400 ;
        RECT 1005.5200 2414.1000 1007.1200 2414.5800 ;
        RECT 1005.5200 2419.5400 1007.1200 2420.0200 ;
        RECT 1005.5200 2424.9800 1007.1200 2425.4600 ;
        RECT 1005.5200 2430.4200 1007.1200 2430.9000 ;
        RECT 1005.5200 2435.8600 1007.1200 2436.3400 ;
        RECT 1005.5200 2441.3000 1007.1200 2441.7800 ;
        RECT 1005.5200 2495.7000 1007.1200 2496.1800 ;
        RECT 1015.5800 2495.7000 1017.1800 2496.1800 ;
        RECT 1005.5200 2446.7400 1007.1200 2447.2200 ;
        RECT 1005.5200 2452.1800 1007.1200 2452.6600 ;
        RECT 1005.5200 2457.6200 1007.1200 2458.1000 ;
        RECT 1005.5200 2468.5000 1007.1200 2468.9800 ;
        RECT 1005.5200 2473.9400 1007.1200 2474.4200 ;
        RECT 1005.5200 2479.3800 1007.1200 2479.8600 ;
        RECT 1005.5200 2484.8200 1007.1200 2485.3000 ;
        RECT 1005.5200 2490.2600 1007.1200 2490.7400 ;
        RECT 1015.5800 2484.8200 1017.1800 2485.3000 ;
        RECT 1015.5800 2490.2600 1017.1800 2490.7400 ;
        RECT 1005.5200 2501.1400 1007.1200 2501.6200 ;
        RECT 1005.5200 2506.5800 1007.1200 2507.0600 ;
        RECT 1015.5800 2501.1400 1017.1800 2501.6200 ;
        RECT 1015.5800 2506.5800 1017.1800 2507.0600 ;
        RECT 1005.5200 2512.0200 1007.1200 2512.5000 ;
        RECT 1005.5200 2517.4600 1007.1200 2517.9400 ;
        RECT 1015.5800 2512.0200 1017.1800 2512.5000 ;
        RECT 1015.5800 2517.4600 1017.1800 2517.9400 ;
        RECT 1005.5200 2522.9000 1007.1200 2523.3800 ;
        RECT 1005.5200 2528.3400 1007.1200 2528.8200 ;
        RECT 1005.5200 2533.7800 1007.1200 2534.2600 ;
        RECT 1015.5800 2522.9000 1017.1800 2523.3800 ;
        RECT 1015.5800 2528.3400 1017.1800 2528.8200 ;
        RECT 1015.5800 2533.7800 1017.1800 2534.2600 ;
        RECT 1005.5200 2539.2200 1007.1200 2539.7000 ;
        RECT 1005.5200 2544.6600 1007.1200 2545.1400 ;
        RECT 1015.5800 2539.2200 1017.1800 2539.7000 ;
        RECT 1015.5800 2544.6600 1017.1800 2545.1400 ;
        RECT 1063.2600 2495.7000 1064.8600 2496.1800 ;
        RECT 1063.2600 2462.2500 1064.8600 2464.8000 ;
        RECT 1063.2600 2483.5700 1064.8600 2485.3000 ;
        RECT 1063.2600 2490.2600 1064.8600 2490.7400 ;
        RECT 1063.2600 2501.1400 1064.8600 2501.6200 ;
        RECT 1063.2600 2506.5800 1064.8600 2507.0600 ;
        RECT 1063.2600 2512.0200 1064.8600 2512.5000 ;
        RECT 1063.2600 2517.4600 1064.8600 2517.9400 ;
        RECT 1063.2600 2522.9000 1064.8600 2523.3800 ;
        RECT 1063.2600 2528.3400 1064.8600 2528.8200 ;
        RECT 1063.2600 2533.7800 1064.8600 2534.2600 ;
        RECT 1075.5800 2522.9000 1077.1800 2523.3800 ;
        RECT 1075.5800 2528.3400 1077.1800 2528.8200 ;
        RECT 1075.5800 2533.7800 1077.1800 2534.2600 ;
        RECT 1063.2600 2539.2200 1064.8600 2539.7000 ;
        RECT 1063.2600 2544.6600 1064.8600 2545.1400 ;
        RECT 1075.5800 2539.2200 1077.1800 2539.7000 ;
        RECT 1075.5800 2544.6600 1077.1800 2545.1400 ;
        RECT 1295.9000 2259.5800 1297.5000 2260.0600 ;
        RECT 1516.1200 2259.5800 1517.7200 2260.0600 ;
        RECT 1283.3400 2461.8900 1285.0800 2464.8000 ;
        RECT 1273.2800 2486.5000 1274.8800 2486.9800 ;
        RECT 1273.2800 2522.9000 1274.8800 2523.3800 ;
        RECT 1273.2800 2528.3400 1274.8800 2528.8200 ;
        RECT 1273.2800 2533.7800 1274.8800 2534.2600 ;
        RECT 1283.3400 2522.9000 1285.0800 2523.3800 ;
        RECT 1283.3400 2528.3400 1285.0800 2528.8200 ;
        RECT 1283.3400 2533.7800 1285.0800 2534.2600 ;
        RECT 1273.2800 2539.2200 1274.8800 2539.7000 ;
        RECT 1273.2800 2544.6600 1274.8800 2545.1400 ;
        RECT 1283.3400 2539.2200 1285.0800 2539.7000 ;
        RECT 1283.3400 2544.6600 1285.0800 2545.1400 ;
        RECT 1295.8000 2522.9000 1297.4000 2523.3800 ;
        RECT 1295.8000 2528.3400 1297.4000 2528.8200 ;
        RECT 1295.8000 2533.7800 1297.4000 2534.2600 ;
        RECT 1295.8000 2539.2200 1297.4000 2539.7000 ;
        RECT 1295.8000 2544.6600 1297.4000 2545.1400 ;
        RECT 1493.5000 2486.5000 1495.1000 2486.9800 ;
        RECT 1493.5000 2522.9000 1495.1000 2523.3800 ;
        RECT 1493.5000 2528.3400 1495.1000 2528.8200 ;
        RECT 1493.5000 2533.7800 1495.1000 2534.2600 ;
        RECT 1493.5000 2539.2200 1495.1000 2539.7000 ;
        RECT 1493.5000 2544.6600 1495.1000 2545.1400 ;
        RECT 1503.5600 2522.9000 1505.1600 2523.3800 ;
        RECT 1503.5600 2528.3400 1505.1600 2528.8200 ;
        RECT 1503.5600 2533.7800 1505.1600 2534.2600 ;
        RECT 1516.0200 2522.9000 1517.6200 2523.3800 ;
        RECT 1516.0200 2528.3400 1517.6200 2528.8200 ;
        RECT 1516.0200 2533.7800 1517.6200 2534.2600 ;
        RECT 1503.5600 2539.2200 1505.1600 2539.7000 ;
        RECT 1503.5600 2544.6600 1505.1600 2545.1400 ;
        RECT 1516.0200 2539.2200 1517.6200 2539.7000 ;
        RECT 1516.0200 2544.6600 1517.6200 2545.1400 ;
        RECT 1053.2000 2550.1000 1054.8000 2550.5800 ;
        RECT 1053.2000 2555.5400 1054.8000 2556.0200 ;
        RECT 1005.5200 2550.1000 1007.1200 2550.5800 ;
        RECT 1005.5200 2555.5400 1007.1200 2556.0200 ;
        RECT 1015.5800 2550.1000 1017.1800 2550.5800 ;
        RECT 1015.5800 2555.5400 1017.1800 2556.0200 ;
        RECT 1063.2600 2550.1000 1064.8600 2550.5800 ;
        RECT 1063.2600 2555.5400 1064.8600 2556.0200 ;
        RECT 1075.5800 2550.1000 1077.1800 2550.5800 ;
        RECT 1075.5800 2555.5400 1077.1800 2556.0200 ;
        RECT 1273.2800 2550.1000 1274.8800 2550.5800 ;
        RECT 1273.2800 2555.5400 1274.8800 2556.0200 ;
        RECT 1283.3400 2550.1000 1285.0800 2550.5800 ;
        RECT 1283.3400 2555.5400 1285.0800 2556.0200 ;
        RECT 1295.8000 2550.1000 1297.4000 2550.5800 ;
        RECT 1295.8000 2555.5400 1297.4000 2556.0200 ;
        RECT 1493.5000 2550.1000 1495.1000 2550.5800 ;
        RECT 1493.5000 2555.5400 1495.1000 2556.0200 ;
        RECT 1503.5600 2550.1000 1505.1600 2550.5800 ;
        RECT 1503.5600 2555.5400 1505.1600 2556.0200 ;
        RECT 1516.0200 2550.1000 1517.6200 2550.5800 ;
        RECT 1516.0200 2555.5400 1517.6200 2556.0200 ;
        RECT 1736.3400 1341.0200 1737.9400 1341.5000 ;
        RECT 1736.3400 1570.6600 1737.9400 1571.1400 ;
        RECT 1944.0000 1543.3300 1945.6000 1545.9800 ;
        RECT 1956.5600 1570.6600 1958.1600 1571.1400 ;
        RECT 2176.7800 1341.0200 2178.3800 1341.5000 ;
        RECT 2434.4200 1341.0200 2436.0200 1341.5000 ;
        RECT 2164.2200 1543.3300 2165.8200 1545.9800 ;
        RECT 2176.7800 1570.6600 2178.3800 1571.1400 ;
        RECT 2434.4200 1570.6600 2436.0200 1571.1400 ;
        RECT 1736.3400 1800.3000 1737.9400 1800.7800 ;
        RECT 1736.3400 2029.9400 1737.9400 2030.4200 ;
        RECT 1944.0000 2002.6100 1945.6000 2005.2600 ;
        RECT 1956.5600 2029.9400 1958.1600 2030.4200 ;
        RECT 2176.7800 1800.3000 2178.3800 1800.7800 ;
        RECT 2434.4200 1800.3000 2436.0200 1800.7800 ;
        RECT 2164.2200 2002.6100 2165.8200 2005.2600 ;
        RECT 2176.7800 2029.9400 2178.3800 2030.4200 ;
        RECT 2444.5800 1973.4600 2446.1800 1973.9400 ;
        RECT 2444.5800 1978.9000 2446.1800 1979.3800 ;
        RECT 2444.5800 1984.3400 2446.1800 1984.8200 ;
        RECT 2444.5800 1989.7800 2446.1800 1990.2600 ;
        RECT 2444.5800 1995.2200 2446.1800 1995.7000 ;
        RECT 2444.5800 2000.6600 2446.1800 2001.1400 ;
        RECT 2444.5800 2007.2900 2446.1800 2007.7700 ;
        RECT 2444.5800 2011.5400 2446.1800 2012.0200 ;
        RECT 2444.5800 2015.7200 2446.1800 2017.4600 ;
        RECT 2495.5200 1973.4600 2497.1200 1973.9400 ;
        RECT 2495.5200 1978.9000 2497.1200 1979.3800 ;
        RECT 2495.5200 1984.3400 2497.1200 1984.8200 ;
        RECT 2495.5200 1989.7800 2497.1200 1990.2600 ;
        RECT 2495.5200 1995.2200 2497.1200 1995.7000 ;
        RECT 2495.5200 2000.6600 2497.1200 2001.1400 ;
        RECT 2495.5200 2006.1000 2497.1200 2006.5800 ;
        RECT 2495.5200 2011.5400 2497.1200 2012.0200 ;
        RECT 2495.5200 2016.9800 2497.1200 2017.4600 ;
        RECT 2434.4200 2029.9400 2436.0200 2030.4200 ;
        RECT 2444.5800 2022.2500 2446.1800 2022.7300 ;
        RECT 2444.5800 2027.8600 2446.1800 2028.3400 ;
        RECT 2444.5800 2033.3000 2446.1800 2033.7800 ;
        RECT 2444.5800 2038.7400 2446.1800 2039.2200 ;
        RECT 2444.5800 2044.1800 2446.1800 2044.6600 ;
        RECT 2444.5800 2049.6200 2446.1800 2050.1000 ;
        RECT 2444.5800 2055.0600 2446.1800 2055.5400 ;
        RECT 2444.5800 2060.5000 2446.1800 2060.9800 ;
        RECT 2444.5800 2065.9400 2446.1800 2066.4200 ;
        RECT 2444.5800 2071.3800 2446.1800 2071.8600 ;
        RECT 2495.5200 2022.4200 2497.1200 2022.9000 ;
        RECT 2495.5200 2027.8600 2497.1200 2028.3400 ;
        RECT 2495.5200 2033.3000 2497.1200 2033.7800 ;
        RECT 2495.5200 2038.7400 2497.1200 2039.2200 ;
        RECT 2495.5200 2044.1800 2497.1200 2044.6600 ;
        RECT 2495.5200 2049.6200 2497.1200 2050.1000 ;
        RECT 2495.5200 2055.0600 2497.1200 2055.5400 ;
        RECT 2495.5200 2060.5000 2497.1200 2060.9800 ;
        RECT 2495.5200 2065.9400 2497.1200 2066.4200 ;
        RECT 2495.5200 2071.3800 2497.1200 2071.8600 ;
        RECT 2444.5800 2087.7000 2446.1800 2088.1800 ;
        RECT 2444.5800 2076.8200 2446.1800 2077.3000 ;
        RECT 2444.5800 2082.2600 2446.1800 2082.7400 ;
        RECT 2444.5800 2093.1400 2446.1800 2093.6200 ;
        RECT 2444.5800 2098.5800 2446.1800 2099.0600 ;
        RECT 2444.5800 2104.0200 2446.1800 2104.5000 ;
        RECT 2444.5800 2109.4600 2446.1800 2109.9400 ;
        RECT 2444.5800 2114.9000 2446.1800 2115.3800 ;
        RECT 2444.5800 2120.3400 2446.1800 2120.8200 ;
        RECT 2444.5800 2125.7800 2446.1800 2126.2600 ;
        RECT 2495.5200 2087.7000 2497.1200 2088.1800 ;
        RECT 2495.5200 2076.8200 2497.1200 2077.3000 ;
        RECT 2495.5200 2082.2600 2497.1200 2082.7400 ;
        RECT 2495.5200 2093.1400 2497.1200 2093.6200 ;
        RECT 2495.5200 2098.5800 2497.1200 2099.0600 ;
        RECT 2495.5200 2104.0200 2497.1200 2104.5000 ;
        RECT 2495.5200 2109.4600 2497.1200 2109.9400 ;
        RECT 2495.5200 2114.9000 2497.1200 2115.3800 ;
        RECT 2495.5200 2120.3400 2497.1200 2120.8200 ;
        RECT 2495.5200 2125.7800 2497.1200 2126.2600 ;
        RECT 3303.1200 1288.0200 3304.7200 1288.5000 ;
        RECT 3303.1200 1293.4600 3304.7200 1293.9400 ;
        RECT 3303.1200 1298.9000 3304.7200 1299.3800 ;
        RECT 3303.1200 1304.3400 3304.7200 1304.8200 ;
        RECT 3303.1200 1309.7800 3304.7200 1310.2600 ;
        RECT 3303.1200 1315.2200 3304.7200 1315.7000 ;
        RECT 3303.1200 1320.6600 3304.7200 1321.1400 ;
        RECT 3303.1200 1326.1000 3304.7200 1326.5800 ;
        RECT 3303.1200 1331.5400 3304.7200 1332.0200 ;
        RECT 3303.1200 1336.9800 3304.7200 1337.4600 ;
        RECT 3365.4200 1288.0200 3368.4200 1288.5000 ;
        RECT 3365.4200 1293.4600 3368.4200 1293.9400 ;
        RECT 3365.4200 1298.9000 3368.4200 1299.3800 ;
        RECT 3365.4200 1304.3400 3368.4200 1304.8200 ;
        RECT 3365.4200 1309.7800 3368.4200 1310.2600 ;
        RECT 3365.4200 1315.2200 3368.4200 1315.7000 ;
        RECT 3365.4200 1320.6600 3368.4200 1321.1400 ;
        RECT 3365.4200 1326.1000 3368.4200 1326.5800 ;
        RECT 3365.4200 1331.5400 3368.4200 1332.0200 ;
        RECT 3365.4200 1336.9800 3368.4200 1337.4600 ;
        RECT 3303.1200 1342.4200 3304.7200 1342.9000 ;
        RECT 3303.1200 1347.8600 3304.7200 1348.3400 ;
        RECT 3303.1200 1353.3000 3304.7200 1353.7800 ;
        RECT 3303.1200 1358.7400 3304.7200 1359.2200 ;
        RECT 3303.1200 1364.1800 3304.7200 1364.6600 ;
        RECT 3303.1200 1369.6200 3304.7200 1370.1000 ;
        RECT 3303.1200 1375.0600 3304.7200 1375.5400 ;
        RECT 3303.1200 1380.5000 3304.7200 1380.9800 ;
        RECT 3303.1200 1385.9400 3304.7200 1386.4200 ;
        RECT 3365.4200 1342.4200 3368.4200 1342.9000 ;
        RECT 3365.4200 1347.8600 3368.4200 1348.3400 ;
        RECT 3365.4200 1353.3000 3368.4200 1353.7800 ;
        RECT 3365.4200 1358.7400 3368.4200 1359.2200 ;
        RECT 3365.4200 1364.1800 3368.4200 1364.6600 ;
        RECT 3365.4200 1369.6200 3368.4200 1370.1000 ;
        RECT 3365.4200 1375.0600 3368.4200 1375.5400 ;
        RECT 3365.4200 1380.5000 3368.4200 1380.9800 ;
        RECT 3365.4200 1385.9400 3368.4200 1386.4200 ;
        RECT 3303.1200 1391.3800 3304.7200 1391.8600 ;
        RECT 3303.1200 1396.8200 3304.7200 1397.3000 ;
        RECT 3303.1200 1402.2600 3304.7200 1402.7400 ;
        RECT 3303.1200 1407.7000 3304.7200 1408.1800 ;
        RECT 3303.1200 1413.1400 3304.7200 1413.6200 ;
        RECT 3303.1200 1429.4600 3304.7200 1429.9400 ;
        RECT 3303.1200 1418.5800 3304.7200 1419.0600 ;
        RECT 3303.1200 1424.0200 3304.7200 1424.5000 ;
        RECT 3303.1200 1434.9000 3304.7200 1435.3800 ;
        RECT 3303.1200 1440.3400 3304.7200 1440.8200 ;
        RECT 3365.4200 1391.3800 3368.4200 1391.8600 ;
        RECT 3365.4200 1396.8200 3368.4200 1397.3000 ;
        RECT 3365.4200 1402.2600 3368.4200 1402.7400 ;
        RECT 3365.4200 1407.7000 3368.4200 1408.1800 ;
        RECT 3365.4200 1413.1400 3368.4200 1413.6200 ;
        RECT 3365.4200 1429.4600 3368.4200 1429.9400 ;
        RECT 3365.4200 1418.5800 3368.4200 1419.0600 ;
        RECT 3365.4200 1424.0200 3368.4200 1424.5000 ;
        RECT 3365.4200 1434.9000 3368.4200 1435.3800 ;
        RECT 3365.4200 1440.3400 3368.4200 1440.8200 ;
        RECT 3303.1200 1445.7800 3304.7200 1446.2600 ;
        RECT 3303.1200 1451.2200 3304.7200 1451.7000 ;
        RECT 3303.1200 1456.6600 3304.7200 1457.1400 ;
        RECT 3303.1200 1462.1000 3304.7200 1462.5800 ;
        RECT 3303.1200 1467.5400 3304.7200 1468.0200 ;
        RECT 3303.1200 1472.9800 3304.7200 1473.4600 ;
        RECT 3303.1200 1478.4200 3304.7200 1478.9000 ;
        RECT 3303.1200 1483.8600 3304.7200 1484.3400 ;
        RECT 3303.1200 1489.3000 3304.7200 1489.7800 ;
        RECT 3303.1200 1494.7400 3304.7200 1495.2200 ;
        RECT 3365.4200 1445.7800 3368.4200 1446.2600 ;
        RECT 3365.4200 1451.2200 3368.4200 1451.7000 ;
        RECT 3365.4200 1456.6600 3368.4200 1457.1400 ;
        RECT 3365.4200 1462.1000 3368.4200 1462.5800 ;
        RECT 3365.4200 1467.5400 3368.4200 1468.0200 ;
        RECT 3365.4200 1472.9800 3368.4200 1473.4600 ;
        RECT 3365.4200 1478.4200 3368.4200 1478.9000 ;
        RECT 3365.4200 1483.8600 3368.4200 1484.3400 ;
        RECT 3365.4200 1489.3000 3368.4200 1489.7800 ;
        RECT 3365.4200 1494.7400 3368.4200 1495.2200 ;
        RECT 3303.1200 1500.1800 3304.7200 1500.6600 ;
        RECT 3303.1200 1505.6200 3304.7200 1506.1000 ;
        RECT 3303.1200 1511.0600 3304.7200 1511.5400 ;
        RECT 3303.1200 1516.5000 3304.7200 1516.9800 ;
        RECT 3303.1200 1521.9400 3304.7200 1522.4200 ;
        RECT 3303.1200 1527.3800 3304.7200 1527.8600 ;
        RECT 3303.1200 1532.8200 3304.7200 1533.3000 ;
        RECT 3303.1200 1538.2600 3304.7200 1538.7400 ;
        RECT 3303.1200 1543.7000 3304.7200 1544.1800 ;
        RECT 3365.4200 1500.1800 3368.4200 1500.6600 ;
        RECT 3365.4200 1505.6200 3368.4200 1506.1000 ;
        RECT 3365.4200 1511.0600 3368.4200 1511.5400 ;
        RECT 3365.4200 1516.5000 3368.4200 1516.9800 ;
        RECT 3365.4200 1521.9400 3368.4200 1522.4200 ;
        RECT 3365.4200 1527.3800 3368.4200 1527.8600 ;
        RECT 3365.4200 1532.8200 3368.4200 1533.3000 ;
        RECT 3365.4200 1538.2600 3368.4200 1538.7400 ;
        RECT 3365.4200 1543.7000 3368.4200 1544.1800 ;
        RECT 3303.1200 1549.1400 3304.7200 1549.6200 ;
        RECT 3303.1200 1554.5800 3304.7200 1555.0600 ;
        RECT 3303.1200 1560.0200 3304.7200 1560.5000 ;
        RECT 3303.1200 1565.4600 3304.7200 1565.9400 ;
        RECT 3303.1200 1570.9000 3304.7200 1571.3800 ;
        RECT 3303.1200 1587.2200 3304.7200 1587.7000 ;
        RECT 3303.1200 1576.3400 3304.7200 1576.8200 ;
        RECT 3303.1200 1581.7800 3304.7200 1582.2600 ;
        RECT 3303.1200 1592.6600 3304.7200 1593.1400 ;
        RECT 3303.1200 1598.1000 3304.7200 1598.5800 ;
        RECT 3365.4200 1549.1400 3368.4200 1549.6200 ;
        RECT 3365.4200 1554.5800 3368.4200 1555.0600 ;
        RECT 3365.4200 1560.0200 3368.4200 1560.5000 ;
        RECT 3365.4200 1565.4600 3368.4200 1565.9400 ;
        RECT 3365.4200 1570.9000 3368.4200 1571.3800 ;
        RECT 3365.4200 1587.2200 3368.4200 1587.7000 ;
        RECT 3365.4200 1576.3400 3368.4200 1576.8200 ;
        RECT 3365.4200 1581.7800 3368.4200 1582.2600 ;
        RECT 3365.4200 1592.6600 3368.4200 1593.1400 ;
        RECT 3365.4200 1598.1000 3368.4200 1598.5800 ;
        RECT 3303.1200 1603.5400 3304.7200 1604.0200 ;
        RECT 3303.1200 1608.9800 3304.7200 1609.4600 ;
        RECT 3303.1200 1614.4200 3304.7200 1614.9000 ;
        RECT 3303.1200 1619.8600 3304.7200 1620.3400 ;
        RECT 3303.1200 1625.3000 3304.7200 1625.7800 ;
        RECT 3303.1200 1630.7400 3304.7200 1631.2200 ;
        RECT 3303.1200 1636.1800 3304.7200 1636.6600 ;
        RECT 3303.1200 1641.6200 3304.7200 1642.1000 ;
        RECT 3303.1200 1647.0600 3304.7200 1647.5400 ;
        RECT 3303.1200 1652.5000 3304.7200 1652.9800 ;
        RECT 3365.4200 1603.5400 3368.4200 1604.0200 ;
        RECT 3365.4200 1608.9800 3368.4200 1609.4600 ;
        RECT 3365.4200 1614.4200 3368.4200 1614.9000 ;
        RECT 3365.4200 1619.8600 3368.4200 1620.3400 ;
        RECT 3365.4200 1625.3000 3368.4200 1625.7800 ;
        RECT 3365.4200 1630.7400 3368.4200 1631.2200 ;
        RECT 3365.4200 1636.1800 3368.4200 1636.6600 ;
        RECT 3365.4200 1641.6200 3368.4200 1642.1000 ;
        RECT 3365.4200 1647.0600 3368.4200 1647.5400 ;
        RECT 3365.4200 1652.5000 3368.4200 1652.9800 ;
        RECT 3303.1200 1679.7000 3304.7200 1680.1800 ;
        RECT 3303.1200 1657.9400 3304.7200 1658.4200 ;
        RECT 3303.1200 1663.3800 3304.7200 1663.8600 ;
        RECT 3303.1200 1668.8200 3304.7200 1669.3000 ;
        RECT 3303.1200 1674.2600 3304.7200 1674.7400 ;
        RECT 3303.1200 1685.1400 3304.7200 1685.6200 ;
        RECT 3303.1200 1690.5800 3304.7200 1691.0600 ;
        RECT 3303.1200 1696.0200 3304.7200 1696.5000 ;
        RECT 3303.1200 1701.4600 3304.7200 1701.9400 ;
        RECT 3365.4200 1679.7000 3368.4200 1680.1800 ;
        RECT 3365.4200 1657.9400 3368.4200 1658.4200 ;
        RECT 3365.4200 1663.3800 3368.4200 1663.8600 ;
        RECT 3365.4200 1668.8200 3368.4200 1669.3000 ;
        RECT 3365.4200 1674.2600 3368.4200 1674.7400 ;
        RECT 3365.4200 1685.1400 3368.4200 1685.6200 ;
        RECT 3365.4200 1690.5800 3368.4200 1691.0600 ;
        RECT 3365.4200 1696.0200 3368.4200 1696.5000 ;
        RECT 3365.4200 1701.4600 3368.4200 1701.9400 ;
        RECT 3303.1200 1706.9000 3304.7200 1707.3800 ;
        RECT 3303.1200 1712.3400 3304.7200 1712.8200 ;
        RECT 3303.1200 1717.7800 3304.7200 1718.2600 ;
        RECT 3303.1200 1723.2200 3304.7200 1723.7000 ;
        RECT 3303.1200 1728.6600 3304.7200 1729.1400 ;
        RECT 3303.1200 1734.1000 3304.7200 1734.5800 ;
        RECT 3303.1200 1739.5400 3304.7200 1740.0200 ;
        RECT 3303.1200 1744.9800 3304.7200 1745.4600 ;
        RECT 3303.1200 1750.4200 3304.7200 1750.9000 ;
        RECT 3303.1200 1755.8600 3304.7200 1756.3400 ;
        RECT 3365.4200 1706.9000 3368.4200 1707.3800 ;
        RECT 3365.4200 1712.3400 3368.4200 1712.8200 ;
        RECT 3365.4200 1717.7800 3368.4200 1718.2600 ;
        RECT 3365.4200 1723.2200 3368.4200 1723.7000 ;
        RECT 3365.4200 1728.6600 3368.4200 1729.1400 ;
        RECT 3365.4200 1734.1000 3368.4200 1734.5800 ;
        RECT 3365.4200 1739.5400 3368.4200 1740.0200 ;
        RECT 3365.4200 1744.9800 3368.4200 1745.4600 ;
        RECT 3365.4200 1750.4200 3368.4200 1750.9000 ;
        RECT 3365.4200 1755.8600 3368.4200 1756.3400 ;
        RECT 3303.1200 1761.3000 3304.7200 1761.7800 ;
        RECT 3303.1200 1766.7400 3304.7200 1767.2200 ;
        RECT 3303.1200 1772.1800 3304.7200 1772.6600 ;
        RECT 3303.1200 1777.6200 3304.7200 1778.1000 ;
        RECT 3303.1200 1783.0600 3304.7200 1783.5400 ;
        RECT 3303.1200 1788.5000 3304.7200 1788.9800 ;
        RECT 3303.1200 1793.9400 3304.7200 1794.4200 ;
        RECT 3303.1200 1799.3800 3304.7200 1799.8600 ;
        RECT 3303.1200 1804.8200 3304.7200 1805.3000 ;
        RECT 3303.1200 1810.2600 3304.7200 1810.7400 ;
        RECT 3365.4200 1761.3000 3368.4200 1761.7800 ;
        RECT 3365.4200 1766.7400 3368.4200 1767.2200 ;
        RECT 3365.4200 1772.1800 3368.4200 1772.6600 ;
        RECT 3365.4200 1777.6200 3368.4200 1778.1000 ;
        RECT 3365.4200 1783.0600 3368.4200 1783.5400 ;
        RECT 3365.4200 1788.5000 3368.4200 1788.9800 ;
        RECT 3365.4200 1793.9400 3368.4200 1794.4200 ;
        RECT 3365.4200 1799.3800 3368.4200 1799.8600 ;
        RECT 3365.4200 1804.8200 3368.4200 1805.3000 ;
        RECT 3365.4200 1810.2600 3368.4200 1810.7400 ;
        RECT 3303.1200 1837.4600 3304.7200 1837.9400 ;
        RECT 3303.1200 1815.7000 3304.7200 1816.1800 ;
        RECT 3303.1200 1821.1400 3304.7200 1821.6200 ;
        RECT 3303.1200 1826.5800 3304.7200 1827.0600 ;
        RECT 3303.1200 1832.0200 3304.7200 1832.5000 ;
        RECT 3303.1200 1842.9000 3304.7200 1843.3800 ;
        RECT 3303.1200 1848.3400 3304.7200 1848.8200 ;
        RECT 3303.1200 1853.7800 3304.7200 1854.2600 ;
        RECT 3303.1200 1859.2200 3304.7200 1859.7000 ;
        RECT 3365.4200 1837.4600 3368.4200 1837.9400 ;
        RECT 3365.4200 1815.7000 3368.4200 1816.1800 ;
        RECT 3365.4200 1821.1400 3368.4200 1821.6200 ;
        RECT 3365.4200 1826.5800 3368.4200 1827.0600 ;
        RECT 3365.4200 1832.0200 3368.4200 1832.5000 ;
        RECT 3365.4200 1842.9000 3368.4200 1843.3800 ;
        RECT 3365.4200 1848.3400 3368.4200 1848.8200 ;
        RECT 3365.4200 1853.7800 3368.4200 1854.2600 ;
        RECT 3365.4200 1859.2200 3368.4200 1859.7000 ;
        RECT 3303.1200 1864.6600 3304.7200 1865.1400 ;
        RECT 3303.1200 1870.1000 3304.7200 1870.5800 ;
        RECT 3303.1200 1875.5400 3304.7200 1876.0200 ;
        RECT 3303.1200 1880.9800 3304.7200 1881.4600 ;
        RECT 3303.1200 1886.4200 3304.7200 1886.9000 ;
        RECT 3303.1200 1891.8600 3304.7200 1892.3400 ;
        RECT 3303.1200 1897.3000 3304.7200 1897.7800 ;
        RECT 3303.1200 1902.7400 3304.7200 1903.2200 ;
        RECT 3303.1200 1908.1800 3304.7200 1908.6600 ;
        RECT 3303.1200 1913.6200 3304.7200 1914.1000 ;
        RECT 3365.4200 1864.6600 3368.4200 1865.1400 ;
        RECT 3365.4200 1870.1000 3368.4200 1870.5800 ;
        RECT 3365.4200 1875.5400 3368.4200 1876.0200 ;
        RECT 3365.4200 1880.9800 3368.4200 1881.4600 ;
        RECT 3365.4200 1886.4200 3368.4200 1886.9000 ;
        RECT 3365.4200 1891.8600 3368.4200 1892.3400 ;
        RECT 3365.4200 1897.3000 3368.4200 1897.7800 ;
        RECT 3365.4200 1902.7400 3368.4200 1903.2200 ;
        RECT 3365.4200 1908.1800 3368.4200 1908.6600 ;
        RECT 3365.4200 1913.6200 3368.4200 1914.1000 ;
        RECT 3303.1200 1929.9400 3304.7200 1930.4200 ;
        RECT 3303.1200 1919.0600 3304.7200 1919.5400 ;
        RECT 3303.1200 1924.5000 3304.7200 1924.9800 ;
        RECT 3303.1200 1935.3800 3304.7200 1935.8600 ;
        RECT 3303.1200 1940.8200 3304.7200 1941.3000 ;
        RECT 3303.1200 1946.2600 3304.7200 1946.7400 ;
        RECT 3303.1200 1951.7000 3304.7200 1952.1800 ;
        RECT 3303.1200 1957.1400 3304.7200 1957.6200 ;
        RECT 3303.1200 1962.5800 3304.7200 1963.0600 ;
        RECT 3303.1200 1968.0200 3304.7200 1968.5000 ;
        RECT 3365.4200 1929.9400 3368.4200 1930.4200 ;
        RECT 3365.4200 1919.0600 3368.4200 1919.5400 ;
        RECT 3365.4200 1924.5000 3368.4200 1924.9800 ;
        RECT 3365.4200 1935.3800 3368.4200 1935.8600 ;
        RECT 3365.4200 1940.8200 3368.4200 1941.3000 ;
        RECT 3365.4200 1946.2600 3368.4200 1946.7400 ;
        RECT 3365.4200 1951.7000 3368.4200 1952.1800 ;
        RECT 3365.4200 1957.1400 3368.4200 1957.6200 ;
        RECT 3365.4200 1962.5800 3368.4200 1963.0600 ;
        RECT 3365.4200 1968.0200 3368.4200 1968.5000 ;
        RECT 3303.1200 1973.4600 3304.7200 1973.9400 ;
        RECT 3303.1200 1978.9000 3304.7200 1979.3800 ;
        RECT 3303.1200 1984.3400 3304.7200 1984.8200 ;
        RECT 3303.1200 1989.7800 3304.7200 1990.2600 ;
        RECT 3303.1200 1995.2200 3304.7200 1995.7000 ;
        RECT 3303.1200 2000.6600 3304.7200 2001.1400 ;
        RECT 3303.1200 2006.1000 3304.7200 2006.5800 ;
        RECT 3303.1200 2011.5400 3304.7200 2012.0200 ;
        RECT 3303.1200 2016.9800 3304.7200 2017.4600 ;
        RECT 3365.4200 1973.4600 3368.4200 1973.9400 ;
        RECT 3365.4200 1978.9000 3368.4200 1979.3800 ;
        RECT 3365.4200 1984.3400 3368.4200 1984.8200 ;
        RECT 3365.4200 1989.7800 3368.4200 1990.2600 ;
        RECT 3365.4200 1995.2200 3368.4200 1995.7000 ;
        RECT 3365.4200 2000.6600 3368.4200 2001.1400 ;
        RECT 3365.4200 2006.1000 3368.4200 2006.5800 ;
        RECT 3365.4200 2011.5400 3368.4200 2012.0200 ;
        RECT 3365.4200 2016.9800 3368.4200 2017.4600 ;
        RECT 3303.1200 2022.4200 3304.7200 2022.9000 ;
        RECT 3303.1200 2027.8600 3304.7200 2028.3400 ;
        RECT 3303.1200 2033.3000 3304.7200 2033.7800 ;
        RECT 3303.1200 2038.7400 3304.7200 2039.2200 ;
        RECT 3303.1200 2044.1800 3304.7200 2044.6600 ;
        RECT 3303.1200 2049.6200 3304.7200 2050.1000 ;
        RECT 3303.1200 2055.0600 3304.7200 2055.5400 ;
        RECT 3303.1200 2060.5000 3304.7200 2060.9800 ;
        RECT 3303.1200 2065.9400 3304.7200 2066.4200 ;
        RECT 3303.1200 2071.3800 3304.7200 2071.8600 ;
        RECT 3365.4200 2022.4200 3368.4200 2022.9000 ;
        RECT 3365.4200 2027.8600 3368.4200 2028.3400 ;
        RECT 3365.4200 2033.3000 3368.4200 2033.7800 ;
        RECT 3365.4200 2038.7400 3368.4200 2039.2200 ;
        RECT 3365.4200 2044.1800 3368.4200 2044.6600 ;
        RECT 3365.4200 2049.6200 3368.4200 2050.1000 ;
        RECT 3365.4200 2055.0600 3368.4200 2055.5400 ;
        RECT 3365.4200 2060.5000 3368.4200 2060.9800 ;
        RECT 3365.4200 2065.9400 3368.4200 2066.4200 ;
        RECT 3365.4200 2071.3800 3368.4200 2071.8600 ;
        RECT 3303.1200 2087.7000 3304.7200 2088.1800 ;
        RECT 3303.1200 2076.8200 3304.7200 2077.3000 ;
        RECT 3303.1200 2082.2600 3304.7200 2082.7400 ;
        RECT 3303.1200 2093.1400 3304.7200 2093.6200 ;
        RECT 3303.1200 2098.5800 3304.7200 2099.0600 ;
        RECT 3303.1200 2104.0200 3304.7200 2104.5000 ;
        RECT 3303.1200 2109.4600 3304.7200 2109.9400 ;
        RECT 3303.1200 2114.9000 3304.7200 2115.3800 ;
        RECT 3303.1200 2120.3400 3304.7200 2120.8200 ;
        RECT 3303.1200 2125.7800 3304.7200 2126.2600 ;
        RECT 3365.4200 2087.7000 3368.4200 2088.1800 ;
        RECT 3365.4200 2076.8200 3368.4200 2077.3000 ;
        RECT 3365.4200 2082.2600 3368.4200 2082.7400 ;
        RECT 3365.4200 2093.1400 3368.4200 2093.6200 ;
        RECT 3365.4200 2098.5800 3368.4200 2099.0600 ;
        RECT 3365.4200 2104.0200 3368.4200 2104.5000 ;
        RECT 3365.4200 2109.4600 3368.4200 2109.9400 ;
        RECT 3365.4200 2114.9000 3368.4200 2115.3800 ;
        RECT 3365.4200 2120.3400 3368.4200 2120.8200 ;
        RECT 3365.4200 2125.7800 3368.4200 2126.2600 ;
        RECT 1736.3400 2259.5800 1737.9400 2260.0600 ;
        RECT 1713.7200 2486.5000 1715.3200 2486.9800 ;
        RECT 1723.7800 2522.9000 1725.3800 2523.3800 ;
        RECT 1723.7800 2528.3400 1725.3800 2528.8200 ;
        RECT 1723.7800 2533.7800 1725.3800 2534.2600 ;
        RECT 1713.7200 2522.9000 1715.3200 2523.3800 ;
        RECT 1713.7200 2528.3400 1715.3200 2528.8200 ;
        RECT 1713.7200 2533.7800 1715.3200 2534.2600 ;
        RECT 1736.2400 2522.9000 1737.8400 2523.3800 ;
        RECT 1736.2400 2528.3400 1737.8400 2528.8200 ;
        RECT 1736.2400 2533.7800 1737.8400 2534.2600 ;
        RECT 1723.7800 2539.2200 1725.3800 2539.7000 ;
        RECT 1723.7800 2544.6600 1725.3800 2545.1400 ;
        RECT 1713.7200 2539.2200 1715.3200 2539.7000 ;
        RECT 1713.7200 2544.6600 1715.3200 2545.1400 ;
        RECT 1736.2400 2539.2200 1737.8400 2539.7000 ;
        RECT 1736.2400 2544.6600 1737.8400 2545.1400 ;
        RECT 1933.9400 2486.5000 1935.5400 2486.9800 ;
        RECT 1944.0000 2461.8900 1945.6000 2464.5400 ;
        RECT 1933.9400 2522.9000 1935.5400 2523.3800 ;
        RECT 1933.9400 2528.3400 1935.5400 2528.8200 ;
        RECT 1933.9400 2533.7800 1935.5400 2534.2600 ;
        RECT 1944.0000 2522.9000 1945.6000 2523.3800 ;
        RECT 1944.0000 2528.3400 1945.6000 2528.8200 ;
        RECT 1944.0000 2533.7800 1945.6000 2534.2600 ;
        RECT 1933.9400 2539.2200 1935.5400 2539.7000 ;
        RECT 1933.9400 2544.6600 1935.5400 2545.1400 ;
        RECT 1944.0000 2539.2200 1945.6000 2539.7000 ;
        RECT 1944.0000 2544.6600 1945.6000 2545.1400 ;
        RECT 1956.4600 2522.9000 1958.0600 2523.3800 ;
        RECT 1956.4600 2528.3400 1958.0600 2528.8200 ;
        RECT 1956.4600 2533.7800 1958.0600 2534.2600 ;
        RECT 1956.4600 2539.2200 1958.0600 2539.7000 ;
        RECT 1956.4600 2544.6600 1958.0600 2545.1400 ;
        RECT 2444.5800 2337.9400 2446.1800 2338.4200 ;
        RECT 2495.5200 2337.9400 2497.1200 2338.4200 ;
        RECT 2176.7800 2259.5800 2178.3800 2260.0600 ;
        RECT 2444.5800 2232.2500 2446.1800 2234.3300 ;
        RECT 2444.5800 2131.2200 2446.1800 2131.7000 ;
        RECT 2444.5800 2136.6600 2446.1800 2137.1400 ;
        RECT 2444.5800 2142.1000 2446.1800 2142.5800 ;
        RECT 2444.5800 2147.5400 2446.1800 2148.0200 ;
        RECT 2444.5800 2152.9800 2446.1800 2153.4600 ;
        RECT 2444.5800 2158.4200 2446.1800 2158.9000 ;
        RECT 2444.5800 2163.8600 2446.1800 2164.3400 ;
        RECT 2444.5800 2169.3000 2446.1800 2169.7800 ;
        RECT 2444.5800 2174.7400 2446.1800 2175.2200 ;
        RECT 2495.5200 2131.2200 2497.1200 2131.7000 ;
        RECT 2495.5200 2136.6600 2497.1200 2137.1400 ;
        RECT 2495.5200 2142.1000 2497.1200 2142.5800 ;
        RECT 2495.5200 2147.5400 2497.1200 2148.0200 ;
        RECT 2495.5200 2152.9800 2497.1200 2153.4600 ;
        RECT 2495.5200 2158.4200 2497.1200 2158.9000 ;
        RECT 2495.5200 2163.8600 2497.1200 2164.3400 ;
        RECT 2495.5200 2169.3000 2497.1200 2169.7800 ;
        RECT 2495.5200 2174.7400 2497.1200 2175.2200 ;
        RECT 2444.5800 2180.1800 2446.1800 2180.6600 ;
        RECT 2444.5800 2185.6200 2446.1800 2186.1000 ;
        RECT 2444.5800 2191.0600 2446.1800 2191.5400 ;
        RECT 2444.5800 2196.5000 2446.1800 2196.9800 ;
        RECT 2444.5800 2201.9400 2446.1800 2202.4200 ;
        RECT 2444.5800 2207.3800 2446.1800 2207.8600 ;
        RECT 2444.5800 2212.8200 2446.1800 2213.3000 ;
        RECT 2444.5800 2218.2600 2446.1800 2218.7400 ;
        RECT 2444.5800 2223.7000 2446.1800 2224.1800 ;
        RECT 2444.5800 2229.1400 2446.1800 2229.6200 ;
        RECT 2495.5200 2180.1800 2497.1200 2180.6600 ;
        RECT 2495.5200 2185.6200 2497.1200 2186.1000 ;
        RECT 2495.5200 2191.0600 2497.1200 2191.5400 ;
        RECT 2495.5200 2196.5000 2497.1200 2196.9800 ;
        RECT 2495.5200 2201.9400 2497.1200 2202.4200 ;
        RECT 2495.5200 2207.3800 2497.1200 2207.8600 ;
        RECT 2495.5200 2212.8200 2497.1200 2213.3000 ;
        RECT 2495.5200 2218.2600 2497.1200 2218.7400 ;
        RECT 2495.5200 2223.7000 2497.1200 2224.1800 ;
        RECT 2495.5200 2229.1400 2497.1200 2229.6200 ;
        RECT 2444.5800 2240.0200 2446.1800 2240.5000 ;
        RECT 2444.5800 2250.9000 2446.1800 2251.3800 ;
        RECT 2434.4200 2259.5800 2436.0200 2260.0600 ;
        RECT 2444.5800 2261.7800 2446.1800 2262.2600 ;
        RECT 2444.5800 2267.2200 2446.1800 2267.7000 ;
        RECT 2444.5800 2272.6600 2446.1800 2273.1400 ;
        RECT 2444.5800 2278.1000 2446.1800 2278.5800 ;
        RECT 2444.5800 2283.5400 2446.1800 2284.0200 ;
        RECT 2495.5200 2234.5800 2497.1200 2235.0600 ;
        RECT 2495.5200 2240.0200 2497.1200 2240.5000 ;
        RECT 2495.5200 2245.4600 2497.1200 2245.9400 ;
        RECT 2495.5200 2250.9000 2497.1200 2251.3800 ;
        RECT 2495.5200 2256.3400 2497.1200 2256.8200 ;
        RECT 2495.5200 2261.7800 2497.1200 2262.2600 ;
        RECT 2495.5200 2267.2200 2497.1200 2267.7000 ;
        RECT 2495.5200 2272.6600 2497.1200 2273.1400 ;
        RECT 2495.5200 2278.1000 2497.1200 2278.5800 ;
        RECT 2495.5200 2283.5400 2497.1200 2284.0200 ;
        RECT 2444.5800 2288.9800 2446.1800 2289.4600 ;
        RECT 2444.5800 2294.4200 2446.1800 2294.9000 ;
        RECT 2444.5800 2299.8600 2446.1800 2300.3400 ;
        RECT 2444.5800 2305.3000 2446.1800 2305.7800 ;
        RECT 2444.5800 2310.7400 2446.1800 2311.2200 ;
        RECT 2444.5800 2316.1800 2446.1800 2316.6600 ;
        RECT 2444.5800 2321.6200 2446.1800 2322.1000 ;
        RECT 2444.5800 2327.0600 2446.1800 2327.5400 ;
        RECT 2444.5800 2332.5000 2446.1800 2332.9800 ;
        RECT 2495.5200 2288.9800 2497.1200 2289.4600 ;
        RECT 2495.5200 2294.4200 2497.1200 2294.9000 ;
        RECT 2495.5200 2299.8600 2497.1200 2300.3400 ;
        RECT 2495.5200 2305.3000 2497.1200 2305.7800 ;
        RECT 2495.5200 2310.7400 2497.1200 2311.2200 ;
        RECT 2495.5200 2316.1800 2497.1200 2316.6600 ;
        RECT 2495.5200 2321.6200 2497.1200 2322.1000 ;
        RECT 2495.5200 2327.0600 2497.1200 2327.5400 ;
        RECT 2495.5200 2332.5000 2497.1200 2332.9800 ;
        RECT 2154.1600 2486.5000 2155.7600 2486.9800 ;
        RECT 2164.2200 2461.8900 2165.8200 2464.5400 ;
        RECT 2154.1600 2522.9000 2155.7600 2523.3800 ;
        RECT 2154.1600 2528.3400 2155.7600 2528.8200 ;
        RECT 2154.1600 2533.7800 2155.7600 2534.2600 ;
        RECT 2154.1600 2539.2200 2155.7600 2539.7000 ;
        RECT 2154.1600 2544.6600 2155.7600 2545.1400 ;
        RECT 2164.2200 2522.9000 2165.8200 2523.3800 ;
        RECT 2164.2200 2528.3400 2165.8200 2528.8200 ;
        RECT 2164.2200 2533.7800 2165.8200 2534.2600 ;
        RECT 2176.6800 2522.9000 2178.2800 2523.3800 ;
        RECT 2176.6800 2528.3400 2178.2800 2528.8200 ;
        RECT 2176.6800 2533.7800 2178.2800 2534.2600 ;
        RECT 2164.2200 2539.2200 2165.8200 2539.7000 ;
        RECT 2164.2200 2544.6600 2165.8200 2545.1400 ;
        RECT 2176.6800 2539.2200 2178.2800 2539.7000 ;
        RECT 2176.6800 2544.6600 2178.2800 2545.1400 ;
        RECT 2444.5800 2343.3800 2446.1800 2343.8600 ;
        RECT 2444.5800 2348.8200 2446.1800 2349.3000 ;
        RECT 2444.5800 2354.2600 2446.1800 2354.7400 ;
        RECT 2444.5800 2359.7000 2446.1800 2360.1800 ;
        RECT 2444.5800 2365.1400 2446.1800 2365.6200 ;
        RECT 2444.5800 2370.5800 2446.1800 2371.0600 ;
        RECT 2444.5800 2376.0200 2446.1800 2376.5000 ;
        RECT 2444.5800 2381.4600 2446.1800 2381.9400 ;
        RECT 2444.5800 2386.9000 2446.1800 2387.3800 ;
        RECT 2495.5200 2343.3800 2497.1200 2343.8600 ;
        RECT 2495.5200 2348.8200 2497.1200 2349.3000 ;
        RECT 2495.5200 2354.2600 2497.1200 2354.7400 ;
        RECT 2495.5200 2359.7000 2497.1200 2360.1800 ;
        RECT 2495.5200 2365.1400 2497.1200 2365.6200 ;
        RECT 2495.5200 2370.5800 2497.1200 2371.0600 ;
        RECT 2495.5200 2376.0200 2497.1200 2376.5000 ;
        RECT 2495.5200 2381.4600 2497.1200 2381.9400 ;
        RECT 2495.5200 2386.9000 2497.1200 2387.3800 ;
        RECT 2444.5800 2392.3400 2446.1800 2392.8200 ;
        RECT 2444.5800 2397.7800 2446.1800 2398.2600 ;
        RECT 2444.5800 2403.2200 2446.1800 2403.7000 ;
        RECT 2444.5800 2408.6600 2446.1800 2409.1400 ;
        RECT 2444.5800 2414.1000 2446.1800 2414.5800 ;
        RECT 2444.5800 2419.5400 2446.1800 2420.0200 ;
        RECT 2444.5800 2424.9800 2446.1800 2425.4600 ;
        RECT 2444.5800 2430.4200 2446.1800 2430.9000 ;
        RECT 2444.5800 2435.8600 2446.1800 2436.3400 ;
        RECT 2444.5800 2441.3000 2446.1800 2441.7800 ;
        RECT 2495.5200 2392.3400 2497.1200 2392.8200 ;
        RECT 2495.5200 2397.7800 2497.1200 2398.2600 ;
        RECT 2495.5200 2403.2200 2497.1200 2403.7000 ;
        RECT 2495.5200 2408.6600 2497.1200 2409.1400 ;
        RECT 2495.5200 2414.1000 2497.1200 2414.5800 ;
        RECT 2495.5200 2419.5400 2497.1200 2420.0200 ;
        RECT 2495.5200 2424.9800 2497.1200 2425.4600 ;
        RECT 2495.5200 2430.4200 2497.1200 2430.9000 ;
        RECT 2495.5200 2435.8600 2497.1200 2436.3400 ;
        RECT 2495.5200 2441.3000 2497.1200 2441.7800 ;
        RECT 2384.4400 2495.7000 2386.0400 2496.1800 ;
        RECT 2397.0000 2495.7000 2398.6000 2496.1800 ;
        RECT 2384.4400 2479.3800 2386.0400 2479.8600 ;
        RECT 2374.3800 2486.5000 2375.9800 2486.9800 ;
        RECT 2384.4400 2483.5700 2386.0400 2485.3000 ;
        RECT 2384.4400 2490.2600 2386.0400 2490.7400 ;
        RECT 2397.0000 2479.3800 2398.6000 2479.8600 ;
        RECT 2397.0000 2484.8200 2398.6000 2485.3000 ;
        RECT 2397.0000 2490.2600 2398.6000 2490.7400 ;
        RECT 2384.4400 2501.1400 2386.0400 2501.6200 ;
        RECT 2384.4400 2507.4300 2386.0400 2507.9100 ;
        RECT 2384.4400 2512.0200 2386.0400 2512.5000 ;
        RECT 2384.4400 2517.4600 2386.0400 2517.9400 ;
        RECT 2397.0000 2501.1400 2398.6000 2501.6200 ;
        RECT 2397.0000 2506.5800 2398.6000 2507.0600 ;
        RECT 2397.0000 2512.0200 2398.6000 2512.5000 ;
        RECT 2397.0000 2517.4600 2398.6000 2517.9400 ;
        RECT 2374.3800 2522.9000 2375.9800 2523.3800 ;
        RECT 2374.3800 2528.3400 2375.9800 2528.8200 ;
        RECT 2374.3800 2533.7800 2375.9800 2534.2600 ;
        RECT 2384.4400 2522.9000 2386.0400 2523.3800 ;
        RECT 2384.4400 2528.3400 2386.0400 2528.8200 ;
        RECT 2384.4400 2533.7800 2386.0400 2534.2600 ;
        RECT 2374.3800 2539.2200 2375.9800 2539.7000 ;
        RECT 2374.3800 2544.6600 2375.9800 2545.1400 ;
        RECT 2384.4400 2539.2200 2386.0400 2539.7000 ;
        RECT 2384.4400 2544.6600 2386.0400 2545.1400 ;
        RECT 2397.0000 2533.7800 2398.6000 2534.2600 ;
        RECT 2397.0000 2528.3400 2398.6000 2528.8200 ;
        RECT 2397.0000 2522.9000 2398.6000 2523.3800 ;
        RECT 2397.0000 2544.6600 2398.6000 2545.1400 ;
        RECT 2397.0000 2539.2200 2398.6000 2539.7000 ;
        RECT 2434.4200 2495.7000 2436.0200 2496.1800 ;
        RECT 2444.5800 2495.7000 2446.1800 2496.1800 ;
        RECT 2495.5200 2495.7000 2497.1200 2496.1800 ;
        RECT 2444.5800 2446.7400 2446.1800 2447.2200 ;
        RECT 2444.5800 2452.1800 2446.1800 2452.6600 ;
        RECT 2444.5800 2457.6200 2446.1800 2458.1000 ;
        RECT 2444.5800 2461.8900 2446.1800 2463.5400 ;
        RECT 2444.5800 2468.5000 2446.1800 2468.9800 ;
        RECT 2434.4200 2479.3800 2436.0200 2479.8600 ;
        RECT 2444.5800 2473.9400 2446.1800 2474.4200 ;
        RECT 2444.5800 2479.3800 2446.1800 2479.8600 ;
        RECT 2434.4200 2484.8200 2436.0200 2485.3000 ;
        RECT 2434.4200 2490.2600 2436.0200 2490.7400 ;
        RECT 2444.5800 2484.8200 2446.1800 2485.3000 ;
        RECT 2444.5800 2490.2600 2446.1800 2490.7400 ;
        RECT 2495.5200 2446.7400 2497.1200 2447.2200 ;
        RECT 2495.5200 2452.1800 2497.1200 2452.6600 ;
        RECT 2495.5200 2457.6200 2497.1200 2458.1000 ;
        RECT 2495.5200 2463.0600 2497.1200 2463.5400 ;
        RECT 2495.5200 2468.5000 2497.1200 2468.9800 ;
        RECT 2495.5200 2473.9400 2497.1200 2474.4200 ;
        RECT 2495.5200 2479.3800 2497.1200 2479.8600 ;
        RECT 2495.5200 2484.8200 2497.1200 2485.3000 ;
        RECT 2495.5200 2490.2600 2497.1200 2490.7400 ;
        RECT 2434.4200 2501.1400 2436.0200 2501.6200 ;
        RECT 2434.4200 2506.5800 2436.0200 2507.0600 ;
        RECT 2444.5800 2501.1400 2446.1800 2501.6200 ;
        RECT 2444.5800 2506.5800 2446.1800 2507.0600 ;
        RECT 2434.4200 2512.0200 2436.0200 2512.5000 ;
        RECT 2434.4200 2517.4600 2436.0200 2517.9400 ;
        RECT 2444.5800 2512.0200 2446.1800 2512.5000 ;
        RECT 2444.5800 2517.4600 2446.1800 2517.9400 ;
        RECT 2434.4200 2522.9000 2436.0200 2523.3800 ;
        RECT 2434.4200 2528.3400 2436.0200 2528.8200 ;
        RECT 2434.4200 2533.7800 2436.0200 2534.2600 ;
        RECT 2444.5800 2522.9000 2446.1800 2523.3800 ;
        RECT 2444.5800 2528.3400 2446.1800 2528.8200 ;
        RECT 2444.5800 2533.7800 2446.1800 2534.2600 ;
        RECT 2434.4200 2539.2200 2436.0200 2539.7000 ;
        RECT 2434.4200 2544.6600 2436.0200 2545.1400 ;
        RECT 2444.5800 2539.2200 2446.1800 2539.7000 ;
        RECT 2444.5800 2544.6600 2446.1800 2545.1400 ;
        RECT 2495.5200 2501.1400 2497.1200 2501.6200 ;
        RECT 2495.5200 2506.5800 2497.1200 2507.0600 ;
        RECT 2495.5200 2512.0200 2497.1200 2512.5000 ;
        RECT 2495.5200 2517.4600 2497.1200 2517.9400 ;
        RECT 2495.5200 2522.9000 2497.1200 2523.3800 ;
        RECT 2495.5200 2528.3400 2497.1200 2528.8200 ;
        RECT 2495.5200 2533.7800 2497.1200 2534.2600 ;
        RECT 2495.5200 2539.2200 2497.1200 2539.7000 ;
        RECT 2495.5200 2544.6600 2497.1200 2545.1400 ;
        RECT 1723.7800 2550.1000 1725.3800 2550.5800 ;
        RECT 1723.7800 2555.5400 1725.3800 2556.0200 ;
        RECT 1713.7200 2550.1000 1715.3200 2550.5800 ;
        RECT 1713.7200 2555.5400 1715.3200 2556.0200 ;
        RECT 1736.2400 2550.1000 1737.8400 2550.5800 ;
        RECT 1736.2400 2555.5400 1737.8400 2556.0200 ;
        RECT 1933.9400 2550.1000 1935.5400 2550.5800 ;
        RECT 1933.9400 2555.5400 1935.5400 2556.0200 ;
        RECT 1944.0000 2550.1000 1945.6000 2550.5800 ;
        RECT 1944.0000 2555.5400 1945.6000 2556.0200 ;
        RECT 1956.4600 2550.1000 1958.0600 2550.5800 ;
        RECT 1956.4600 2555.5400 1958.0600 2556.0200 ;
        RECT 2154.1600 2550.1000 2155.7600 2550.5800 ;
        RECT 2154.1600 2555.5400 2155.7600 2556.0200 ;
        RECT 2164.2200 2550.1000 2165.8200 2550.5800 ;
        RECT 2164.2200 2555.5400 2165.8200 2556.0200 ;
        RECT 2176.6800 2550.1000 2178.2800 2550.5800 ;
        RECT 2176.6800 2555.5400 2178.2800 2556.0200 ;
        RECT 2374.3800 2550.1000 2375.9800 2550.5800 ;
        RECT 2374.3800 2555.5400 2375.9800 2556.0200 ;
        RECT 2384.4400 2550.1000 2386.0400 2550.5800 ;
        RECT 2384.4400 2555.5400 2386.0400 2556.0200 ;
        RECT 2397.0000 2550.1000 2398.6000 2550.5800 ;
        RECT 2397.0000 2555.5400 2398.6000 2556.0200 ;
        RECT 2434.4200 2550.1000 2436.0200 2550.5800 ;
        RECT 2434.4200 2555.5400 2436.0200 2556.0200 ;
        RECT 2444.5800 2550.1000 2446.1800 2550.5800 ;
        RECT 2444.5800 2555.5400 2446.1800 2556.0200 ;
        RECT 2495.5200 2550.1000 2497.1200 2550.5800 ;
        RECT 2495.5200 2555.5400 2497.1200 2556.0200 ;
        RECT 3365.4200 2337.9400 3368.4200 2338.4200 ;
        RECT 3303.1200 2337.9400 3304.7200 2338.4200 ;
        RECT 3303.1200 2131.2200 3304.7200 2131.7000 ;
        RECT 3303.1200 2136.6600 3304.7200 2137.1400 ;
        RECT 3303.1200 2142.1000 3304.7200 2142.5800 ;
        RECT 3303.1200 2147.5400 3304.7200 2148.0200 ;
        RECT 3303.1200 2152.9800 3304.7200 2153.4600 ;
        RECT 3303.1200 2158.4200 3304.7200 2158.9000 ;
        RECT 3303.1200 2163.8600 3304.7200 2164.3400 ;
        RECT 3303.1200 2169.3000 3304.7200 2169.7800 ;
        RECT 3303.1200 2174.7400 3304.7200 2175.2200 ;
        RECT 3365.4200 2131.2200 3368.4200 2131.7000 ;
        RECT 3365.4200 2136.6600 3368.4200 2137.1400 ;
        RECT 3365.4200 2142.1000 3368.4200 2142.5800 ;
        RECT 3365.4200 2147.5400 3368.4200 2148.0200 ;
        RECT 3365.4200 2152.9800 3368.4200 2153.4600 ;
        RECT 3365.4200 2158.4200 3368.4200 2158.9000 ;
        RECT 3365.4200 2163.8600 3368.4200 2164.3400 ;
        RECT 3365.4200 2169.3000 3368.4200 2169.7800 ;
        RECT 3365.4200 2174.7400 3368.4200 2175.2200 ;
        RECT 3303.1200 2180.1800 3304.7200 2180.6600 ;
        RECT 3303.1200 2185.6200 3304.7200 2186.1000 ;
        RECT 3303.1200 2191.0600 3304.7200 2191.5400 ;
        RECT 3303.1200 2196.5000 3304.7200 2196.9800 ;
        RECT 3303.1200 2201.9400 3304.7200 2202.4200 ;
        RECT 3303.1200 2207.3800 3304.7200 2207.8600 ;
        RECT 3303.1200 2212.8200 3304.7200 2213.3000 ;
        RECT 3303.1200 2218.2600 3304.7200 2218.7400 ;
        RECT 3303.1200 2223.7000 3304.7200 2224.1800 ;
        RECT 3303.1200 2229.1400 3304.7200 2229.6200 ;
        RECT 3365.4200 2180.1800 3368.4200 2180.6600 ;
        RECT 3365.4200 2185.6200 3368.4200 2186.1000 ;
        RECT 3365.4200 2191.0600 3368.4200 2191.5400 ;
        RECT 3365.4200 2196.5000 3368.4200 2196.9800 ;
        RECT 3365.4200 2201.9400 3368.4200 2202.4200 ;
        RECT 3365.4200 2207.3800 3368.4200 2207.8600 ;
        RECT 3365.4200 2212.8200 3368.4200 2213.3000 ;
        RECT 3365.4200 2218.2600 3368.4200 2218.7400 ;
        RECT 3365.4200 2223.7000 3368.4200 2224.1800 ;
        RECT 3365.4200 2229.1400 3368.4200 2229.6200 ;
        RECT 3303.1200 2234.5800 3304.7200 2235.0600 ;
        RECT 3303.1200 2240.0200 3304.7200 2240.5000 ;
        RECT 3303.1200 2245.4600 3304.7200 2245.9400 ;
        RECT 3303.1200 2250.9000 3304.7200 2251.3800 ;
        RECT 3303.1200 2256.3400 3304.7200 2256.8200 ;
        RECT 3303.1200 2261.7800 3304.7200 2262.2600 ;
        RECT 3303.1200 2267.2200 3304.7200 2267.7000 ;
        RECT 3303.1200 2272.6600 3304.7200 2273.1400 ;
        RECT 3303.1200 2278.1000 3304.7200 2278.5800 ;
        RECT 3303.1200 2283.5400 3304.7200 2284.0200 ;
        RECT 3365.4200 2234.5800 3368.4200 2235.0600 ;
        RECT 3365.4200 2240.0200 3368.4200 2240.5000 ;
        RECT 3365.4200 2245.4600 3368.4200 2245.9400 ;
        RECT 3365.4200 2250.9000 3368.4200 2251.3800 ;
        RECT 3365.4200 2256.3400 3368.4200 2256.8200 ;
        RECT 3365.4200 2261.7800 3368.4200 2262.2600 ;
        RECT 3365.4200 2267.2200 3368.4200 2267.7000 ;
        RECT 3365.4200 2272.6600 3368.4200 2273.1400 ;
        RECT 3365.4200 2278.1000 3368.4200 2278.5800 ;
        RECT 3365.4200 2283.5400 3368.4200 2284.0200 ;
        RECT 3303.1200 2288.9800 3304.7200 2289.4600 ;
        RECT 3303.1200 2294.4200 3304.7200 2294.9000 ;
        RECT 3303.1200 2299.8600 3304.7200 2300.3400 ;
        RECT 3303.1200 2305.3000 3304.7200 2305.7800 ;
        RECT 3303.1200 2310.7400 3304.7200 2311.2200 ;
        RECT 3303.1200 2316.1800 3304.7200 2316.6600 ;
        RECT 3303.1200 2321.6200 3304.7200 2322.1000 ;
        RECT 3303.1200 2327.0600 3304.7200 2327.5400 ;
        RECT 3303.1200 2332.5000 3304.7200 2332.9800 ;
        RECT 3365.4200 2288.9800 3368.4200 2289.4600 ;
        RECT 3365.4200 2294.4200 3368.4200 2294.9000 ;
        RECT 3365.4200 2299.8600 3368.4200 2300.3400 ;
        RECT 3365.4200 2305.3000 3368.4200 2305.7800 ;
        RECT 3365.4200 2310.7400 3368.4200 2311.2200 ;
        RECT 3365.4200 2316.1800 3368.4200 2316.6600 ;
        RECT 3365.4200 2321.6200 3368.4200 2322.1000 ;
        RECT 3365.4200 2327.0600 3368.4200 2327.5400 ;
        RECT 3365.4200 2332.5000 3368.4200 2332.9800 ;
        RECT 3303.1200 2343.3800 3304.7200 2343.8600 ;
        RECT 3303.1200 2348.8200 3304.7200 2349.3000 ;
        RECT 3303.1200 2354.2600 3304.7200 2354.7400 ;
        RECT 3303.1200 2359.7000 3304.7200 2360.1800 ;
        RECT 3303.1200 2365.1400 3304.7200 2365.6200 ;
        RECT 3303.1200 2370.5800 3304.7200 2371.0600 ;
        RECT 3303.1200 2376.0200 3304.7200 2376.5000 ;
        RECT 3303.1200 2381.4600 3304.7200 2381.9400 ;
        RECT 3303.1200 2386.9000 3304.7200 2387.3800 ;
        RECT 3365.4200 2343.3800 3368.4200 2343.8600 ;
        RECT 3365.4200 2348.8200 3368.4200 2349.3000 ;
        RECT 3365.4200 2354.2600 3368.4200 2354.7400 ;
        RECT 3365.4200 2359.7000 3368.4200 2360.1800 ;
        RECT 3365.4200 2365.1400 3368.4200 2365.6200 ;
        RECT 3365.4200 2370.5800 3368.4200 2371.0600 ;
        RECT 3365.4200 2376.0200 3368.4200 2376.5000 ;
        RECT 3365.4200 2381.4600 3368.4200 2381.9400 ;
        RECT 3365.4200 2386.9000 3368.4200 2387.3800 ;
        RECT 3303.1200 2392.3400 3304.7200 2392.8200 ;
        RECT 3303.1200 2397.7800 3304.7200 2398.2600 ;
        RECT 3303.1200 2403.2200 3304.7200 2403.7000 ;
        RECT 3303.1200 2408.6600 3304.7200 2409.1400 ;
        RECT 3303.1200 2414.1000 3304.7200 2414.5800 ;
        RECT 3303.1200 2419.5400 3304.7200 2420.0200 ;
        RECT 3303.1200 2424.9800 3304.7200 2425.4600 ;
        RECT 3303.1200 2430.4200 3304.7200 2430.9000 ;
        RECT 3303.1200 2435.8600 3304.7200 2436.3400 ;
        RECT 3303.1200 2441.3000 3304.7200 2441.7800 ;
        RECT 3365.4200 2392.3400 3368.4200 2392.8200 ;
        RECT 3365.4200 2397.7800 3368.4200 2398.2600 ;
        RECT 3365.4200 2403.2200 3368.4200 2403.7000 ;
        RECT 3365.4200 2408.6600 3368.4200 2409.1400 ;
        RECT 3365.4200 2414.1000 3368.4200 2414.5800 ;
        RECT 3365.4200 2419.5400 3368.4200 2420.0200 ;
        RECT 3365.4200 2424.9800 3368.4200 2425.4600 ;
        RECT 3365.4200 2430.4200 3368.4200 2430.9000 ;
        RECT 3365.4200 2435.8600 3368.4200 2436.3400 ;
        RECT 3365.4200 2441.3000 3368.4200 2441.7800 ;
        RECT 3365.4200 2495.7000 3368.4200 2496.1800 ;
        RECT 3303.1200 2495.7000 3304.7200 2496.1800 ;
        RECT 3303.1200 2446.7400 3304.7200 2447.2200 ;
        RECT 3303.1200 2452.1800 3304.7200 2452.6600 ;
        RECT 3303.1200 2457.6200 3304.7200 2458.1000 ;
        RECT 3303.1200 2463.0600 3304.7200 2463.5400 ;
        RECT 3303.1200 2468.5000 3304.7200 2468.9800 ;
        RECT 3303.1200 2473.9400 3304.7200 2474.4200 ;
        RECT 3303.1200 2479.3800 3304.7200 2479.8600 ;
        RECT 3303.1200 2484.8200 3304.7200 2485.3000 ;
        RECT 3303.1200 2490.2600 3304.7200 2490.7400 ;
        RECT 3365.4200 2446.7400 3368.4200 2447.2200 ;
        RECT 3365.4200 2452.1800 3368.4200 2452.6600 ;
        RECT 3365.4200 2457.6200 3368.4200 2458.1000 ;
        RECT 3365.4200 2463.0600 3368.4200 2463.5400 ;
        RECT 3365.4200 2468.5000 3368.4200 2468.9800 ;
        RECT 3365.4200 2473.9400 3368.4200 2474.4200 ;
        RECT 3365.4200 2479.3800 3368.4200 2479.8600 ;
        RECT 3365.4200 2484.8200 3368.4200 2485.3000 ;
        RECT 3365.4200 2490.2600 3368.4200 2490.7400 ;
        RECT 3303.1200 2501.1400 3304.7200 2501.6200 ;
        RECT 3303.1200 2506.5800 3304.7200 2507.0600 ;
        RECT 3303.1200 2512.0200 3304.7200 2512.5000 ;
        RECT 3303.1200 2517.4600 3304.7200 2517.9400 ;
        RECT 3303.1200 2522.9000 3304.7200 2523.3800 ;
        RECT 3303.1200 2528.3400 3304.7200 2528.8200 ;
        RECT 3303.1200 2533.7800 3304.7200 2534.2600 ;
        RECT 3303.1200 2539.2200 3304.7200 2539.7000 ;
        RECT 3303.1200 2544.6600 3304.7200 2545.1400 ;
        RECT 3365.4200 2501.1400 3368.4200 2501.6200 ;
        RECT 3365.4200 2506.5800 3368.4200 2507.0600 ;
        RECT 3365.4200 2512.0200 3368.4200 2512.5000 ;
        RECT 3365.4200 2517.4600 3368.4200 2517.9400 ;
        RECT 3365.4200 2522.9000 3368.4200 2523.3800 ;
        RECT 3365.4200 2528.3400 3368.4200 2528.8200 ;
        RECT 3365.4200 2533.7800 3368.4200 2534.2600 ;
        RECT 3365.4200 2539.2200 3368.4200 2539.7000 ;
        RECT 3365.4200 2544.6600 3368.4200 2545.1400 ;
        RECT 3303.1200 2550.1000 3304.7200 2550.5800 ;
        RECT 3303.1200 2555.5400 3304.7200 2556.0200 ;
        RECT 3365.4200 2550.1000 3368.4200 2550.5800 ;
        RECT 3365.4200 2555.5400 3368.4200 2556.0200 ;
      LAYER met4 ;
        RECT 155.5200 638.1400 157.1200 2017.5800 ;
        RECT 963.1200 638.1400 964.7200 2017.5800 ;
        RECT 1005.5200 178.8600 1007.1200 2567.7200 ;
        RECT 1063.2600 2.0000 1064.8600 2567.7200 ;
        RECT 1283.3400 2.0000 1284.9400 2567.7200 ;
        RECT 1283.4800 2.0000 1285.0800 2567.7200 ;
        RECT 1503.5600 2.0000 1505.1600 2567.7200 ;
        RECT 2.0000 2.0000 5.0000 2567.7200 ;
        RECT 1723.7800 2.0000 1725.3800 2567.7200 ;
        RECT 1944.0000 2.0000 1945.6000 2567.7200 ;
        RECT 2164.2200 2.0000 2165.8200 2567.7200 ;
        RECT 2384.4400 2.0000 2386.0400 2567.7200 ;
        RECT 2444.5800 2.0000 2446.1800 2567.7200 ;
        RECT 2495.5200 2.0000 2497.1200 2567.7200 ;
        RECT 3303.1200 2.0000 3304.7200 2567.7200 ;
        RECT 3365.4200 2.0000 3368.4200 2567.7200 ;
        RECT 505.5200 178.8600 507.1200 639.7400 ;
        RECT 663.1200 178.8600 664.7200 639.7400 ;
        RECT 1053.2000 178.8600 1054.8000 184.2600 ;
        RECT 1015.5800 178.8600 1017.1800 184.2600 ;
        RECT 1015.5800 178.8600 1017.1800 193.3200 ;
        RECT 1075.7200 172.6600 1077.3200 179.0000 ;
        RECT 1075.8200 178.8600 1077.4200 184.2600 ;
        RECT 1075.7200 138.6000 1077.3200 144.0000 ;
        RECT 1075.8200 187.0550 1077.4200 193.0800 ;
        RECT 1053.2000 402.3000 1054.8000 410.1000 ;
        RECT 1053.2000 408.5000 1054.8000 413.9000 ;
        RECT 1015.5800 408.5000 1017.1800 422.9600 ;
        RECT 1015.5800 402.3000 1017.1800 410.1000 ;
        RECT 1015.5800 408.5000 1017.1800 413.9000 ;
        RECT 1295.9000 178.6000 1297.5000 184.0000 ;
        RECT 1273.4200 172.6600 1275.0200 179.0000 ;
        RECT 1273.3200 178.8600 1274.9200 184.2600 ;
        RECT 1273.4200 138.6000 1275.0200 150.3400 ;
        RECT 1273.4200 138.6000 1275.0200 144.0000 ;
        RECT 1295.8000 138.3400 1297.4000 143.7400 ;
        RECT 1295.8000 172.4000 1297.4000 178.6700 ;
        RECT 1295.9000 186.7950 1297.5000 192.8200 ;
        RECT 1493.4000 178.6000 1495.0000 184.0000 ;
        RECT 1516.1200 178.6000 1517.7200 184.0000 ;
        RECT 1493.5000 138.3400 1495.1000 150.0800 ;
        RECT 1493.5000 138.3400 1495.1000 143.7400 ;
        RECT 1516.0200 138.3400 1517.6200 143.7400 ;
        RECT 1493.5000 172.4000 1495.1000 178.6700 ;
        RECT 1516.0200 172.4000 1517.6200 178.6700 ;
        RECT 1516.1200 186.7950 1517.7200 192.8200 ;
        RECT 1295.9000 408.2400 1297.5000 413.6400 ;
        RECT 1295.9000 402.0400 1297.5000 409.8400 ;
        RECT 1295.9000 416.4350 1297.5000 422.4600 ;
        RECT 1516.1200 402.0400 1517.7200 409.8400 ;
        RECT 1493.4000 402.0400 1495.0000 409.8400 ;
        RECT 1516.1200 408.2400 1517.7200 413.6400 ;
        RECT 1493.4000 408.2400 1495.0000 413.6400 ;
        RECT 1516.1200 416.4350 1517.7200 422.4600 ;
        RECT 1516.1200 861.3200 1517.7200 869.1200 ;
        RECT 1295.9000 861.3200 1297.5000 869.1200 ;
        RECT 1493.4000 861.3200 1495.0000 869.1200 ;
        RECT 1015.5800 861.5800 1017.1800 869.3800 ;
        RECT 1053.2000 861.5800 1054.8000 869.3800 ;
        RECT 1053.2000 638.1400 1054.8000 643.5400 ;
        RECT 1053.2000 631.9400 1054.8000 639.7400 ;
        RECT 1015.5800 631.9400 1017.1800 639.7400 ;
        RECT 1015.5800 638.1400 1017.1800 652.6000 ;
        RECT 1015.5800 638.1400 1017.1800 643.5400 ;
        RECT 1075.8200 638.1400 1077.4200 643.5400 ;
        RECT 1075.8200 632.4800 1077.4200 639.7400 ;
        RECT 1075.8200 646.3350 1077.4200 652.3600 ;
        RECT 1273.3200 638.1400 1274.9200 643.5400 ;
        RECT 1273.3200 632.4800 1274.9200 639.7400 ;
        RECT 1295.9000 631.6800 1297.5000 639.4800 ;
        RECT 1295.9000 646.0750 1297.5000 652.1000 ;
        RECT 1295.9000 637.8800 1297.5000 643.2800 ;
        RECT 1493.4000 631.6800 1495.0000 639.4800 ;
        RECT 1493.4000 637.8800 1495.0000 643.2800 ;
        RECT 1516.1200 631.6800 1517.7200 639.4800 ;
        RECT 1516.1200 646.0750 1517.7200 652.1000 ;
        RECT 1516.1200 637.8800 1517.7200 643.2800 ;
        RECT 1015.5800 867.7800 1017.1800 882.2400 ;
        RECT 1015.5800 867.7800 1017.1800 873.1800 ;
        RECT 1053.2000 867.7800 1054.8000 873.1800 ;
        RECT 1053.2000 1097.4200 1054.8000 1102.8200 ;
        RECT 1053.2000 1091.2200 1054.8000 1099.0200 ;
        RECT 1015.5800 1097.4200 1017.1800 1102.8200 ;
        RECT 1015.5800 1097.4200 1017.1800 1111.8800 ;
        RECT 1015.5800 1091.2200 1017.1800 1099.0200 ;
        RECT 1075.8200 1097.4200 1077.4200 1102.8200 ;
        RECT 1075.8200 1091.7600 1077.4200 1099.0200 ;
        RECT 1075.8200 1105.6150 1077.4200 1111.6400 ;
        RECT 1295.9000 867.5200 1297.5000 872.9200 ;
        RECT 1295.9000 875.7150 1297.5000 881.7400 ;
        RECT 1493.4000 867.5200 1495.0000 872.9200 ;
        RECT 1516.1200 867.5200 1517.7200 872.9200 ;
        RECT 1516.1200 875.7150 1517.7200 881.7400 ;
        RECT 1295.9000 1097.1600 1297.5000 1102.5600 ;
        RECT 1273.3200 1097.4200 1274.9200 1102.8200 ;
        RECT 1273.3200 1091.7600 1274.9200 1099.0200 ;
        RECT 1295.9000 1090.9600 1297.5000 1098.7600 ;
        RECT 1295.9000 1105.3550 1297.5000 1111.3800 ;
        RECT 1516.1200 1097.1600 1517.7200 1102.5600 ;
        RECT 1493.4000 1097.1600 1495.0000 1102.5600 ;
        RECT 1516.1200 1090.9600 1517.7200 1098.7600 ;
        RECT 1493.4000 1090.9600 1495.0000 1098.7600 ;
        RECT 1516.1200 1105.3550 1517.7200 1111.3800 ;
        RECT 1713.6200 178.6000 1715.2200 184.0000 ;
        RECT 1736.3400 178.6000 1737.9400 184.0000 ;
        RECT 1713.7200 138.3400 1715.3200 143.7400 ;
        RECT 1713.7200 138.3400 1715.3200 150.0800 ;
        RECT 1736.2400 138.3400 1737.8400 143.7400 ;
        RECT 1736.2400 172.4000 1737.8400 178.6700 ;
        RECT 1713.7200 172.4000 1715.3200 178.6700 ;
        RECT 1736.3400 186.7950 1737.9400 192.8200 ;
        RECT 1956.5600 178.6000 1958.1600 184.0000 ;
        RECT 1933.8400 178.6000 1935.4400 184.0000 ;
        RECT 1933.9400 138.3400 1935.5400 143.7400 ;
        RECT 1933.9400 138.3400 1935.5400 150.0800 ;
        RECT 1933.9400 172.4000 1935.5400 178.6700 ;
        RECT 1956.4600 172.4000 1958.0600 178.6700 ;
        RECT 1956.4600 138.3400 1958.0600 143.7400 ;
        RECT 1956.5600 186.7950 1958.1600 192.8200 ;
        RECT 1736.3400 416.4350 1737.9400 422.4600 ;
        RECT 1736.3400 402.0400 1737.9400 409.8400 ;
        RECT 1736.3400 408.2400 1737.9400 413.6400 ;
        RECT 1713.6200 408.2400 1715.2200 413.6400 ;
        RECT 1713.6200 402.0400 1715.2200 409.8400 ;
        RECT 1933.8400 408.2400 1935.4400 413.6400 ;
        RECT 1933.8400 402.0400 1935.4400 409.8400 ;
        RECT 2154.0600 178.6000 2155.6600 184.0000 ;
        RECT 2176.7800 178.6000 2178.3800 184.0000 ;
        RECT 2154.1600 138.3400 2155.7600 150.0800 ;
        RECT 2154.1600 172.4000 2155.7600 178.6700 ;
        RECT 2154.1600 138.3400 2155.7600 143.7400 ;
        RECT 2176.6800 138.3400 2178.2800 143.7400 ;
        RECT 2176.6800 172.4000 2178.2800 178.6700 ;
        RECT 2176.7800 186.7950 2178.3800 192.8200 ;
        RECT 2397.0000 178.6000 2398.6000 184.0000 ;
        RECT 2374.2800 178.6000 2375.8800 184.0000 ;
        RECT 2374.3800 138.3400 2375.9800 143.7400 ;
        RECT 2374.3800 138.3400 2375.9800 150.0800 ;
        RECT 2374.3800 172.4000 2375.9800 178.6700 ;
        RECT 2434.4200 178.6000 2436.0200 193.0600 ;
        RECT 2434.4200 178.6000 2436.0200 184.0000 ;
        RECT 2176.7800 416.4350 2178.3800 422.4600 ;
        RECT 2176.7800 402.0400 2178.3800 409.8400 ;
        RECT 2176.7800 408.2400 2178.3800 413.6400 ;
        RECT 2397.0000 408.2400 2398.6000 413.6400 ;
        RECT 2397.0000 402.0400 2398.6000 409.8400 ;
        RECT 2374.2800 402.0400 2375.8800 409.8400 ;
        RECT 2374.2800 408.2400 2375.8800 413.6400 ;
        RECT 2434.4200 408.2400 2436.0200 422.7000 ;
        RECT 2434.4200 402.0400 2436.0200 409.8400 ;
        RECT 2434.4200 408.2400 2436.0200 413.6400 ;
        RECT 1736.3400 861.3200 1737.9400 869.1200 ;
        RECT 1933.8400 861.3200 1935.4400 869.1200 ;
        RECT 1713.6200 861.3200 1715.2200 869.1200 ;
        RECT 2434.4200 861.3200 2436.0200 869.1200 ;
        RECT 2397.0000 861.3200 2398.6000 869.1200 ;
        RECT 2176.7800 861.3200 2178.3800 869.1200 ;
        RECT 2374.2800 861.3200 2375.8800 869.1200 ;
        RECT 1736.3400 631.6800 1737.9400 639.4800 ;
        RECT 1736.3400 646.0750 1737.9400 652.1000 ;
        RECT 1736.3400 637.8800 1737.9400 643.2800 ;
        RECT 1713.6200 637.8800 1715.2200 643.2800 ;
        RECT 1713.6200 631.6800 1715.2200 639.4800 ;
        RECT 1933.8400 637.8800 1935.4400 643.2800 ;
        RECT 1933.8400 631.6800 1935.4400 639.4800 ;
        RECT 1956.5600 637.8800 1958.1600 643.2800 ;
        RECT 1956.5600 646.0750 1958.1600 652.1000 ;
        RECT 1956.5600 632.2200 1958.1600 639.4800 ;
        RECT 2154.0600 637.8800 2155.6600 643.2800 ;
        RECT 2154.0600 632.2200 2155.6600 639.4800 ;
        RECT 2176.7800 631.6800 2178.3800 639.4800 ;
        RECT 2176.7800 637.8800 2178.3800 643.2800 ;
        RECT 2176.7800 646.0750 2178.3800 652.1000 ;
        RECT 2397.0000 631.6800 2398.6000 639.4800 ;
        RECT 2397.0000 637.8800 2398.6000 643.2800 ;
        RECT 2374.2800 637.8800 2375.8800 643.2800 ;
        RECT 2374.2800 631.6800 2375.8800 639.4800 ;
        RECT 2434.4200 637.8800 2436.0200 643.2800 ;
        RECT 2434.4200 637.8800 2436.0200 652.3400 ;
        RECT 2434.4200 631.6800 2436.0200 639.4800 ;
        RECT 1713.6200 867.5200 1715.2200 872.9200 ;
        RECT 1736.3400 867.5200 1737.9400 872.9200 ;
        RECT 1736.3400 875.7150 1737.9400 881.7400 ;
        RECT 1933.8400 867.5200 1935.4400 872.9200 ;
        RECT 1736.3400 1090.9600 1737.9400 1098.7600 ;
        RECT 1736.3400 1097.1600 1737.9400 1102.5600 ;
        RECT 1736.3400 1105.3550 1737.9400 1111.3800 ;
        RECT 1713.6200 1097.1600 1715.2200 1102.5600 ;
        RECT 1713.6200 1090.9600 1715.2200 1098.7600 ;
        RECT 1933.8400 1097.1600 1935.4400 1102.5600 ;
        RECT 1933.8400 1090.9600 1935.4400 1098.7600 ;
        RECT 1956.5600 1105.3550 1958.1600 1111.3800 ;
        RECT 1956.5600 1097.1600 1958.1600 1102.5600 ;
        RECT 1956.5600 1091.5000 1958.1600 1098.7600 ;
        RECT 2176.7800 867.5200 2178.3800 872.9200 ;
        RECT 2176.7800 875.7150 2178.3800 881.7400 ;
        RECT 2397.0000 867.5200 2398.6000 872.9200 ;
        RECT 2434.4200 867.5200 2436.0200 872.9200 ;
        RECT 2434.4200 867.5200 2436.0200 881.9800 ;
        RECT 2374.2800 867.5200 2375.8800 872.9200 ;
        RECT 2154.0600 1097.1600 2155.6600 1102.5600 ;
        RECT 2154.0600 1091.5000 2155.6600 1098.7600 ;
        RECT 2176.7800 1097.1600 2178.3800 1102.5600 ;
        RECT 2176.7800 1090.9600 2178.3800 1098.7600 ;
        RECT 2176.7800 1105.3550 2178.3800 1111.3800 ;
        RECT 2397.0000 1097.1600 2398.6000 1102.5600 ;
        RECT 2374.2800 1097.1600 2375.8800 1102.5600 ;
        RECT 2397.0000 1090.9600 2398.6000 1098.7600 ;
        RECT 2374.2800 1090.9600 2375.8800 1098.7600 ;
        RECT 2434.4200 1097.1600 2436.0200 1102.5600 ;
        RECT 2434.4200 1097.1600 2436.0200 1111.6200 ;
        RECT 2434.4200 1090.9600 2436.0200 1098.7600 ;
        RECT 1053.2000 1327.0600 1054.8000 1332.4600 ;
        RECT 1053.2000 1320.8600 1054.8000 1328.6600 ;
        RECT 1015.5800 1320.8600 1017.1800 1328.6600 ;
        RECT 1015.5800 1327.0600 1017.1800 1332.4600 ;
        RECT 1015.5800 1327.0600 1017.1800 1341.5200 ;
        RECT 1053.2000 1550.5000 1054.8000 1558.3000 ;
        RECT 1053.2000 1556.7000 1054.8000 1562.1000 ;
        RECT 1015.5800 1550.5000 1017.1800 1558.3000 ;
        RECT 1015.5800 1556.7000 1017.1800 1571.1600 ;
        RECT 1015.5800 1556.7000 1017.1800 1562.1000 ;
        RECT 1075.8200 1564.8950 1077.4200 1570.9200 ;
        RECT 1075.8200 1551.0400 1077.4200 1558.3000 ;
        RECT 1075.8200 1556.7000 1077.4200 1562.1000 ;
        RECT 1295.9000 1326.8000 1297.5000 1332.2000 ;
        RECT 1295.9000 1320.6000 1297.5000 1328.4000 ;
        RECT 1295.9000 1334.9950 1297.5000 1341.0200 ;
        RECT 1516.1200 1334.9950 1517.7200 1341.0200 ;
        RECT 1493.4000 1326.8000 1495.0000 1332.2000 ;
        RECT 1516.1200 1326.8000 1517.7200 1332.2000 ;
        RECT 1493.4000 1320.6000 1495.0000 1328.4000 ;
        RECT 1516.1200 1320.6000 1517.7200 1328.4000 ;
        RECT 1273.3200 1556.7000 1274.9200 1562.1000 ;
        RECT 1273.3200 1551.0400 1274.9200 1558.3000 ;
        RECT 1295.9000 1556.4400 1297.5000 1561.8400 ;
        RECT 1295.9000 1564.6350 1297.5000 1570.6600 ;
        RECT 1295.9000 1550.2400 1297.5000 1558.0400 ;
        RECT 1493.4000 1556.4400 1495.0000 1561.8400 ;
        RECT 1516.1200 1556.4400 1517.7200 1561.8400 ;
        RECT 1516.1200 1564.6350 1517.7200 1570.6600 ;
        RECT 1516.1200 1550.2400 1517.7200 1558.0400 ;
        RECT 1493.4000 1550.2400 1495.0000 1558.0400 ;
        RECT 1053.2000 1786.3400 1054.8000 1791.7400 ;
        RECT 1053.2000 1780.1400 1054.8000 1787.9400 ;
        RECT 1015.5800 1780.1400 1017.1800 1787.9400 ;
        RECT 1015.5800 1786.3400 1017.1800 1791.7400 ;
        RECT 1015.5800 1786.3400 1017.1800 1800.8000 ;
        RECT 1053.2000 2015.9800 1054.8000 2021.3800 ;
        RECT 1053.2000 2009.7800 1054.8000 2017.5800 ;
        RECT 1015.5800 2015.9800 1017.1800 2030.4400 ;
        RECT 1015.5800 2015.9800 1017.1800 2021.3800 ;
        RECT 1015.5800 2009.7800 1017.1800 2017.5800 ;
        RECT 1075.8200 2015.9800 1077.4200 2021.3800 ;
        RECT 1075.8200 2010.3200 1077.4200 2017.5800 ;
        RECT 1075.8200 2024.1750 1077.4200 2030.2000 ;
        RECT 1295.9000 1786.0800 1297.5000 1791.4800 ;
        RECT 1295.9000 1794.2750 1297.5000 1800.3000 ;
        RECT 1295.9000 1779.8800 1297.5000 1787.6800 ;
        RECT 1516.1200 1779.8800 1517.7200 1787.6800 ;
        RECT 1493.4000 1779.8800 1495.0000 1787.6800 ;
        RECT 1516.1200 1794.2750 1517.7200 1800.3000 ;
        RECT 1516.1200 1786.0800 1517.7200 1791.4800 ;
        RECT 1493.4000 1786.0800 1495.0000 1791.4800 ;
        RECT 1273.3200 2015.9800 1274.9200 2021.3800 ;
        RECT 1273.3200 2010.3200 1274.9200 2017.5800 ;
        RECT 1295.9000 2009.5200 1297.5000 2017.3200 ;
        RECT 1295.9000 2015.7200 1297.5000 2021.1200 ;
        RECT 1295.9000 2023.9150 1297.5000 2029.9400 ;
        RECT 1516.1200 2009.5200 1517.7200 2017.3200 ;
        RECT 1493.4000 2009.5200 1495.0000 2017.3200 ;
        RECT 1516.1200 2015.7200 1517.7200 2021.1200 ;
        RECT 1493.4000 2015.7200 1495.0000 2021.1200 ;
        RECT 1516.1200 2023.9150 1517.7200 2029.9400 ;
        RECT 1295.8000 2509.0600 1297.4000 2567.7200 ;
        RECT 1493.5000 2509.0600 1495.1000 2567.7200 ;
        RECT 1516.0200 2509.0600 1517.6200 2567.7200 ;
        RECT 1273.2800 2509.0600 1274.8800 2567.7200 ;
        RECT 1075.5800 2509.0600 1077.1800 2567.7200 ;
        RECT 1015.5800 2469.0600 1017.1800 2567.7200 ;
        RECT 1053.2000 2469.0600 1054.8000 2567.7200 ;
        RECT 1053.2000 2245.6200 1054.8000 2251.0200 ;
        RECT 1053.2000 2239.4200 1054.8000 2247.2200 ;
        RECT 1015.5800 2245.6200 1017.1800 2260.0800 ;
        RECT 1015.5800 2239.4200 1017.1800 2247.2200 ;
        RECT 1015.5800 2245.6200 1017.1800 2251.0200 ;
        RECT 1075.8200 2469.6000 1077.4200 2475.0300 ;
        RECT 1075.5800 2475.0000 1077.1800 2480.4000 ;
        RECT 1295.9000 2245.3600 1297.5000 2250.7600 ;
        RECT 1295.9000 2239.1600 1297.5000 2246.9600 ;
        RECT 1295.9000 2253.5550 1297.5000 2259.5800 ;
        RECT 1493.4000 2245.3600 1495.0000 2250.7600 ;
        RECT 1516.1200 2245.3600 1517.7200 2250.7600 ;
        RECT 1493.4000 2239.1600 1495.0000 2246.9600 ;
        RECT 1516.1200 2239.1600 1517.7200 2246.9600 ;
        RECT 1516.1200 2253.5550 1517.7200 2259.5800 ;
        RECT 1273.3200 2469.6000 1274.9200 2475.0300 ;
        RECT 1295.9000 2468.8000 1297.5000 2475.0300 ;
        RECT 1295.8000 2475.0000 1297.4000 2480.4000 ;
        RECT 1273.2800 2475.0000 1274.8800 2486.7400 ;
        RECT 1273.2800 2475.0000 1274.8800 2480.4000 ;
        RECT 1493.4000 2468.8000 1495.0000 2475.0300 ;
        RECT 1516.1200 2468.8000 1517.7200 2475.0300 ;
        RECT 1516.0200 2475.0000 1517.6200 2480.4000 ;
        RECT 1493.5000 2475.0000 1495.1000 2486.7400 ;
        RECT 1493.5000 2475.0000 1495.1000 2480.4000 ;
        RECT 1736.3400 1334.9950 1737.9400 1341.0200 ;
        RECT 1736.3400 1320.6000 1737.9400 1328.4000 ;
        RECT 1736.3400 1326.8000 1737.9400 1332.2000 ;
        RECT 1713.6200 1326.8000 1715.2200 1332.2000 ;
        RECT 1713.6200 1320.6000 1715.2200 1328.4000 ;
        RECT 1933.8400 1326.8000 1935.4400 1332.2000 ;
        RECT 1933.8400 1320.6000 1935.4400 1328.4000 ;
        RECT 1713.6200 1550.2400 1715.2200 1558.0400 ;
        RECT 1736.3400 1556.4400 1737.9400 1561.8400 ;
        RECT 1736.3400 1564.6350 1737.9400 1570.6600 ;
        RECT 1736.3400 1550.2400 1737.9400 1558.0400 ;
        RECT 1713.6200 1556.4400 1715.2200 1561.8400 ;
        RECT 1933.8400 1550.2400 1935.4400 1558.0400 ;
        RECT 1933.8400 1556.4400 1935.4400 1561.8400 ;
        RECT 1956.5600 1564.6350 1958.1600 1570.6600 ;
        RECT 1956.5600 1556.4400 1958.1600 1561.8400 ;
        RECT 1956.5600 1550.7800 1958.1600 1558.0400 ;
        RECT 2176.7800 1326.8000 2178.3800 1332.2000 ;
        RECT 2176.7800 1320.6000 2178.3800 1328.4000 ;
        RECT 2176.7800 1334.9950 2178.3800 1341.0200 ;
        RECT 2374.2800 1326.8000 2375.8800 1332.2000 ;
        RECT 2374.2800 1320.6000 2375.8800 1328.4000 ;
        RECT 2397.0000 1320.6000 2398.6000 1328.4000 ;
        RECT 2397.0000 1326.8000 2398.6000 1332.2000 ;
        RECT 2434.4200 1326.8000 2436.0200 1341.2600 ;
        RECT 2434.4200 1326.8000 2436.0200 1332.2000 ;
        RECT 2434.4200 1320.6000 2436.0200 1328.4000 ;
        RECT 2154.0600 1550.7800 2155.6600 1558.0400 ;
        RECT 2154.0600 1556.4400 2155.6600 1561.8400 ;
        RECT 2176.7800 1556.4400 2178.3800 1561.8400 ;
        RECT 2176.7800 1564.6350 2178.3800 1570.6600 ;
        RECT 2176.7800 1550.2400 2178.3800 1558.0400 ;
        RECT 2374.2800 1550.2400 2375.8800 1558.0400 ;
        RECT 2397.0000 1556.4400 2398.6000 1561.8400 ;
        RECT 2374.2800 1556.4400 2375.8800 1561.8400 ;
        RECT 2397.0000 1550.2400 2398.6000 1558.0400 ;
        RECT 2434.4200 1556.4400 2436.0200 1561.8400 ;
        RECT 2434.4200 1556.4400 2436.0200 1570.9000 ;
        RECT 2434.4200 1550.2400 2436.0200 1558.0400 ;
        RECT 1736.3400 1779.8800 1737.9400 1787.6800 ;
        RECT 1736.3400 1794.2750 1737.9400 1800.3000 ;
        RECT 1736.3400 1786.0800 1737.9400 1791.4800 ;
        RECT 1713.6200 1786.0800 1715.2200 1791.4800 ;
        RECT 1713.6200 1779.8800 1715.2200 1787.6800 ;
        RECT 1933.8400 1786.0800 1935.4400 1791.4800 ;
        RECT 1933.8400 1779.8800 1935.4400 1787.6800 ;
        RECT 1713.6200 2015.7200 1715.2200 2021.1200 ;
        RECT 1736.3400 2009.5200 1737.9400 2017.3200 ;
        RECT 1736.3400 2015.7200 1737.9400 2021.1200 ;
        RECT 1713.6200 2009.5200 1715.2200 2017.3200 ;
        RECT 1736.3400 2023.9150 1737.9400 2029.9400 ;
        RECT 1933.8400 2015.7200 1935.4400 2021.1200 ;
        RECT 1933.8400 2009.5200 1935.4400 2017.3200 ;
        RECT 1956.5600 2010.0600 1958.1600 2017.3200 ;
        RECT 1956.5600 2015.7200 1958.1600 2021.1200 ;
        RECT 1956.5600 2023.9150 1958.1600 2029.9400 ;
        RECT 2176.7800 1786.0800 2178.3800 1791.4800 ;
        RECT 2176.7800 1794.2750 2178.3800 1800.3000 ;
        RECT 2176.7800 1779.8800 2178.3800 1787.6800 ;
        RECT 2397.0000 1786.0800 2398.6000 1791.4800 ;
        RECT 2374.2800 1786.0800 2375.8800 1791.4800 ;
        RECT 2374.2800 1779.8800 2375.8800 1787.6800 ;
        RECT 2397.0000 1779.8800 2398.6000 1787.6800 ;
        RECT 2434.4200 1786.0800 2436.0200 1800.5400 ;
        RECT 2434.4200 1786.0800 2436.0200 1791.4800 ;
        RECT 2434.4200 1779.8800 2436.0200 1787.6800 ;
        RECT 2154.0600 2015.7200 2155.6600 2021.1200 ;
        RECT 2176.7800 2015.7200 2178.3800 2021.1200 ;
        RECT 2154.0600 2010.0600 2155.6600 2017.3200 ;
        RECT 2176.7800 2009.5200 2178.3800 2017.3200 ;
        RECT 2176.7800 2023.9150 2178.3800 2029.9400 ;
        RECT 2434.4200 2015.7200 2436.0200 2030.1800 ;
        RECT 2397.0000 2009.5200 2398.6000 2017.3200 ;
        RECT 2397.0000 2015.7200 2398.6000 2021.1200 ;
        RECT 2374.2800 2009.5200 2375.8800 2017.3200 ;
        RECT 2374.2800 2015.7200 2375.8800 2021.1200 ;
        RECT 2434.4200 2009.5200 2436.0200 2017.3200 ;
        RECT 2434.4200 2015.7200 2436.0200 2021.1200 ;
        RECT 1736.2400 2509.0600 1737.8400 2567.7200 ;
        RECT 1933.9400 2509.0600 1935.5400 2567.7200 ;
        RECT 1713.7200 2509.0600 1715.3200 2567.7200 ;
        RECT 2434.4200 2468.8000 2436.0200 2567.7200 ;
        RECT 2397.0000 2468.8000 2398.6000 2567.7200 ;
        RECT 1956.4600 2509.0600 1958.0600 2567.7200 ;
        RECT 2154.1600 2509.0600 2155.7600 2567.7200 ;
        RECT 2176.6800 2509.0600 2178.2800 2567.7200 ;
        RECT 2374.3800 2509.0600 2375.9800 2567.7200 ;
        RECT 1736.3400 2253.5550 1737.9400 2259.5800 ;
        RECT 1736.3400 2245.3600 1737.9400 2250.7600 ;
        RECT 1736.3400 2239.1600 1737.9400 2246.9600 ;
        RECT 1713.6200 2245.3600 1715.2200 2250.7600 ;
        RECT 1713.6200 2239.1600 1715.2200 2246.9600 ;
        RECT 1933.8400 2239.1600 1935.4400 2246.9600 ;
        RECT 1933.8400 2245.3600 1935.4400 2250.7600 ;
        RECT 1736.3400 2468.8000 1737.9400 2475.0300 ;
        RECT 1713.6200 2468.8000 1715.2200 2475.0300 ;
        RECT 1736.2400 2475.0000 1737.8400 2480.4000 ;
        RECT 1713.7200 2475.0000 1715.3200 2486.7400 ;
        RECT 1713.7200 2475.0000 1715.3200 2480.4000 ;
        RECT 1933.8400 2468.8000 1935.4400 2475.0300 ;
        RECT 1933.9400 2475.0000 1935.5400 2486.7400 ;
        RECT 1933.9400 2475.0000 1935.5400 2480.4000 ;
        RECT 1956.5600 2469.3400 1958.1600 2475.0300 ;
        RECT 1956.4600 2475.0000 1958.0600 2480.4000 ;
        RECT 2176.7800 2245.3600 2178.3800 2250.7600 ;
        RECT 2176.7800 2253.5550 2178.3800 2259.5800 ;
        RECT 2176.7800 2239.1600 2178.3800 2246.9600 ;
        RECT 2397.0000 2245.3600 2398.6000 2250.7600 ;
        RECT 2397.0000 2239.1600 2398.6000 2246.9600 ;
        RECT 2374.2800 2245.3600 2375.8800 2250.7600 ;
        RECT 2374.2800 2239.1600 2375.8800 2246.9600 ;
        RECT 2434.4200 2245.3600 2436.0200 2259.8200 ;
        RECT 2434.4200 2239.1600 2436.0200 2246.9600 ;
        RECT 2434.4200 2245.3600 2436.0200 2250.7600 ;
        RECT 2154.1600 2475.0000 2155.7600 2486.7400 ;
        RECT 2154.1600 2475.0000 2155.7600 2480.4000 ;
        RECT 2154.0600 2469.3400 2155.6600 2475.0300 ;
        RECT 2176.7800 2468.8000 2178.3800 2475.0300 ;
        RECT 2176.6800 2475.0000 2178.2800 2480.4000 ;
        RECT 2374.2800 2468.8000 2375.8800 2475.0300 ;
        RECT 2374.3800 2475.0000 2375.9800 2486.7400 ;
        RECT 2374.3800 2475.0000 2375.9800 2480.4000 ;
        RECT 1283.3400 20.5000 1285.0800 20.9800 ;
        RECT 1283.3400 2.0000 1285.0800 5.0000 ;
        RECT 1283.3400 9.6200 1285.0800 10.1000 ;
        RECT 1283.3400 15.0600 1285.0800 15.5400 ;
        RECT 1015.5800 193.0800 1017.1800 193.5600 ;
        RECT 1075.8200 193.0800 1077.4200 193.5600 ;
        RECT 1015.5800 422.7200 1017.1800 423.2000 ;
        RECT 1283.3400 25.9400 1285.0800 26.4200 ;
        RECT 1283.3400 31.3800 1285.0800 31.8600 ;
        RECT 1283.3400 36.8200 1285.0800 37.3000 ;
        RECT 1283.3400 42.2600 1285.0800 42.7400 ;
        RECT 1283.3400 47.7000 1285.0800 48.1800 ;
        RECT 1283.3400 53.1400 1285.0800 53.6200 ;
        RECT 1283.3400 58.5800 1285.0800 59.0600 ;
        RECT 1283.3400 64.0200 1285.0800 64.5000 ;
        RECT 1283.3400 69.4600 1285.0800 69.9400 ;
        RECT 1283.3400 74.9000 1285.0800 75.3800 ;
        RECT 1283.3400 80.3400 1285.0800 80.8200 ;
        RECT 1283.3400 85.7800 1285.0800 86.2600 ;
        RECT 1283.3400 91.2200 1285.0800 91.7000 ;
        RECT 1283.3400 96.6600 1285.0800 97.1400 ;
        RECT 1283.3400 112.9800 1285.0800 113.4600 ;
        RECT 1283.3400 102.1000 1285.0800 102.5800 ;
        RECT 1283.3400 107.5400 1285.0800 108.0200 ;
        RECT 1283.3400 118.4200 1285.0800 118.9000 ;
        RECT 1283.3400 123.8600 1285.0800 124.3400 ;
        RECT 1283.3400 178.6000 1285.0800 180.4600 ;
        RECT 1283.3400 138.3400 1285.0800 140.2000 ;
        RECT 1273.4200 150.1000 1275.0200 150.5800 ;
        RECT 1283.3400 129.3000 1285.0800 129.7800 ;
        RECT 1283.3400 146.9100 1285.0800 148.7700 ;
        RECT 1283.3400 166.4400 1285.0800 168.3000 ;
        RECT 1283.3400 188.6300 1285.0800 190.4900 ;
        RECT 1295.9000 192.8200 1297.5000 193.3000 ;
        RECT 1493.5000 149.8400 1495.1000 150.3200 ;
        RECT 1516.1200 192.8200 1517.7200 193.3000 ;
        RECT 1283.3400 408.2400 1285.0800 409.8400 ;
        RECT 1283.3400 395.1300 1285.0800 396.7300 ;
        RECT 1283.3400 418.2700 1285.0800 419.8700 ;
        RECT 1295.9000 422.4600 1297.5000 422.9400 ;
        RECT 1516.1200 422.4600 1517.7200 422.9400 ;
        RECT 1015.5800 652.3600 1017.1800 652.8400 ;
        RECT 1075.8200 652.3600 1077.4200 652.8400 ;
        RECT 1283.3400 624.7700 1285.0800 627.6800 ;
        RECT 1283.3400 637.8800 1285.0800 639.7400 ;
        RECT 1283.3400 647.9100 1285.0800 649.7700 ;
        RECT 1295.9000 652.1000 1297.5000 652.5800 ;
        RECT 1516.1200 652.1000 1517.7200 652.5800 ;
        RECT 1283.3400 854.4100 1285.0800 856.0100 ;
        RECT 1015.5800 882.0000 1017.1800 882.4800 ;
        RECT 1015.5800 1111.6400 1017.1800 1112.1200 ;
        RECT 1075.8200 1111.6400 1077.4200 1112.1200 ;
        RECT 1283.3400 877.5500 1285.0800 879.1500 ;
        RECT 1283.3400 867.5200 1285.0800 869.1200 ;
        RECT 1295.9000 881.7400 1297.5000 882.2200 ;
        RECT 1516.1200 881.7400 1517.7200 882.2200 ;
        RECT 1283.3400 1097.1600 1285.0800 1099.0200 ;
        RECT 1283.3400 1084.0500 1285.0800 1086.9600 ;
        RECT 1283.3400 1107.1900 1285.0800 1109.0500 ;
        RECT 1295.9000 1111.3800 1297.5000 1111.8600 ;
        RECT 1516.1200 1111.3800 1517.7200 1111.8600 ;
        RECT 1713.7200 149.8400 1715.3200 150.3200 ;
        RECT 1736.3400 192.8200 1737.9400 193.3000 ;
        RECT 1933.9400 149.8400 1935.5400 150.3200 ;
        RECT 1956.5600 192.8200 1958.1600 193.3000 ;
        RECT 1736.3400 422.4600 1737.9400 422.9400 ;
        RECT 2154.1600 149.8400 2155.7600 150.3200 ;
        RECT 2176.7800 192.8200 2178.3800 193.3000 ;
        RECT 2374.3800 149.8400 2375.9800 150.3200 ;
        RECT 2434.4200 192.8200 2436.0200 193.3000 ;
        RECT 2176.7800 422.4600 2178.3800 422.9400 ;
        RECT 2434.4200 422.4600 2436.0200 422.9400 ;
        RECT 1736.3400 652.1000 1737.9400 652.5800 ;
        RECT 1956.5600 652.1000 1958.1600 652.5800 ;
        RECT 2176.7800 652.1000 2178.3800 652.5800 ;
        RECT 2434.4200 652.1000 2436.0200 652.5800 ;
        RECT 1736.3400 881.7400 1737.9400 882.2200 ;
        RECT 1736.3400 1111.3800 1737.9400 1111.8600 ;
        RECT 1956.5600 1111.3800 1958.1600 1111.8600 ;
        RECT 2176.7800 881.7400 2178.3800 882.2200 ;
        RECT 2434.4200 881.7400 2436.0200 882.2200 ;
        RECT 2176.7800 1111.3800 2178.3800 1111.8600 ;
        RECT 2434.4200 1111.3800 2436.0200 1111.8600 ;
        RECT 1015.5800 1341.2800 1017.1800 1341.7600 ;
        RECT 1015.5800 1570.9200 1017.1800 1571.4000 ;
        RECT 1075.8200 1570.9200 1077.4200 1571.4000 ;
        RECT 1283.3400 1326.8000 1285.0800 1328.4000 ;
        RECT 1283.3400 1336.8300 1285.0800 1338.4300 ;
        RECT 1283.3400 1313.6900 1285.0800 1315.2900 ;
        RECT 1295.9000 1341.0200 1297.5000 1341.5000 ;
        RECT 1516.1200 1341.0200 1517.7200 1341.5000 ;
        RECT 1283.3400 1543.3300 1285.0800 1546.2400 ;
        RECT 1295.9000 1570.6600 1297.5000 1571.1400 ;
        RECT 1283.3400 1556.4400 1285.0800 1558.3000 ;
        RECT 1283.3400 1566.4700 1285.0800 1568.3300 ;
        RECT 1516.1200 1570.6600 1517.7200 1571.1400 ;
        RECT 1015.5800 1800.5600 1017.1800 1801.0400 ;
        RECT 1015.5800 2030.2000 1017.1800 2030.6800 ;
        RECT 1075.8200 2030.2000 1077.4200 2030.6800 ;
        RECT 1283.3400 1786.0800 1285.0800 1787.6800 ;
        RECT 1283.3400 1772.9700 1285.0800 1774.5700 ;
        RECT 1283.3400 1796.1100 1285.0800 1797.7100 ;
        RECT 1295.9000 1800.3000 1297.5000 1800.7800 ;
        RECT 1516.1200 1800.3000 1517.7200 1800.7800 ;
        RECT 1283.3400 2015.7200 1285.0800 2017.5800 ;
        RECT 1283.3400 2002.6100 1285.0800 2005.5200 ;
        RECT 1283.3400 2025.7500 1285.0800 2027.6100 ;
        RECT 1295.9000 2029.9400 1297.5000 2030.4200 ;
        RECT 1516.1200 2029.9400 1517.7200 2030.4200 ;
        RECT 1015.5800 2259.8400 1017.1800 2260.3200 ;
        RECT 1283.3400 2245.3600 1285.0800 2246.9600 ;
        RECT 1283.3400 2255.3900 1285.0800 2256.9900 ;
        RECT 1283.3400 2232.2500 1285.0800 2233.8500 ;
        RECT 1295.9000 2259.5800 1297.5000 2260.0600 ;
        RECT 1516.1200 2259.5800 1517.7200 2260.0600 ;
        RECT 1283.3400 2461.8900 1285.0800 2464.8000 ;
        RECT 1283.3400 2475.0000 1285.0800 2476.6000 ;
        RECT 1283.3400 2483.5700 1285.0800 2485.1700 ;
        RECT 1273.2800 2486.5000 1274.8800 2486.9800 ;
        RECT 1283.3400 2503.1000 1285.0800 2504.7000 ;
        RECT 1283.3400 2522.9000 1285.0800 2523.3800 ;
        RECT 1283.3400 2528.3400 1285.0800 2528.8200 ;
        RECT 1283.3400 2533.7800 1285.0800 2534.2600 ;
        RECT 1283.3400 2539.2200 1285.0800 2539.7000 ;
        RECT 1283.3400 2544.6600 1285.0800 2545.1400 ;
        RECT 1493.5000 2486.5000 1495.1000 2486.9800 ;
        RECT 1283.3400 2550.1000 1285.0800 2550.5800 ;
        RECT 1283.3400 2555.5400 1285.0800 2556.0200 ;
        RECT 1283.3400 2564.7200 1285.0800 2567.7200 ;
        RECT 1736.3400 1341.0200 1737.9400 1341.5000 ;
        RECT 1736.3400 1570.6600 1737.9400 1571.1400 ;
        RECT 1956.5600 1570.6600 1958.1600 1571.1400 ;
        RECT 2176.7800 1341.0200 2178.3800 1341.5000 ;
        RECT 2434.4200 1341.0200 2436.0200 1341.5000 ;
        RECT 2176.7800 1570.6600 2178.3800 1571.1400 ;
        RECT 2434.4200 1570.6600 2436.0200 1571.1400 ;
        RECT 1736.3400 1800.3000 1737.9400 1800.7800 ;
        RECT 1736.3400 2029.9400 1737.9400 2030.4200 ;
        RECT 1956.5600 2029.9400 1958.1600 2030.4200 ;
        RECT 2176.7800 1800.3000 2178.3800 1800.7800 ;
        RECT 2434.4200 1800.3000 2436.0200 1800.7800 ;
        RECT 2176.7800 2029.9400 2178.3800 2030.4200 ;
        RECT 2434.4200 2029.9400 2436.0200 2030.4200 ;
        RECT 1736.3400 2259.5800 1737.9400 2260.0600 ;
        RECT 1713.7200 2486.5000 1715.3200 2486.9800 ;
        RECT 1933.9400 2486.5000 1935.5400 2486.9800 ;
        RECT 2176.7800 2259.5800 2178.3800 2260.0600 ;
        RECT 2434.4200 2259.5800 2436.0200 2260.0600 ;
        RECT 2154.1600 2486.5000 2155.7600 2486.9800 ;
        RECT 2374.3800 2486.5000 2375.9800 2486.9800 ;
        RECT 1075.8200 186.2550 1077.4200 187.8550 ;
        RECT 1295.9000 185.9950 1297.5000 187.5950 ;
        RECT 1516.1200 185.9950 1517.7200 187.5950 ;
        RECT 1295.9000 415.6350 1297.5000 417.2350 ;
        RECT 1516.1200 415.6350 1517.7200 417.2350 ;
        RECT 647.8800 505.3800 649.4800 506.9800 ;
        RECT 1075.8200 645.5350 1077.4200 647.1350 ;
        RECT 1295.9000 645.2750 1297.5000 646.8750 ;
        RECT 1516.1200 645.2750 1517.7200 646.8750 ;
        RECT 1075.8200 1104.8150 1077.4200 1106.4150 ;
        RECT 1295.9000 874.9150 1297.5000 876.5150 ;
        RECT 1516.1200 874.9150 1517.7200 876.5150 ;
        RECT 1295.9000 1104.5550 1297.5000 1106.1550 ;
        RECT 1516.1200 1104.5550 1517.7200 1106.1550 ;
        RECT 1736.3400 185.9950 1737.9400 187.5950 ;
        RECT 1956.5600 185.9950 1958.1600 187.5950 ;
        RECT 1736.3400 415.6350 1737.9400 417.2350 ;
        RECT 2176.7800 185.9950 2178.3800 187.5950 ;
        RECT 2176.7800 415.6350 2178.3800 417.2350 ;
        RECT 1736.3400 645.2750 1737.9400 646.8750 ;
        RECT 1956.5600 645.2750 1958.1600 646.8750 ;
        RECT 2176.7800 645.2750 2178.3800 646.8750 ;
        RECT 1736.3400 874.9150 1737.9400 876.5150 ;
        RECT 1736.3400 1104.5550 1737.9400 1106.1550 ;
        RECT 1956.5600 1104.5550 1958.1600 1106.1550 ;
        RECT 2176.7800 874.9150 2178.3800 876.5150 ;
        RECT 2176.7800 1104.5550 2178.3800 1106.1550 ;
        RECT 1075.8200 1564.0950 1077.4200 1565.6950 ;
        RECT 1295.9000 1334.1950 1297.5000 1335.7950 ;
        RECT 1516.1200 1334.1950 1517.7200 1335.7950 ;
        RECT 1295.9000 1563.8350 1297.5000 1565.4350 ;
        RECT 1516.1200 1563.8350 1517.7200 1565.4350 ;
        RECT 947.8800 1930.9000 949.4800 1932.5000 ;
        RECT 1075.8200 2023.3750 1077.4200 2024.9750 ;
        RECT 1295.9000 1793.4750 1297.5000 1795.0750 ;
        RECT 1516.1200 1793.4750 1517.7200 1795.0750 ;
        RECT 1295.9000 2023.1150 1297.5000 2024.7150 ;
        RECT 1516.1200 2023.1150 1517.7200 2024.7150 ;
        RECT 1295.9000 2252.7550 1297.5000 2254.3550 ;
        RECT 1516.1200 2252.7550 1517.7200 2254.3550 ;
        RECT 1736.3400 1334.1950 1737.9400 1335.7950 ;
        RECT 1736.3400 1563.8350 1737.9400 1565.4350 ;
        RECT 1956.5600 1563.8350 1958.1600 1565.4350 ;
        RECT 2176.7800 1334.1950 2178.3800 1335.7950 ;
        RECT 2176.7800 1563.8350 2178.3800 1565.4350 ;
        RECT 1736.3400 1793.4750 1737.9400 1795.0750 ;
        RECT 1736.3400 2023.1150 1737.9400 2024.7150 ;
        RECT 1956.5600 2023.1150 1958.1600 2024.7150 ;
        RECT 2176.7800 1793.4750 2178.3800 1795.0750 ;
        RECT 2176.7800 2023.1150 2178.3800 2024.7150 ;
        RECT 3287.8800 1930.9000 3289.4800 1932.5000 ;
        RECT 1736.3400 2252.7550 1737.9400 2254.3550 ;
        RECT 2176.7800 2252.7550 2178.3800 2254.3550 ;
    END
# end of P/G power stripe data as pin


# P/G pin shape extracted from block 'core_sram'
    PORT
      LAYER met4 ;
        RECT 171.0800 1930.9000 949.4800 1932.5000 ;
    END
# end of P/G pin shape extracted from block 'core_sram'


# P/G pin shape extracted from block 'core_sram'
    PORT
      LAYER met4 ;
        RECT 2511.0800 1930.9000 3289.4800 1932.5000 ;
    END
# end of P/G pin shape extracted from block 'core_sram'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 183.4600 1054.8000 403.1000 ;
        RECT 1015.5800 183.4600 1017.1800 403.1000 ;
      LAYER met3 ;
        RECT 1053.2000 378.0400 1054.8000 378.5200 ;
        RECT 1053.2000 383.4800 1054.8000 383.9600 ;
        RECT 1053.2000 388.9200 1054.8000 389.4000 ;
        RECT 1053.2000 367.1600 1054.8000 367.6400 ;
        RECT 1053.2000 372.6000 1054.8000 373.0800 ;
        RECT 1053.2000 350.8400 1054.8000 351.3200 ;
        RECT 1053.2000 356.2800 1054.8000 356.7600 ;
        RECT 1053.2000 361.7200 1054.8000 362.2000 ;
        RECT 1053.2000 334.5200 1054.8000 335.0000 ;
        RECT 1053.2000 339.9600 1054.8000 340.4400 ;
        RECT 1053.2000 345.4000 1054.8000 345.8800 ;
        RECT 1053.2000 323.6400 1054.8000 324.1200 ;
        RECT 1053.2000 329.0800 1054.8000 329.5600 ;
        RECT 1053.2000 307.3200 1054.8000 307.8000 ;
        RECT 1053.2000 312.7600 1054.8000 313.2400 ;
        RECT 1053.2000 318.2000 1054.8000 318.6800 ;
        RECT 1053.2000 296.4400 1054.8000 296.9200 ;
        RECT 1053.2000 301.8800 1054.8000 302.3600 ;
        RECT 1015.5800 378.0400 1017.1800 378.5200 ;
        RECT 1015.5800 383.4800 1017.1800 383.9600 ;
        RECT 1015.5800 388.9200 1017.1800 389.4000 ;
        RECT 1015.5800 367.1600 1017.1800 367.6400 ;
        RECT 1015.5800 372.6000 1017.1800 373.0800 ;
        RECT 1015.5800 350.8400 1017.1800 351.3200 ;
        RECT 1015.5800 356.2800 1017.1800 356.7600 ;
        RECT 1015.5800 361.7200 1017.1800 362.2000 ;
        RECT 1015.5800 334.5200 1017.1800 335.0000 ;
        RECT 1015.5800 339.9600 1017.1800 340.4400 ;
        RECT 1015.5800 345.4000 1017.1800 345.8800 ;
        RECT 1015.5800 323.6400 1017.1800 324.1200 ;
        RECT 1015.5800 329.0800 1017.1800 329.5600 ;
        RECT 1015.5800 307.3200 1017.1800 307.8000 ;
        RECT 1015.5800 312.7600 1017.1800 313.2400 ;
        RECT 1015.5800 318.2000 1017.1800 318.6800 ;
        RECT 1015.5800 296.4400 1017.1800 296.9200 ;
        RECT 1015.5800 301.8800 1017.1800 302.3600 ;
        RECT 1053.2000 280.1200 1054.8000 280.6000 ;
        RECT 1053.2000 285.5600 1054.8000 286.0400 ;
        RECT 1053.2000 291.0000 1054.8000 291.4800 ;
        RECT 1053.2000 269.2400 1054.8000 269.7200 ;
        RECT 1053.2000 274.6800 1054.8000 275.1600 ;
        RECT 1053.2000 252.9200 1054.8000 253.4000 ;
        RECT 1053.2000 258.3600 1054.8000 258.8400 ;
        RECT 1053.2000 263.8000 1054.8000 264.2800 ;
        RECT 1053.2000 242.0400 1054.8000 242.5200 ;
        RECT 1053.2000 247.4800 1054.8000 247.9600 ;
        RECT 1053.2000 225.7200 1054.8000 226.2000 ;
        RECT 1053.2000 231.1600 1054.8000 231.6400 ;
        RECT 1053.2000 236.6000 1054.8000 237.0800 ;
        RECT 1053.2000 214.8400 1054.8000 215.3200 ;
        RECT 1053.2000 220.2800 1054.8000 220.7600 ;
        RECT 1053.2000 198.5200 1054.8000 199.0000 ;
        RECT 1053.2000 203.9600 1054.8000 204.4400 ;
        RECT 1053.2000 209.4000 1054.8000 209.8800 ;
        RECT 1053.2000 193.0800 1054.8000 193.5600 ;
        RECT 1015.5800 280.1200 1017.1800 280.6000 ;
        RECT 1015.5800 285.5600 1017.1800 286.0400 ;
        RECT 1015.5800 291.0000 1017.1800 291.4800 ;
        RECT 1015.5800 269.2400 1017.1800 269.7200 ;
        RECT 1015.5800 274.6800 1017.1800 275.1600 ;
        RECT 1015.5800 252.9200 1017.1800 253.4000 ;
        RECT 1015.5800 258.3600 1017.1800 258.8400 ;
        RECT 1015.5800 263.8000 1017.1800 264.2800 ;
        RECT 1015.5800 242.0400 1017.1800 242.5200 ;
        RECT 1015.5800 247.4800 1017.1800 247.9600 ;
        RECT 1015.5800 225.7200 1017.1800 226.2000 ;
        RECT 1015.5800 231.1600 1017.1800 231.6400 ;
        RECT 1015.5800 236.6000 1017.1800 237.0800 ;
        RECT 1015.5800 214.8400 1017.1800 215.3200 ;
        RECT 1015.5800 220.2800 1017.1800 220.7600 ;
        RECT 1015.5800 198.5200 1017.1800 199.0000 ;
        RECT 1015.5800 203.9600 1017.1800 204.4400 ;
        RECT 1015.5800 209.4000 1017.1800 209.8800 ;
        RECT 1015.5800 193.0800 1017.1800 193.5600 ;
        RECT 1010.1200 395.4900 1060.2600 397.0900 ;
        RECT 1010.1200 188.7900 1060.2600 190.3900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 183.4600 1017.1800 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 401.5000 1017.1800 403.1000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 183.4600 1054.8000 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 401.5000 1054.8000 403.1000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 188.7900 1011.7200 190.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 188.7900 1060.2600 190.3900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 395.4900 1011.7200 397.0900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 395.4900 1060.2600 397.0900 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 2250.2200 1054.8000 2469.8600 ;
        RECT 1015.5800 2250.2200 1017.1800 2469.8600 ;
      LAYER met3 ;
        RECT 1053.2000 2444.8000 1054.8000 2445.2800 ;
        RECT 1053.2000 2450.2400 1054.8000 2450.7200 ;
        RECT 1053.2000 2455.6800 1054.8000 2456.1600 ;
        RECT 1053.2000 2433.9200 1054.8000 2434.4000 ;
        RECT 1053.2000 2439.3600 1054.8000 2439.8400 ;
        RECT 1053.2000 2417.6000 1054.8000 2418.0800 ;
        RECT 1053.2000 2423.0400 1054.8000 2423.5200 ;
        RECT 1053.2000 2428.4800 1054.8000 2428.9600 ;
        RECT 1053.2000 2401.2800 1054.8000 2401.7600 ;
        RECT 1053.2000 2406.7200 1054.8000 2407.2000 ;
        RECT 1053.2000 2412.1600 1054.8000 2412.6400 ;
        RECT 1053.2000 2390.4000 1054.8000 2390.8800 ;
        RECT 1053.2000 2395.8400 1054.8000 2396.3200 ;
        RECT 1053.2000 2374.0800 1054.8000 2374.5600 ;
        RECT 1053.2000 2379.5200 1054.8000 2380.0000 ;
        RECT 1053.2000 2384.9600 1054.8000 2385.4400 ;
        RECT 1053.2000 2363.2000 1054.8000 2363.6800 ;
        RECT 1053.2000 2368.6400 1054.8000 2369.1200 ;
        RECT 1015.5800 2444.8000 1017.1800 2445.2800 ;
        RECT 1015.5800 2450.2400 1017.1800 2450.7200 ;
        RECT 1015.5800 2455.6800 1017.1800 2456.1600 ;
        RECT 1015.5800 2433.9200 1017.1800 2434.4000 ;
        RECT 1015.5800 2439.3600 1017.1800 2439.8400 ;
        RECT 1015.5800 2417.6000 1017.1800 2418.0800 ;
        RECT 1015.5800 2423.0400 1017.1800 2423.5200 ;
        RECT 1015.5800 2428.4800 1017.1800 2428.9600 ;
        RECT 1015.5800 2401.2800 1017.1800 2401.7600 ;
        RECT 1015.5800 2406.7200 1017.1800 2407.2000 ;
        RECT 1015.5800 2412.1600 1017.1800 2412.6400 ;
        RECT 1015.5800 2390.4000 1017.1800 2390.8800 ;
        RECT 1015.5800 2395.8400 1017.1800 2396.3200 ;
        RECT 1015.5800 2374.0800 1017.1800 2374.5600 ;
        RECT 1015.5800 2379.5200 1017.1800 2380.0000 ;
        RECT 1015.5800 2384.9600 1017.1800 2385.4400 ;
        RECT 1015.5800 2363.2000 1017.1800 2363.6800 ;
        RECT 1015.5800 2368.6400 1017.1800 2369.1200 ;
        RECT 1053.2000 2346.8800 1054.8000 2347.3600 ;
        RECT 1053.2000 2352.3200 1054.8000 2352.8000 ;
        RECT 1053.2000 2357.7600 1054.8000 2358.2400 ;
        RECT 1053.2000 2336.0000 1054.8000 2336.4800 ;
        RECT 1053.2000 2341.4400 1054.8000 2341.9200 ;
        RECT 1053.2000 2319.6800 1054.8000 2320.1600 ;
        RECT 1053.2000 2325.1200 1054.8000 2325.6000 ;
        RECT 1053.2000 2330.5600 1054.8000 2331.0400 ;
        RECT 1053.2000 2308.8000 1054.8000 2309.2800 ;
        RECT 1053.2000 2314.2400 1054.8000 2314.7200 ;
        RECT 1053.2000 2292.4800 1054.8000 2292.9600 ;
        RECT 1053.2000 2297.9200 1054.8000 2298.4000 ;
        RECT 1053.2000 2303.3600 1054.8000 2303.8400 ;
        RECT 1053.2000 2281.6000 1054.8000 2282.0800 ;
        RECT 1053.2000 2287.0400 1054.8000 2287.5200 ;
        RECT 1053.2000 2265.2800 1054.8000 2265.7600 ;
        RECT 1053.2000 2270.7200 1054.8000 2271.2000 ;
        RECT 1053.2000 2276.1600 1054.8000 2276.6400 ;
        RECT 1053.2000 2259.8400 1054.8000 2260.3200 ;
        RECT 1015.5800 2346.8800 1017.1800 2347.3600 ;
        RECT 1015.5800 2352.3200 1017.1800 2352.8000 ;
        RECT 1015.5800 2357.7600 1017.1800 2358.2400 ;
        RECT 1015.5800 2336.0000 1017.1800 2336.4800 ;
        RECT 1015.5800 2341.4400 1017.1800 2341.9200 ;
        RECT 1015.5800 2319.6800 1017.1800 2320.1600 ;
        RECT 1015.5800 2325.1200 1017.1800 2325.6000 ;
        RECT 1015.5800 2330.5600 1017.1800 2331.0400 ;
        RECT 1015.5800 2308.8000 1017.1800 2309.2800 ;
        RECT 1015.5800 2314.2400 1017.1800 2314.7200 ;
        RECT 1015.5800 2292.4800 1017.1800 2292.9600 ;
        RECT 1015.5800 2297.9200 1017.1800 2298.4000 ;
        RECT 1015.5800 2303.3600 1017.1800 2303.8400 ;
        RECT 1015.5800 2281.6000 1017.1800 2282.0800 ;
        RECT 1015.5800 2287.0400 1017.1800 2287.5200 ;
        RECT 1015.5800 2265.2800 1017.1800 2265.7600 ;
        RECT 1015.5800 2270.7200 1017.1800 2271.2000 ;
        RECT 1015.5800 2276.1600 1017.1800 2276.6400 ;
        RECT 1015.5800 2259.8400 1017.1800 2260.3200 ;
        RECT 1010.1200 2462.2500 1060.2600 2463.8500 ;
        RECT 1010.1200 2255.5500 1060.2600 2257.1500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 2250.2200 1017.1800 2251.8200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 2468.2600 1017.1800 2469.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 2250.2200 1054.8000 2251.8200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 2468.2600 1054.8000 2469.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2255.5500 1011.7200 2257.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2255.5500 1060.2600 2257.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2462.2500 1011.7200 2463.8500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2462.2500 1060.2600 2463.8500 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 2020.5800 1054.8000 2240.2200 ;
        RECT 1015.5800 2020.5800 1017.1800 2240.2200 ;
      LAYER met3 ;
        RECT 1053.2000 2215.1600 1054.8000 2215.6400 ;
        RECT 1053.2000 2220.6000 1054.8000 2221.0800 ;
        RECT 1053.2000 2226.0400 1054.8000 2226.5200 ;
        RECT 1053.2000 2204.2800 1054.8000 2204.7600 ;
        RECT 1053.2000 2209.7200 1054.8000 2210.2000 ;
        RECT 1053.2000 2187.9600 1054.8000 2188.4400 ;
        RECT 1053.2000 2193.4000 1054.8000 2193.8800 ;
        RECT 1053.2000 2198.8400 1054.8000 2199.3200 ;
        RECT 1053.2000 2171.6400 1054.8000 2172.1200 ;
        RECT 1053.2000 2177.0800 1054.8000 2177.5600 ;
        RECT 1053.2000 2182.5200 1054.8000 2183.0000 ;
        RECT 1053.2000 2160.7600 1054.8000 2161.2400 ;
        RECT 1053.2000 2166.2000 1054.8000 2166.6800 ;
        RECT 1053.2000 2144.4400 1054.8000 2144.9200 ;
        RECT 1053.2000 2149.8800 1054.8000 2150.3600 ;
        RECT 1053.2000 2155.3200 1054.8000 2155.8000 ;
        RECT 1053.2000 2133.5600 1054.8000 2134.0400 ;
        RECT 1053.2000 2139.0000 1054.8000 2139.4800 ;
        RECT 1015.5800 2215.1600 1017.1800 2215.6400 ;
        RECT 1015.5800 2220.6000 1017.1800 2221.0800 ;
        RECT 1015.5800 2226.0400 1017.1800 2226.5200 ;
        RECT 1015.5800 2204.2800 1017.1800 2204.7600 ;
        RECT 1015.5800 2209.7200 1017.1800 2210.2000 ;
        RECT 1015.5800 2187.9600 1017.1800 2188.4400 ;
        RECT 1015.5800 2193.4000 1017.1800 2193.8800 ;
        RECT 1015.5800 2198.8400 1017.1800 2199.3200 ;
        RECT 1015.5800 2171.6400 1017.1800 2172.1200 ;
        RECT 1015.5800 2177.0800 1017.1800 2177.5600 ;
        RECT 1015.5800 2182.5200 1017.1800 2183.0000 ;
        RECT 1015.5800 2160.7600 1017.1800 2161.2400 ;
        RECT 1015.5800 2166.2000 1017.1800 2166.6800 ;
        RECT 1015.5800 2144.4400 1017.1800 2144.9200 ;
        RECT 1015.5800 2149.8800 1017.1800 2150.3600 ;
        RECT 1015.5800 2155.3200 1017.1800 2155.8000 ;
        RECT 1015.5800 2133.5600 1017.1800 2134.0400 ;
        RECT 1015.5800 2139.0000 1017.1800 2139.4800 ;
        RECT 1053.2000 2117.2400 1054.8000 2117.7200 ;
        RECT 1053.2000 2122.6800 1054.8000 2123.1600 ;
        RECT 1053.2000 2128.1200 1054.8000 2128.6000 ;
        RECT 1053.2000 2106.3600 1054.8000 2106.8400 ;
        RECT 1053.2000 2111.8000 1054.8000 2112.2800 ;
        RECT 1053.2000 2090.0400 1054.8000 2090.5200 ;
        RECT 1053.2000 2095.4800 1054.8000 2095.9600 ;
        RECT 1053.2000 2100.9200 1054.8000 2101.4000 ;
        RECT 1053.2000 2079.1600 1054.8000 2079.6400 ;
        RECT 1053.2000 2084.6000 1054.8000 2085.0800 ;
        RECT 1053.2000 2062.8400 1054.8000 2063.3200 ;
        RECT 1053.2000 2068.2800 1054.8000 2068.7600 ;
        RECT 1053.2000 2073.7200 1054.8000 2074.2000 ;
        RECT 1053.2000 2051.9600 1054.8000 2052.4400 ;
        RECT 1053.2000 2057.4000 1054.8000 2057.8800 ;
        RECT 1053.2000 2035.6400 1054.8000 2036.1200 ;
        RECT 1053.2000 2041.0800 1054.8000 2041.5600 ;
        RECT 1053.2000 2046.5200 1054.8000 2047.0000 ;
        RECT 1053.2000 2030.2000 1054.8000 2030.6800 ;
        RECT 1015.5800 2117.2400 1017.1800 2117.7200 ;
        RECT 1015.5800 2122.6800 1017.1800 2123.1600 ;
        RECT 1015.5800 2128.1200 1017.1800 2128.6000 ;
        RECT 1015.5800 2106.3600 1017.1800 2106.8400 ;
        RECT 1015.5800 2111.8000 1017.1800 2112.2800 ;
        RECT 1015.5800 2090.0400 1017.1800 2090.5200 ;
        RECT 1015.5800 2095.4800 1017.1800 2095.9600 ;
        RECT 1015.5800 2100.9200 1017.1800 2101.4000 ;
        RECT 1015.5800 2079.1600 1017.1800 2079.6400 ;
        RECT 1015.5800 2084.6000 1017.1800 2085.0800 ;
        RECT 1015.5800 2062.8400 1017.1800 2063.3200 ;
        RECT 1015.5800 2068.2800 1017.1800 2068.7600 ;
        RECT 1015.5800 2073.7200 1017.1800 2074.2000 ;
        RECT 1015.5800 2051.9600 1017.1800 2052.4400 ;
        RECT 1015.5800 2057.4000 1017.1800 2057.8800 ;
        RECT 1015.5800 2035.6400 1017.1800 2036.1200 ;
        RECT 1015.5800 2041.0800 1017.1800 2041.5600 ;
        RECT 1015.5800 2046.5200 1017.1800 2047.0000 ;
        RECT 1015.5800 2030.2000 1017.1800 2030.6800 ;
        RECT 1010.1200 2232.6100 1060.2600 2234.2100 ;
        RECT 1010.1200 2025.9100 1060.2600 2027.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 2020.5800 1017.1800 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 2238.6200 1017.1800 2240.2200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 2020.5800 1054.8000 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 2238.6200 1054.8000 2240.2200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2025.9100 1011.7200 2027.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2025.9100 1060.2600 2027.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2232.6100 1011.7200 2234.2100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2232.6100 1060.2600 2234.2100 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 1790.9400 1054.8000 2010.5800 ;
        RECT 1015.5800 1790.9400 1017.1800 2010.5800 ;
      LAYER met3 ;
        RECT 1053.2000 1985.5200 1054.8000 1986.0000 ;
        RECT 1053.2000 1990.9600 1054.8000 1991.4400 ;
        RECT 1053.2000 1996.4000 1054.8000 1996.8800 ;
        RECT 1053.2000 1974.6400 1054.8000 1975.1200 ;
        RECT 1053.2000 1980.0800 1054.8000 1980.5600 ;
        RECT 1053.2000 1958.3200 1054.8000 1958.8000 ;
        RECT 1053.2000 1963.7600 1054.8000 1964.2400 ;
        RECT 1053.2000 1969.2000 1054.8000 1969.6800 ;
        RECT 1053.2000 1942.0000 1054.8000 1942.4800 ;
        RECT 1053.2000 1947.4400 1054.8000 1947.9200 ;
        RECT 1053.2000 1952.8800 1054.8000 1953.3600 ;
        RECT 1053.2000 1931.1200 1054.8000 1931.6000 ;
        RECT 1053.2000 1936.5600 1054.8000 1937.0400 ;
        RECT 1053.2000 1914.8000 1054.8000 1915.2800 ;
        RECT 1053.2000 1920.2400 1054.8000 1920.7200 ;
        RECT 1053.2000 1925.6800 1054.8000 1926.1600 ;
        RECT 1053.2000 1903.9200 1054.8000 1904.4000 ;
        RECT 1053.2000 1909.3600 1054.8000 1909.8400 ;
        RECT 1015.5800 1985.5200 1017.1800 1986.0000 ;
        RECT 1015.5800 1990.9600 1017.1800 1991.4400 ;
        RECT 1015.5800 1996.4000 1017.1800 1996.8800 ;
        RECT 1015.5800 1974.6400 1017.1800 1975.1200 ;
        RECT 1015.5800 1980.0800 1017.1800 1980.5600 ;
        RECT 1015.5800 1958.3200 1017.1800 1958.8000 ;
        RECT 1015.5800 1963.7600 1017.1800 1964.2400 ;
        RECT 1015.5800 1969.2000 1017.1800 1969.6800 ;
        RECT 1015.5800 1942.0000 1017.1800 1942.4800 ;
        RECT 1015.5800 1947.4400 1017.1800 1947.9200 ;
        RECT 1015.5800 1952.8800 1017.1800 1953.3600 ;
        RECT 1015.5800 1931.1200 1017.1800 1931.6000 ;
        RECT 1015.5800 1936.5600 1017.1800 1937.0400 ;
        RECT 1015.5800 1914.8000 1017.1800 1915.2800 ;
        RECT 1015.5800 1920.2400 1017.1800 1920.7200 ;
        RECT 1015.5800 1925.6800 1017.1800 1926.1600 ;
        RECT 1015.5800 1903.9200 1017.1800 1904.4000 ;
        RECT 1015.5800 1909.3600 1017.1800 1909.8400 ;
        RECT 1053.2000 1887.6000 1054.8000 1888.0800 ;
        RECT 1053.2000 1893.0400 1054.8000 1893.5200 ;
        RECT 1053.2000 1898.4800 1054.8000 1898.9600 ;
        RECT 1053.2000 1876.7200 1054.8000 1877.2000 ;
        RECT 1053.2000 1882.1600 1054.8000 1882.6400 ;
        RECT 1053.2000 1860.4000 1054.8000 1860.8800 ;
        RECT 1053.2000 1865.8400 1054.8000 1866.3200 ;
        RECT 1053.2000 1871.2800 1054.8000 1871.7600 ;
        RECT 1053.2000 1849.5200 1054.8000 1850.0000 ;
        RECT 1053.2000 1854.9600 1054.8000 1855.4400 ;
        RECT 1053.2000 1833.2000 1054.8000 1833.6800 ;
        RECT 1053.2000 1838.6400 1054.8000 1839.1200 ;
        RECT 1053.2000 1844.0800 1054.8000 1844.5600 ;
        RECT 1053.2000 1822.3200 1054.8000 1822.8000 ;
        RECT 1053.2000 1827.7600 1054.8000 1828.2400 ;
        RECT 1053.2000 1806.0000 1054.8000 1806.4800 ;
        RECT 1053.2000 1811.4400 1054.8000 1811.9200 ;
        RECT 1053.2000 1816.8800 1054.8000 1817.3600 ;
        RECT 1053.2000 1800.5600 1054.8000 1801.0400 ;
        RECT 1015.5800 1887.6000 1017.1800 1888.0800 ;
        RECT 1015.5800 1893.0400 1017.1800 1893.5200 ;
        RECT 1015.5800 1898.4800 1017.1800 1898.9600 ;
        RECT 1015.5800 1876.7200 1017.1800 1877.2000 ;
        RECT 1015.5800 1882.1600 1017.1800 1882.6400 ;
        RECT 1015.5800 1860.4000 1017.1800 1860.8800 ;
        RECT 1015.5800 1865.8400 1017.1800 1866.3200 ;
        RECT 1015.5800 1871.2800 1017.1800 1871.7600 ;
        RECT 1015.5800 1849.5200 1017.1800 1850.0000 ;
        RECT 1015.5800 1854.9600 1017.1800 1855.4400 ;
        RECT 1015.5800 1833.2000 1017.1800 1833.6800 ;
        RECT 1015.5800 1838.6400 1017.1800 1839.1200 ;
        RECT 1015.5800 1844.0800 1017.1800 1844.5600 ;
        RECT 1015.5800 1822.3200 1017.1800 1822.8000 ;
        RECT 1015.5800 1827.7600 1017.1800 1828.2400 ;
        RECT 1015.5800 1806.0000 1017.1800 1806.4800 ;
        RECT 1015.5800 1811.4400 1017.1800 1811.9200 ;
        RECT 1015.5800 1816.8800 1017.1800 1817.3600 ;
        RECT 1015.5800 1800.5600 1017.1800 1801.0400 ;
        RECT 1010.1200 2002.9700 1060.2600 2004.5700 ;
        RECT 1010.1200 1796.2700 1060.2600 1797.8700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1790.9400 1017.1800 1792.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 2008.9800 1017.1800 2010.5800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1790.9400 1054.8000 1792.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 2008.9800 1054.8000 2010.5800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1796.2700 1011.7200 1797.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1796.2700 1060.2600 1797.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 2002.9700 1011.7200 2004.5700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 2002.9700 1060.2600 2004.5700 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 1561.3000 1054.8000 1780.9400 ;
        RECT 1015.5800 1561.3000 1017.1800 1780.9400 ;
      LAYER met3 ;
        RECT 1053.2000 1755.8800 1054.8000 1756.3600 ;
        RECT 1053.2000 1761.3200 1054.8000 1761.8000 ;
        RECT 1053.2000 1766.7600 1054.8000 1767.2400 ;
        RECT 1053.2000 1745.0000 1054.8000 1745.4800 ;
        RECT 1053.2000 1750.4400 1054.8000 1750.9200 ;
        RECT 1053.2000 1728.6800 1054.8000 1729.1600 ;
        RECT 1053.2000 1734.1200 1054.8000 1734.6000 ;
        RECT 1053.2000 1739.5600 1054.8000 1740.0400 ;
        RECT 1053.2000 1712.3600 1054.8000 1712.8400 ;
        RECT 1053.2000 1717.8000 1054.8000 1718.2800 ;
        RECT 1053.2000 1723.2400 1054.8000 1723.7200 ;
        RECT 1053.2000 1701.4800 1054.8000 1701.9600 ;
        RECT 1053.2000 1706.9200 1054.8000 1707.4000 ;
        RECT 1053.2000 1685.1600 1054.8000 1685.6400 ;
        RECT 1053.2000 1690.6000 1054.8000 1691.0800 ;
        RECT 1053.2000 1696.0400 1054.8000 1696.5200 ;
        RECT 1053.2000 1674.2800 1054.8000 1674.7600 ;
        RECT 1053.2000 1679.7200 1054.8000 1680.2000 ;
        RECT 1015.5800 1755.8800 1017.1800 1756.3600 ;
        RECT 1015.5800 1761.3200 1017.1800 1761.8000 ;
        RECT 1015.5800 1766.7600 1017.1800 1767.2400 ;
        RECT 1015.5800 1745.0000 1017.1800 1745.4800 ;
        RECT 1015.5800 1750.4400 1017.1800 1750.9200 ;
        RECT 1015.5800 1728.6800 1017.1800 1729.1600 ;
        RECT 1015.5800 1734.1200 1017.1800 1734.6000 ;
        RECT 1015.5800 1739.5600 1017.1800 1740.0400 ;
        RECT 1015.5800 1712.3600 1017.1800 1712.8400 ;
        RECT 1015.5800 1717.8000 1017.1800 1718.2800 ;
        RECT 1015.5800 1723.2400 1017.1800 1723.7200 ;
        RECT 1015.5800 1701.4800 1017.1800 1701.9600 ;
        RECT 1015.5800 1706.9200 1017.1800 1707.4000 ;
        RECT 1015.5800 1685.1600 1017.1800 1685.6400 ;
        RECT 1015.5800 1690.6000 1017.1800 1691.0800 ;
        RECT 1015.5800 1696.0400 1017.1800 1696.5200 ;
        RECT 1015.5800 1674.2800 1017.1800 1674.7600 ;
        RECT 1015.5800 1679.7200 1017.1800 1680.2000 ;
        RECT 1053.2000 1657.9600 1054.8000 1658.4400 ;
        RECT 1053.2000 1663.4000 1054.8000 1663.8800 ;
        RECT 1053.2000 1668.8400 1054.8000 1669.3200 ;
        RECT 1053.2000 1647.0800 1054.8000 1647.5600 ;
        RECT 1053.2000 1652.5200 1054.8000 1653.0000 ;
        RECT 1053.2000 1630.7600 1054.8000 1631.2400 ;
        RECT 1053.2000 1636.2000 1054.8000 1636.6800 ;
        RECT 1053.2000 1641.6400 1054.8000 1642.1200 ;
        RECT 1053.2000 1619.8800 1054.8000 1620.3600 ;
        RECT 1053.2000 1625.3200 1054.8000 1625.8000 ;
        RECT 1053.2000 1603.5600 1054.8000 1604.0400 ;
        RECT 1053.2000 1609.0000 1054.8000 1609.4800 ;
        RECT 1053.2000 1614.4400 1054.8000 1614.9200 ;
        RECT 1053.2000 1592.6800 1054.8000 1593.1600 ;
        RECT 1053.2000 1598.1200 1054.8000 1598.6000 ;
        RECT 1053.2000 1576.3600 1054.8000 1576.8400 ;
        RECT 1053.2000 1581.8000 1054.8000 1582.2800 ;
        RECT 1053.2000 1587.2400 1054.8000 1587.7200 ;
        RECT 1053.2000 1570.9200 1054.8000 1571.4000 ;
        RECT 1015.5800 1657.9600 1017.1800 1658.4400 ;
        RECT 1015.5800 1663.4000 1017.1800 1663.8800 ;
        RECT 1015.5800 1668.8400 1017.1800 1669.3200 ;
        RECT 1015.5800 1647.0800 1017.1800 1647.5600 ;
        RECT 1015.5800 1652.5200 1017.1800 1653.0000 ;
        RECT 1015.5800 1630.7600 1017.1800 1631.2400 ;
        RECT 1015.5800 1636.2000 1017.1800 1636.6800 ;
        RECT 1015.5800 1641.6400 1017.1800 1642.1200 ;
        RECT 1015.5800 1619.8800 1017.1800 1620.3600 ;
        RECT 1015.5800 1625.3200 1017.1800 1625.8000 ;
        RECT 1015.5800 1603.5600 1017.1800 1604.0400 ;
        RECT 1015.5800 1609.0000 1017.1800 1609.4800 ;
        RECT 1015.5800 1614.4400 1017.1800 1614.9200 ;
        RECT 1015.5800 1592.6800 1017.1800 1593.1600 ;
        RECT 1015.5800 1598.1200 1017.1800 1598.6000 ;
        RECT 1015.5800 1576.3600 1017.1800 1576.8400 ;
        RECT 1015.5800 1581.8000 1017.1800 1582.2800 ;
        RECT 1015.5800 1587.2400 1017.1800 1587.7200 ;
        RECT 1015.5800 1570.9200 1017.1800 1571.4000 ;
        RECT 1010.1200 1773.3300 1060.2600 1774.9300 ;
        RECT 1010.1200 1566.6300 1060.2600 1568.2300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1561.3000 1017.1800 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1779.3400 1017.1800 1780.9400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1561.3000 1054.8000 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1779.3400 1054.8000 1780.9400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1566.6300 1011.7200 1568.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1566.6300 1060.2600 1568.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1773.3300 1011.7200 1774.9300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1773.3300 1060.2600 1774.9300 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 1331.6600 1054.8000 1551.3000 ;
        RECT 1015.5800 1331.6600 1017.1800 1551.3000 ;
      LAYER met3 ;
        RECT 1053.2000 1526.2400 1054.8000 1526.7200 ;
        RECT 1053.2000 1531.6800 1054.8000 1532.1600 ;
        RECT 1053.2000 1537.1200 1054.8000 1537.6000 ;
        RECT 1053.2000 1515.3600 1054.8000 1515.8400 ;
        RECT 1053.2000 1520.8000 1054.8000 1521.2800 ;
        RECT 1053.2000 1499.0400 1054.8000 1499.5200 ;
        RECT 1053.2000 1504.4800 1054.8000 1504.9600 ;
        RECT 1053.2000 1509.9200 1054.8000 1510.4000 ;
        RECT 1053.2000 1482.7200 1054.8000 1483.2000 ;
        RECT 1053.2000 1488.1600 1054.8000 1488.6400 ;
        RECT 1053.2000 1493.6000 1054.8000 1494.0800 ;
        RECT 1053.2000 1471.8400 1054.8000 1472.3200 ;
        RECT 1053.2000 1477.2800 1054.8000 1477.7600 ;
        RECT 1053.2000 1455.5200 1054.8000 1456.0000 ;
        RECT 1053.2000 1460.9600 1054.8000 1461.4400 ;
        RECT 1053.2000 1466.4000 1054.8000 1466.8800 ;
        RECT 1053.2000 1444.6400 1054.8000 1445.1200 ;
        RECT 1053.2000 1450.0800 1054.8000 1450.5600 ;
        RECT 1015.5800 1526.2400 1017.1800 1526.7200 ;
        RECT 1015.5800 1531.6800 1017.1800 1532.1600 ;
        RECT 1015.5800 1537.1200 1017.1800 1537.6000 ;
        RECT 1015.5800 1515.3600 1017.1800 1515.8400 ;
        RECT 1015.5800 1520.8000 1017.1800 1521.2800 ;
        RECT 1015.5800 1499.0400 1017.1800 1499.5200 ;
        RECT 1015.5800 1504.4800 1017.1800 1504.9600 ;
        RECT 1015.5800 1509.9200 1017.1800 1510.4000 ;
        RECT 1015.5800 1482.7200 1017.1800 1483.2000 ;
        RECT 1015.5800 1488.1600 1017.1800 1488.6400 ;
        RECT 1015.5800 1493.6000 1017.1800 1494.0800 ;
        RECT 1015.5800 1471.8400 1017.1800 1472.3200 ;
        RECT 1015.5800 1477.2800 1017.1800 1477.7600 ;
        RECT 1015.5800 1455.5200 1017.1800 1456.0000 ;
        RECT 1015.5800 1460.9600 1017.1800 1461.4400 ;
        RECT 1015.5800 1466.4000 1017.1800 1466.8800 ;
        RECT 1015.5800 1444.6400 1017.1800 1445.1200 ;
        RECT 1015.5800 1450.0800 1017.1800 1450.5600 ;
        RECT 1053.2000 1428.3200 1054.8000 1428.8000 ;
        RECT 1053.2000 1433.7600 1054.8000 1434.2400 ;
        RECT 1053.2000 1439.2000 1054.8000 1439.6800 ;
        RECT 1053.2000 1417.4400 1054.8000 1417.9200 ;
        RECT 1053.2000 1422.8800 1054.8000 1423.3600 ;
        RECT 1053.2000 1401.1200 1054.8000 1401.6000 ;
        RECT 1053.2000 1406.5600 1054.8000 1407.0400 ;
        RECT 1053.2000 1412.0000 1054.8000 1412.4800 ;
        RECT 1053.2000 1390.2400 1054.8000 1390.7200 ;
        RECT 1053.2000 1395.6800 1054.8000 1396.1600 ;
        RECT 1053.2000 1373.9200 1054.8000 1374.4000 ;
        RECT 1053.2000 1379.3600 1054.8000 1379.8400 ;
        RECT 1053.2000 1384.8000 1054.8000 1385.2800 ;
        RECT 1053.2000 1363.0400 1054.8000 1363.5200 ;
        RECT 1053.2000 1368.4800 1054.8000 1368.9600 ;
        RECT 1053.2000 1346.7200 1054.8000 1347.2000 ;
        RECT 1053.2000 1352.1600 1054.8000 1352.6400 ;
        RECT 1053.2000 1357.6000 1054.8000 1358.0800 ;
        RECT 1053.2000 1341.2800 1054.8000 1341.7600 ;
        RECT 1015.5800 1428.3200 1017.1800 1428.8000 ;
        RECT 1015.5800 1433.7600 1017.1800 1434.2400 ;
        RECT 1015.5800 1439.2000 1017.1800 1439.6800 ;
        RECT 1015.5800 1417.4400 1017.1800 1417.9200 ;
        RECT 1015.5800 1422.8800 1017.1800 1423.3600 ;
        RECT 1015.5800 1401.1200 1017.1800 1401.6000 ;
        RECT 1015.5800 1406.5600 1017.1800 1407.0400 ;
        RECT 1015.5800 1412.0000 1017.1800 1412.4800 ;
        RECT 1015.5800 1390.2400 1017.1800 1390.7200 ;
        RECT 1015.5800 1395.6800 1017.1800 1396.1600 ;
        RECT 1015.5800 1373.9200 1017.1800 1374.4000 ;
        RECT 1015.5800 1379.3600 1017.1800 1379.8400 ;
        RECT 1015.5800 1384.8000 1017.1800 1385.2800 ;
        RECT 1015.5800 1363.0400 1017.1800 1363.5200 ;
        RECT 1015.5800 1368.4800 1017.1800 1368.9600 ;
        RECT 1015.5800 1346.7200 1017.1800 1347.2000 ;
        RECT 1015.5800 1352.1600 1017.1800 1352.6400 ;
        RECT 1015.5800 1357.6000 1017.1800 1358.0800 ;
        RECT 1015.5800 1341.2800 1017.1800 1341.7600 ;
        RECT 1010.1200 1543.6900 1060.2600 1545.2900 ;
        RECT 1010.1200 1336.9900 1060.2600 1338.5900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1331.6600 1017.1800 1333.2600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1549.7000 1017.1800 1551.3000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1331.6600 1054.8000 1333.2600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1549.7000 1054.8000 1551.3000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1336.9900 1011.7200 1338.5900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1336.9900 1060.2600 1338.5900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1543.6900 1011.7200 1545.2900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1543.6900 1060.2600 1545.2900 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 1102.0200 1054.8000 1321.6600 ;
        RECT 1015.5800 1102.0200 1017.1800 1321.6600 ;
      LAYER met3 ;
        RECT 1053.2000 1296.6000 1054.8000 1297.0800 ;
        RECT 1053.2000 1302.0400 1054.8000 1302.5200 ;
        RECT 1053.2000 1307.4800 1054.8000 1307.9600 ;
        RECT 1053.2000 1285.7200 1054.8000 1286.2000 ;
        RECT 1053.2000 1291.1600 1054.8000 1291.6400 ;
        RECT 1053.2000 1269.4000 1054.8000 1269.8800 ;
        RECT 1053.2000 1274.8400 1054.8000 1275.3200 ;
        RECT 1053.2000 1280.2800 1054.8000 1280.7600 ;
        RECT 1053.2000 1253.0800 1054.8000 1253.5600 ;
        RECT 1053.2000 1258.5200 1054.8000 1259.0000 ;
        RECT 1053.2000 1263.9600 1054.8000 1264.4400 ;
        RECT 1053.2000 1242.2000 1054.8000 1242.6800 ;
        RECT 1053.2000 1247.6400 1054.8000 1248.1200 ;
        RECT 1053.2000 1225.8800 1054.8000 1226.3600 ;
        RECT 1053.2000 1231.3200 1054.8000 1231.8000 ;
        RECT 1053.2000 1236.7600 1054.8000 1237.2400 ;
        RECT 1053.2000 1215.0000 1054.8000 1215.4800 ;
        RECT 1053.2000 1220.4400 1054.8000 1220.9200 ;
        RECT 1015.5800 1296.6000 1017.1800 1297.0800 ;
        RECT 1015.5800 1302.0400 1017.1800 1302.5200 ;
        RECT 1015.5800 1307.4800 1017.1800 1307.9600 ;
        RECT 1015.5800 1285.7200 1017.1800 1286.2000 ;
        RECT 1015.5800 1291.1600 1017.1800 1291.6400 ;
        RECT 1015.5800 1269.4000 1017.1800 1269.8800 ;
        RECT 1015.5800 1274.8400 1017.1800 1275.3200 ;
        RECT 1015.5800 1280.2800 1017.1800 1280.7600 ;
        RECT 1015.5800 1253.0800 1017.1800 1253.5600 ;
        RECT 1015.5800 1258.5200 1017.1800 1259.0000 ;
        RECT 1015.5800 1263.9600 1017.1800 1264.4400 ;
        RECT 1015.5800 1242.2000 1017.1800 1242.6800 ;
        RECT 1015.5800 1247.6400 1017.1800 1248.1200 ;
        RECT 1015.5800 1225.8800 1017.1800 1226.3600 ;
        RECT 1015.5800 1231.3200 1017.1800 1231.8000 ;
        RECT 1015.5800 1236.7600 1017.1800 1237.2400 ;
        RECT 1015.5800 1215.0000 1017.1800 1215.4800 ;
        RECT 1015.5800 1220.4400 1017.1800 1220.9200 ;
        RECT 1053.2000 1198.6800 1054.8000 1199.1600 ;
        RECT 1053.2000 1204.1200 1054.8000 1204.6000 ;
        RECT 1053.2000 1209.5600 1054.8000 1210.0400 ;
        RECT 1053.2000 1187.8000 1054.8000 1188.2800 ;
        RECT 1053.2000 1193.2400 1054.8000 1193.7200 ;
        RECT 1053.2000 1171.4800 1054.8000 1171.9600 ;
        RECT 1053.2000 1176.9200 1054.8000 1177.4000 ;
        RECT 1053.2000 1182.3600 1054.8000 1182.8400 ;
        RECT 1053.2000 1160.6000 1054.8000 1161.0800 ;
        RECT 1053.2000 1166.0400 1054.8000 1166.5200 ;
        RECT 1053.2000 1144.2800 1054.8000 1144.7600 ;
        RECT 1053.2000 1149.7200 1054.8000 1150.2000 ;
        RECT 1053.2000 1155.1600 1054.8000 1155.6400 ;
        RECT 1053.2000 1133.4000 1054.8000 1133.8800 ;
        RECT 1053.2000 1138.8400 1054.8000 1139.3200 ;
        RECT 1053.2000 1117.0800 1054.8000 1117.5600 ;
        RECT 1053.2000 1122.5200 1054.8000 1123.0000 ;
        RECT 1053.2000 1127.9600 1054.8000 1128.4400 ;
        RECT 1053.2000 1111.6400 1054.8000 1112.1200 ;
        RECT 1015.5800 1198.6800 1017.1800 1199.1600 ;
        RECT 1015.5800 1204.1200 1017.1800 1204.6000 ;
        RECT 1015.5800 1209.5600 1017.1800 1210.0400 ;
        RECT 1015.5800 1187.8000 1017.1800 1188.2800 ;
        RECT 1015.5800 1193.2400 1017.1800 1193.7200 ;
        RECT 1015.5800 1171.4800 1017.1800 1171.9600 ;
        RECT 1015.5800 1176.9200 1017.1800 1177.4000 ;
        RECT 1015.5800 1182.3600 1017.1800 1182.8400 ;
        RECT 1015.5800 1160.6000 1017.1800 1161.0800 ;
        RECT 1015.5800 1166.0400 1017.1800 1166.5200 ;
        RECT 1015.5800 1144.2800 1017.1800 1144.7600 ;
        RECT 1015.5800 1149.7200 1017.1800 1150.2000 ;
        RECT 1015.5800 1155.1600 1017.1800 1155.6400 ;
        RECT 1015.5800 1133.4000 1017.1800 1133.8800 ;
        RECT 1015.5800 1138.8400 1017.1800 1139.3200 ;
        RECT 1015.5800 1117.0800 1017.1800 1117.5600 ;
        RECT 1015.5800 1122.5200 1017.1800 1123.0000 ;
        RECT 1015.5800 1127.9600 1017.1800 1128.4400 ;
        RECT 1015.5800 1111.6400 1017.1800 1112.1200 ;
        RECT 1010.1200 1314.0500 1060.2600 1315.6500 ;
        RECT 1010.1200 1107.3500 1060.2600 1108.9500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1102.0200 1017.1800 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1320.0600 1017.1800 1321.6600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1102.0200 1054.8000 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1320.0600 1054.8000 1321.6600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1107.3500 1011.7200 1108.9500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1107.3500 1060.2600 1108.9500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1314.0500 1011.7200 1315.6500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1314.0500 1060.2600 1315.6500 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 872.3800 1054.8000 1092.0200 ;
        RECT 1015.5800 872.3800 1017.1800 1092.0200 ;
      LAYER met3 ;
        RECT 1053.2000 1066.9600 1054.8000 1067.4400 ;
        RECT 1053.2000 1072.4000 1054.8000 1072.8800 ;
        RECT 1053.2000 1077.8400 1054.8000 1078.3200 ;
        RECT 1053.2000 1056.0800 1054.8000 1056.5600 ;
        RECT 1053.2000 1061.5200 1054.8000 1062.0000 ;
        RECT 1053.2000 1039.7600 1054.8000 1040.2400 ;
        RECT 1053.2000 1045.2000 1054.8000 1045.6800 ;
        RECT 1053.2000 1050.6400 1054.8000 1051.1200 ;
        RECT 1053.2000 1023.4400 1054.8000 1023.9200 ;
        RECT 1053.2000 1028.8800 1054.8000 1029.3600 ;
        RECT 1053.2000 1034.3200 1054.8000 1034.8000 ;
        RECT 1053.2000 1012.5600 1054.8000 1013.0400 ;
        RECT 1053.2000 1018.0000 1054.8000 1018.4800 ;
        RECT 1053.2000 996.2400 1054.8000 996.7200 ;
        RECT 1053.2000 1001.6800 1054.8000 1002.1600 ;
        RECT 1053.2000 1007.1200 1054.8000 1007.6000 ;
        RECT 1053.2000 985.3600 1054.8000 985.8400 ;
        RECT 1053.2000 990.8000 1054.8000 991.2800 ;
        RECT 1015.5800 1066.9600 1017.1800 1067.4400 ;
        RECT 1015.5800 1072.4000 1017.1800 1072.8800 ;
        RECT 1015.5800 1077.8400 1017.1800 1078.3200 ;
        RECT 1015.5800 1056.0800 1017.1800 1056.5600 ;
        RECT 1015.5800 1061.5200 1017.1800 1062.0000 ;
        RECT 1015.5800 1039.7600 1017.1800 1040.2400 ;
        RECT 1015.5800 1045.2000 1017.1800 1045.6800 ;
        RECT 1015.5800 1050.6400 1017.1800 1051.1200 ;
        RECT 1015.5800 1023.4400 1017.1800 1023.9200 ;
        RECT 1015.5800 1028.8800 1017.1800 1029.3600 ;
        RECT 1015.5800 1034.3200 1017.1800 1034.8000 ;
        RECT 1015.5800 1012.5600 1017.1800 1013.0400 ;
        RECT 1015.5800 1018.0000 1017.1800 1018.4800 ;
        RECT 1015.5800 996.2400 1017.1800 996.7200 ;
        RECT 1015.5800 1001.6800 1017.1800 1002.1600 ;
        RECT 1015.5800 1007.1200 1017.1800 1007.6000 ;
        RECT 1015.5800 985.3600 1017.1800 985.8400 ;
        RECT 1015.5800 990.8000 1017.1800 991.2800 ;
        RECT 1053.2000 969.0400 1054.8000 969.5200 ;
        RECT 1053.2000 974.4800 1054.8000 974.9600 ;
        RECT 1053.2000 979.9200 1054.8000 980.4000 ;
        RECT 1053.2000 958.1600 1054.8000 958.6400 ;
        RECT 1053.2000 963.6000 1054.8000 964.0800 ;
        RECT 1053.2000 941.8400 1054.8000 942.3200 ;
        RECT 1053.2000 947.2800 1054.8000 947.7600 ;
        RECT 1053.2000 952.7200 1054.8000 953.2000 ;
        RECT 1053.2000 930.9600 1054.8000 931.4400 ;
        RECT 1053.2000 936.4000 1054.8000 936.8800 ;
        RECT 1053.2000 914.6400 1054.8000 915.1200 ;
        RECT 1053.2000 920.0800 1054.8000 920.5600 ;
        RECT 1053.2000 925.5200 1054.8000 926.0000 ;
        RECT 1053.2000 903.7600 1054.8000 904.2400 ;
        RECT 1053.2000 909.2000 1054.8000 909.6800 ;
        RECT 1053.2000 887.4400 1054.8000 887.9200 ;
        RECT 1053.2000 892.8800 1054.8000 893.3600 ;
        RECT 1053.2000 898.3200 1054.8000 898.8000 ;
        RECT 1053.2000 882.0000 1054.8000 882.4800 ;
        RECT 1015.5800 969.0400 1017.1800 969.5200 ;
        RECT 1015.5800 974.4800 1017.1800 974.9600 ;
        RECT 1015.5800 979.9200 1017.1800 980.4000 ;
        RECT 1015.5800 958.1600 1017.1800 958.6400 ;
        RECT 1015.5800 963.6000 1017.1800 964.0800 ;
        RECT 1015.5800 941.8400 1017.1800 942.3200 ;
        RECT 1015.5800 947.2800 1017.1800 947.7600 ;
        RECT 1015.5800 952.7200 1017.1800 953.2000 ;
        RECT 1015.5800 930.9600 1017.1800 931.4400 ;
        RECT 1015.5800 936.4000 1017.1800 936.8800 ;
        RECT 1015.5800 914.6400 1017.1800 915.1200 ;
        RECT 1015.5800 920.0800 1017.1800 920.5600 ;
        RECT 1015.5800 925.5200 1017.1800 926.0000 ;
        RECT 1015.5800 903.7600 1017.1800 904.2400 ;
        RECT 1015.5800 909.2000 1017.1800 909.6800 ;
        RECT 1015.5800 887.4400 1017.1800 887.9200 ;
        RECT 1015.5800 892.8800 1017.1800 893.3600 ;
        RECT 1015.5800 898.3200 1017.1800 898.8000 ;
        RECT 1015.5800 882.0000 1017.1800 882.4800 ;
        RECT 1010.1200 1084.4100 1060.2600 1086.0100 ;
        RECT 1010.1200 877.7100 1060.2600 879.3100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 872.3800 1017.1800 873.9800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 1090.4200 1017.1800 1092.0200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 872.3800 1054.8000 873.9800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 1090.4200 1054.8000 1092.0200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 877.7100 1011.7200 879.3100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 877.7100 1060.2600 879.3100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 1084.4100 1011.7200 1086.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 1084.4100 1060.2600 1086.0100 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 642.7400 1054.8000 862.3800 ;
        RECT 1015.5800 642.7400 1017.1800 862.3800 ;
      LAYER met3 ;
        RECT 1053.2000 837.3200 1054.8000 837.8000 ;
        RECT 1053.2000 842.7600 1054.8000 843.2400 ;
        RECT 1053.2000 848.2000 1054.8000 848.6800 ;
        RECT 1053.2000 826.4400 1054.8000 826.9200 ;
        RECT 1053.2000 831.8800 1054.8000 832.3600 ;
        RECT 1053.2000 810.1200 1054.8000 810.6000 ;
        RECT 1053.2000 815.5600 1054.8000 816.0400 ;
        RECT 1053.2000 821.0000 1054.8000 821.4800 ;
        RECT 1053.2000 793.8000 1054.8000 794.2800 ;
        RECT 1053.2000 799.2400 1054.8000 799.7200 ;
        RECT 1053.2000 804.6800 1054.8000 805.1600 ;
        RECT 1053.2000 782.9200 1054.8000 783.4000 ;
        RECT 1053.2000 788.3600 1054.8000 788.8400 ;
        RECT 1053.2000 766.6000 1054.8000 767.0800 ;
        RECT 1053.2000 772.0400 1054.8000 772.5200 ;
        RECT 1053.2000 777.4800 1054.8000 777.9600 ;
        RECT 1053.2000 755.7200 1054.8000 756.2000 ;
        RECT 1053.2000 761.1600 1054.8000 761.6400 ;
        RECT 1015.5800 837.3200 1017.1800 837.8000 ;
        RECT 1015.5800 842.7600 1017.1800 843.2400 ;
        RECT 1015.5800 848.2000 1017.1800 848.6800 ;
        RECT 1015.5800 826.4400 1017.1800 826.9200 ;
        RECT 1015.5800 831.8800 1017.1800 832.3600 ;
        RECT 1015.5800 810.1200 1017.1800 810.6000 ;
        RECT 1015.5800 815.5600 1017.1800 816.0400 ;
        RECT 1015.5800 821.0000 1017.1800 821.4800 ;
        RECT 1015.5800 793.8000 1017.1800 794.2800 ;
        RECT 1015.5800 799.2400 1017.1800 799.7200 ;
        RECT 1015.5800 804.6800 1017.1800 805.1600 ;
        RECT 1015.5800 782.9200 1017.1800 783.4000 ;
        RECT 1015.5800 788.3600 1017.1800 788.8400 ;
        RECT 1015.5800 766.6000 1017.1800 767.0800 ;
        RECT 1015.5800 772.0400 1017.1800 772.5200 ;
        RECT 1015.5800 777.4800 1017.1800 777.9600 ;
        RECT 1015.5800 755.7200 1017.1800 756.2000 ;
        RECT 1015.5800 761.1600 1017.1800 761.6400 ;
        RECT 1053.2000 739.4000 1054.8000 739.8800 ;
        RECT 1053.2000 744.8400 1054.8000 745.3200 ;
        RECT 1053.2000 750.2800 1054.8000 750.7600 ;
        RECT 1053.2000 728.5200 1054.8000 729.0000 ;
        RECT 1053.2000 733.9600 1054.8000 734.4400 ;
        RECT 1053.2000 712.2000 1054.8000 712.6800 ;
        RECT 1053.2000 717.6400 1054.8000 718.1200 ;
        RECT 1053.2000 723.0800 1054.8000 723.5600 ;
        RECT 1053.2000 701.3200 1054.8000 701.8000 ;
        RECT 1053.2000 706.7600 1054.8000 707.2400 ;
        RECT 1053.2000 685.0000 1054.8000 685.4800 ;
        RECT 1053.2000 690.4400 1054.8000 690.9200 ;
        RECT 1053.2000 695.8800 1054.8000 696.3600 ;
        RECT 1053.2000 674.1200 1054.8000 674.6000 ;
        RECT 1053.2000 679.5600 1054.8000 680.0400 ;
        RECT 1053.2000 657.8000 1054.8000 658.2800 ;
        RECT 1053.2000 663.2400 1054.8000 663.7200 ;
        RECT 1053.2000 668.6800 1054.8000 669.1600 ;
        RECT 1053.2000 652.3600 1054.8000 652.8400 ;
        RECT 1015.5800 739.4000 1017.1800 739.8800 ;
        RECT 1015.5800 744.8400 1017.1800 745.3200 ;
        RECT 1015.5800 750.2800 1017.1800 750.7600 ;
        RECT 1015.5800 728.5200 1017.1800 729.0000 ;
        RECT 1015.5800 733.9600 1017.1800 734.4400 ;
        RECT 1015.5800 712.2000 1017.1800 712.6800 ;
        RECT 1015.5800 717.6400 1017.1800 718.1200 ;
        RECT 1015.5800 723.0800 1017.1800 723.5600 ;
        RECT 1015.5800 701.3200 1017.1800 701.8000 ;
        RECT 1015.5800 706.7600 1017.1800 707.2400 ;
        RECT 1015.5800 685.0000 1017.1800 685.4800 ;
        RECT 1015.5800 690.4400 1017.1800 690.9200 ;
        RECT 1015.5800 695.8800 1017.1800 696.3600 ;
        RECT 1015.5800 674.1200 1017.1800 674.6000 ;
        RECT 1015.5800 679.5600 1017.1800 680.0400 ;
        RECT 1015.5800 657.8000 1017.1800 658.2800 ;
        RECT 1015.5800 663.2400 1017.1800 663.7200 ;
        RECT 1015.5800 668.6800 1017.1800 669.1600 ;
        RECT 1015.5800 652.3600 1017.1800 652.8400 ;
        RECT 1010.1200 854.7700 1060.2600 856.3700 ;
        RECT 1010.1200 648.0700 1060.2600 649.6700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 642.7400 1017.1800 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 860.7800 1017.1800 862.3800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 642.7400 1054.8000 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 860.7800 1054.8000 862.3800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 648.0700 1011.7200 649.6700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 648.0700 1060.2600 649.6700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 854.7700 1011.7200 856.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 854.7700 1060.2600 856.3700 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'W_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 1053.2000 413.1000 1054.8000 632.7400 ;
        RECT 1015.5800 413.1000 1017.1800 632.7400 ;
      LAYER met3 ;
        RECT 1053.2000 607.6800 1054.8000 608.1600 ;
        RECT 1053.2000 613.1200 1054.8000 613.6000 ;
        RECT 1053.2000 618.5600 1054.8000 619.0400 ;
        RECT 1053.2000 596.8000 1054.8000 597.2800 ;
        RECT 1053.2000 602.2400 1054.8000 602.7200 ;
        RECT 1053.2000 580.4800 1054.8000 580.9600 ;
        RECT 1053.2000 585.9200 1054.8000 586.4000 ;
        RECT 1053.2000 591.3600 1054.8000 591.8400 ;
        RECT 1053.2000 564.1600 1054.8000 564.6400 ;
        RECT 1053.2000 569.6000 1054.8000 570.0800 ;
        RECT 1053.2000 575.0400 1054.8000 575.5200 ;
        RECT 1053.2000 553.2800 1054.8000 553.7600 ;
        RECT 1053.2000 558.7200 1054.8000 559.2000 ;
        RECT 1053.2000 536.9600 1054.8000 537.4400 ;
        RECT 1053.2000 542.4000 1054.8000 542.8800 ;
        RECT 1053.2000 547.8400 1054.8000 548.3200 ;
        RECT 1053.2000 526.0800 1054.8000 526.5600 ;
        RECT 1053.2000 531.5200 1054.8000 532.0000 ;
        RECT 1015.5800 607.6800 1017.1800 608.1600 ;
        RECT 1015.5800 613.1200 1017.1800 613.6000 ;
        RECT 1015.5800 618.5600 1017.1800 619.0400 ;
        RECT 1015.5800 596.8000 1017.1800 597.2800 ;
        RECT 1015.5800 602.2400 1017.1800 602.7200 ;
        RECT 1015.5800 580.4800 1017.1800 580.9600 ;
        RECT 1015.5800 585.9200 1017.1800 586.4000 ;
        RECT 1015.5800 591.3600 1017.1800 591.8400 ;
        RECT 1015.5800 564.1600 1017.1800 564.6400 ;
        RECT 1015.5800 569.6000 1017.1800 570.0800 ;
        RECT 1015.5800 575.0400 1017.1800 575.5200 ;
        RECT 1015.5800 553.2800 1017.1800 553.7600 ;
        RECT 1015.5800 558.7200 1017.1800 559.2000 ;
        RECT 1015.5800 536.9600 1017.1800 537.4400 ;
        RECT 1015.5800 542.4000 1017.1800 542.8800 ;
        RECT 1015.5800 547.8400 1017.1800 548.3200 ;
        RECT 1015.5800 526.0800 1017.1800 526.5600 ;
        RECT 1015.5800 531.5200 1017.1800 532.0000 ;
        RECT 1053.2000 509.7600 1054.8000 510.2400 ;
        RECT 1053.2000 515.2000 1054.8000 515.6800 ;
        RECT 1053.2000 520.6400 1054.8000 521.1200 ;
        RECT 1053.2000 498.8800 1054.8000 499.3600 ;
        RECT 1053.2000 504.3200 1054.8000 504.8000 ;
        RECT 1053.2000 482.5600 1054.8000 483.0400 ;
        RECT 1053.2000 488.0000 1054.8000 488.4800 ;
        RECT 1053.2000 493.4400 1054.8000 493.9200 ;
        RECT 1053.2000 471.6800 1054.8000 472.1600 ;
        RECT 1053.2000 477.1200 1054.8000 477.6000 ;
        RECT 1053.2000 455.3600 1054.8000 455.8400 ;
        RECT 1053.2000 460.8000 1054.8000 461.2800 ;
        RECT 1053.2000 466.2400 1054.8000 466.7200 ;
        RECT 1053.2000 444.4800 1054.8000 444.9600 ;
        RECT 1053.2000 449.9200 1054.8000 450.4000 ;
        RECT 1053.2000 428.1600 1054.8000 428.6400 ;
        RECT 1053.2000 433.6000 1054.8000 434.0800 ;
        RECT 1053.2000 439.0400 1054.8000 439.5200 ;
        RECT 1053.2000 422.7200 1054.8000 423.2000 ;
        RECT 1015.5800 509.7600 1017.1800 510.2400 ;
        RECT 1015.5800 515.2000 1017.1800 515.6800 ;
        RECT 1015.5800 520.6400 1017.1800 521.1200 ;
        RECT 1015.5800 498.8800 1017.1800 499.3600 ;
        RECT 1015.5800 504.3200 1017.1800 504.8000 ;
        RECT 1015.5800 482.5600 1017.1800 483.0400 ;
        RECT 1015.5800 488.0000 1017.1800 488.4800 ;
        RECT 1015.5800 493.4400 1017.1800 493.9200 ;
        RECT 1015.5800 471.6800 1017.1800 472.1600 ;
        RECT 1015.5800 477.1200 1017.1800 477.6000 ;
        RECT 1015.5800 455.3600 1017.1800 455.8400 ;
        RECT 1015.5800 460.8000 1017.1800 461.2800 ;
        RECT 1015.5800 466.2400 1017.1800 466.7200 ;
        RECT 1015.5800 444.4800 1017.1800 444.9600 ;
        RECT 1015.5800 449.9200 1017.1800 450.4000 ;
        RECT 1015.5800 428.1600 1017.1800 428.6400 ;
        RECT 1015.5800 433.6000 1017.1800 434.0800 ;
        RECT 1015.5800 439.0400 1017.1800 439.5200 ;
        RECT 1015.5800 422.7200 1017.1800 423.2000 ;
        RECT 1010.1200 625.1300 1060.2600 626.7300 ;
        RECT 1010.1200 418.4300 1060.2600 420.0300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 413.1000 1017.1800 414.7000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1015.5800 631.1400 1017.1800 632.7400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 413.1000 1054.8000 414.7000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1053.2000 631.1400 1054.8000 632.7400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 418.4300 1011.7200 420.0300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 418.4300 1060.2600 420.0300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1010.1200 625.1300 1011.7200 626.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1058.6600 625.1300 1060.2600 626.7300 ;
    END
# end of P/G pin shape extracted from block 'W_CPU_IO'


# P/G pin shape extracted from block 'N_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1075.5800 2479.6000 1077.1800 2509.8600 ;
        RECT 1273.2800 2479.6000 1274.8800 2509.8600 ;
      LAYER met3 ;
        RECT 1273.2800 2497.3800 1274.8800 2497.8600 ;
        RECT 1075.5800 2497.3800 1077.1800 2497.8600 ;
        RECT 1273.2800 2491.9400 1274.8800 2492.4200 ;
        RECT 1273.2800 2486.5000 1274.8800 2486.9800 ;
        RECT 1075.5800 2491.9400 1077.1800 2492.4200 ;
        RECT 1075.5800 2486.5000 1077.1800 2486.9800 ;
        RECT 1070.1200 2503.1000 1280.3400 2504.7000 ;
        RECT 1070.1200 2483.5700 1280.3400 2485.1700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.5800 2479.6000 1077.1800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.5800 2508.2600 1077.1800 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.2800 2479.6000 1274.8800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.2800 2508.2600 1274.8800 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.1200 2483.5700 1071.7200 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.7400 2483.5700 1280.3400 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.1200 2503.1000 1071.7200 2504.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.7400 2503.1000 1280.3400 2504.7000 ;
    END
# end of P/G pin shape extracted from block 'N_term_DSP'


# P/G pin shape extracted from block 'S_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1075.7200 143.2000 1077.3200 173.4600 ;
        RECT 1273.4200 143.2000 1275.0200 173.4600 ;
      LAYER met3 ;
        RECT 1273.4200 160.9800 1275.0200 161.4600 ;
        RECT 1075.7200 160.9800 1077.3200 161.4600 ;
        RECT 1273.4200 155.5400 1275.0200 156.0200 ;
        RECT 1273.4200 150.1000 1275.0200 150.5800 ;
        RECT 1075.7200 155.5400 1077.3200 156.0200 ;
        RECT 1075.7200 150.1000 1077.3200 150.5800 ;
        RECT 1070.2600 166.7000 1280.4800 168.3000 ;
        RECT 1070.2600 147.1700 1280.4800 148.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.7200 143.2000 1077.3200 144.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.7200 171.8600 1077.3200 173.4600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.4200 143.2000 1275.0200 144.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.4200 171.8600 1275.0200 173.4600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 147.1700 1071.8600 148.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 147.1700 1280.4800 148.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 166.7000 1071.8600 168.3000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 166.7000 1280.4800 168.3000 ;
    END
# end of P/G pin shape extracted from block 'S_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1075.8200 2020.5800 1077.4200 2470.4000 ;
        RECT 1273.3200 2020.5800 1274.9200 2470.4000 ;
        RECT 1083.5800 2026.0100 1085.1800 2464.8000 ;
        RECT 1128.5800 2026.0100 1130.1800 2464.8000 ;
        RECT 1173.5800 2026.0100 1175.1800 2464.8000 ;
        RECT 1218.5800 2026.0100 1220.1800 2464.8000 ;
        RECT 1263.5800 2026.0100 1265.1800 2464.8000 ;
      LAYER met3 ;
        RECT 1273.3200 2459.9600 1274.9200 2460.4400 ;
        RECT 1273.3200 2454.5200 1274.9200 2455.0000 ;
        RECT 1273.3200 2449.0800 1274.9200 2449.5600 ;
        RECT 1273.3200 2443.6400 1274.9200 2444.1200 ;
        RECT 1273.3200 2438.2000 1274.9200 2438.6800 ;
        RECT 1273.3200 2432.7600 1274.9200 2433.2400 ;
        RECT 1273.3200 2427.3200 1274.9200 2427.8000 ;
        RECT 1273.3200 2421.8800 1274.9200 2422.3600 ;
        RECT 1273.3200 2416.4400 1274.9200 2416.9200 ;
        RECT 1273.3200 2411.0000 1274.9200 2411.4800 ;
        RECT 1273.3200 2405.5600 1274.9200 2406.0400 ;
        RECT 1273.3200 2400.1200 1274.9200 2400.6000 ;
        RECT 1273.3200 2394.6800 1274.9200 2395.1600 ;
        RECT 1273.3200 2389.2400 1274.9200 2389.7200 ;
        RECT 1273.3200 2383.8000 1274.9200 2384.2800 ;
        RECT 1273.3200 2378.3600 1274.9200 2378.8400 ;
        RECT 1273.3200 2372.9200 1274.9200 2373.4000 ;
        RECT 1273.3200 2367.4800 1274.9200 2367.9600 ;
        RECT 1273.3200 2362.0400 1274.9200 2362.5200 ;
        RECT 1273.3200 2356.6000 1274.9200 2357.0800 ;
        RECT 1273.3200 2351.1600 1274.9200 2351.6400 ;
        RECT 1273.3200 2345.7200 1274.9200 2346.2000 ;
        RECT 1273.3200 2340.2800 1274.9200 2340.7600 ;
        RECT 1273.3200 2334.8400 1274.9200 2335.3200 ;
        RECT 1273.3200 2323.9600 1274.9200 2324.4400 ;
        RECT 1273.3200 2318.5200 1274.9200 2319.0000 ;
        RECT 1273.3200 2313.0800 1274.9200 2313.5600 ;
        RECT 1273.3200 2307.6400 1274.9200 2308.1200 ;
        RECT 1273.3200 2302.2000 1274.9200 2302.6800 ;
        RECT 1273.3200 2329.4000 1274.9200 2329.8800 ;
        RECT 1273.3200 2296.7600 1274.9200 2297.2400 ;
        RECT 1273.3200 2291.3200 1274.9200 2291.8000 ;
        RECT 1273.3200 2285.8800 1274.9200 2286.3600 ;
        RECT 1273.3200 2280.4400 1274.9200 2280.9200 ;
        RECT 1273.3200 2275.0000 1274.9200 2275.4800 ;
        RECT 1273.3200 2269.5600 1274.9200 2270.0400 ;
        RECT 1273.3200 2264.1200 1274.9200 2264.6000 ;
        RECT 1273.3200 2258.6800 1274.9200 2259.1600 ;
        RECT 1273.3200 2253.2400 1274.9200 2253.7200 ;
        RECT 1273.3200 2247.8000 1274.9200 2248.2800 ;
        RECT 1075.8200 2459.9600 1077.4200 2460.4400 ;
        RECT 1075.8200 2454.5200 1077.4200 2455.0000 ;
        RECT 1075.8200 2449.0800 1077.4200 2449.5600 ;
        RECT 1075.8200 2443.6400 1077.4200 2444.1200 ;
        RECT 1075.8200 2438.2000 1077.4200 2438.6800 ;
        RECT 1075.8200 2432.7600 1077.4200 2433.2400 ;
        RECT 1075.8200 2427.3200 1077.4200 2427.8000 ;
        RECT 1075.8200 2421.8800 1077.4200 2422.3600 ;
        RECT 1075.8200 2416.4400 1077.4200 2416.9200 ;
        RECT 1075.8200 2411.0000 1077.4200 2411.4800 ;
        RECT 1075.8200 2405.5600 1077.4200 2406.0400 ;
        RECT 1075.8200 2400.1200 1077.4200 2400.6000 ;
        RECT 1075.8200 2394.6800 1077.4200 2395.1600 ;
        RECT 1075.8200 2389.2400 1077.4200 2389.7200 ;
        RECT 1075.8200 2383.8000 1077.4200 2384.2800 ;
        RECT 1075.8200 2378.3600 1077.4200 2378.8400 ;
        RECT 1075.8200 2372.9200 1077.4200 2373.4000 ;
        RECT 1075.8200 2367.4800 1077.4200 2367.9600 ;
        RECT 1075.8200 2362.0400 1077.4200 2362.5200 ;
        RECT 1075.8200 2356.6000 1077.4200 2357.0800 ;
        RECT 1075.8200 2351.1600 1077.4200 2351.6400 ;
        RECT 1075.8200 2345.7200 1077.4200 2346.2000 ;
        RECT 1075.8200 2340.2800 1077.4200 2340.7600 ;
        RECT 1075.8200 2334.8400 1077.4200 2335.3200 ;
        RECT 1075.8200 2323.9600 1077.4200 2324.4400 ;
        RECT 1075.8200 2318.5200 1077.4200 2319.0000 ;
        RECT 1075.8200 2313.0800 1077.4200 2313.5600 ;
        RECT 1075.8200 2307.6400 1077.4200 2308.1200 ;
        RECT 1075.8200 2302.2000 1077.4200 2302.6800 ;
        RECT 1075.8200 2329.4000 1077.4200 2329.8800 ;
        RECT 1075.8200 2296.7600 1077.4200 2297.2400 ;
        RECT 1075.8200 2291.3200 1077.4200 2291.8000 ;
        RECT 1075.8200 2285.8800 1077.4200 2286.3600 ;
        RECT 1075.8200 2280.4400 1077.4200 2280.9200 ;
        RECT 1075.8200 2275.0000 1077.4200 2275.4800 ;
        RECT 1075.8200 2269.5600 1077.4200 2270.0400 ;
        RECT 1075.8200 2264.1200 1077.4200 2264.6000 ;
        RECT 1075.8200 2258.6800 1077.4200 2259.1600 ;
        RECT 1075.8200 2253.2400 1077.4200 2253.7200 ;
        RECT 1075.8200 2247.8000 1077.4200 2248.2800 ;
        RECT 1273.3200 2242.3600 1274.9200 2242.8400 ;
        RECT 1273.3200 2236.9200 1274.9200 2237.4000 ;
        RECT 1273.3200 2231.4800 1274.9200 2231.9600 ;
        RECT 1273.3200 2226.0400 1274.9200 2226.5200 ;
        RECT 1273.3200 2220.6000 1274.9200 2221.0800 ;
        RECT 1273.3200 2215.1600 1274.9200 2215.6400 ;
        RECT 1273.3200 2209.7200 1274.9200 2210.2000 ;
        RECT 1273.3200 2204.2800 1274.9200 2204.7600 ;
        RECT 1273.3200 2198.8400 1274.9200 2199.3200 ;
        RECT 1273.3200 2193.4000 1274.9200 2193.8800 ;
        RECT 1273.3200 2187.9600 1274.9200 2188.4400 ;
        RECT 1273.3200 2182.5200 1274.9200 2183.0000 ;
        RECT 1273.3200 2177.0800 1274.9200 2177.5600 ;
        RECT 1273.3200 2171.6400 1274.9200 2172.1200 ;
        RECT 1273.3200 2166.2000 1274.9200 2166.6800 ;
        RECT 1273.3200 2155.3200 1274.9200 2155.8000 ;
        RECT 1273.3200 2149.8800 1274.9200 2150.3600 ;
        RECT 1273.3200 2144.4400 1274.9200 2144.9200 ;
        RECT 1273.3200 2139.0000 1274.9200 2139.4800 ;
        RECT 1273.3200 2133.5600 1274.9200 2134.0400 ;
        RECT 1273.3200 2160.7600 1274.9200 2161.2400 ;
        RECT 1273.3200 2128.1200 1274.9200 2128.6000 ;
        RECT 1273.3200 2122.6800 1274.9200 2123.1600 ;
        RECT 1273.3200 2117.2400 1274.9200 2117.7200 ;
        RECT 1273.3200 2111.8000 1274.9200 2112.2800 ;
        RECT 1273.3200 2106.3600 1274.9200 2106.8400 ;
        RECT 1273.3200 2100.9200 1274.9200 2101.4000 ;
        RECT 1273.3200 2095.4800 1274.9200 2095.9600 ;
        RECT 1273.3200 2090.0400 1274.9200 2090.5200 ;
        RECT 1273.3200 2084.6000 1274.9200 2085.0800 ;
        RECT 1273.3200 2079.1600 1274.9200 2079.6400 ;
        RECT 1273.3200 2073.7200 1274.9200 2074.2000 ;
        RECT 1273.3200 2068.2800 1274.9200 2068.7600 ;
        RECT 1273.3200 2062.8400 1274.9200 2063.3200 ;
        RECT 1273.3200 2057.4000 1274.9200 2057.8800 ;
        RECT 1273.3200 2051.9600 1274.9200 2052.4400 ;
        RECT 1273.3200 2046.5200 1274.9200 2047.0000 ;
        RECT 1273.3200 2041.0800 1274.9200 2041.5600 ;
        RECT 1273.3200 2035.6400 1274.9200 2036.1200 ;
        RECT 1273.3200 2030.2000 1274.9200 2030.6800 ;
        RECT 1075.8200 2242.3600 1077.4200 2242.8400 ;
        RECT 1075.8200 2236.9200 1077.4200 2237.4000 ;
        RECT 1075.8200 2231.4800 1077.4200 2231.9600 ;
        RECT 1075.8200 2226.0400 1077.4200 2226.5200 ;
        RECT 1075.8200 2220.6000 1077.4200 2221.0800 ;
        RECT 1075.8200 2215.1600 1077.4200 2215.6400 ;
        RECT 1075.8200 2209.7200 1077.4200 2210.2000 ;
        RECT 1075.8200 2204.2800 1077.4200 2204.7600 ;
        RECT 1075.8200 2198.8400 1077.4200 2199.3200 ;
        RECT 1075.8200 2193.4000 1077.4200 2193.8800 ;
        RECT 1075.8200 2187.9600 1077.4200 2188.4400 ;
        RECT 1075.8200 2182.5200 1077.4200 2183.0000 ;
        RECT 1075.8200 2177.0800 1077.4200 2177.5600 ;
        RECT 1075.8200 2171.6400 1077.4200 2172.1200 ;
        RECT 1075.8200 2166.2000 1077.4200 2166.6800 ;
        RECT 1075.8200 2155.3200 1077.4200 2155.8000 ;
        RECT 1075.8200 2149.8800 1077.4200 2150.3600 ;
        RECT 1075.8200 2144.4400 1077.4200 2144.9200 ;
        RECT 1075.8200 2139.0000 1077.4200 2139.4800 ;
        RECT 1075.8200 2133.5600 1077.4200 2134.0400 ;
        RECT 1075.8200 2160.7600 1077.4200 2161.2400 ;
        RECT 1075.8200 2128.1200 1077.4200 2128.6000 ;
        RECT 1075.8200 2122.6800 1077.4200 2123.1600 ;
        RECT 1075.8200 2117.2400 1077.4200 2117.7200 ;
        RECT 1075.8200 2111.8000 1077.4200 2112.2800 ;
        RECT 1075.8200 2106.3600 1077.4200 2106.8400 ;
        RECT 1075.8200 2100.9200 1077.4200 2101.4000 ;
        RECT 1075.8200 2095.4800 1077.4200 2095.9600 ;
        RECT 1075.8200 2090.0400 1077.4200 2090.5200 ;
        RECT 1075.8200 2084.6000 1077.4200 2085.0800 ;
        RECT 1075.8200 2079.1600 1077.4200 2079.6400 ;
        RECT 1075.8200 2073.7200 1077.4200 2074.2000 ;
        RECT 1075.8200 2068.2800 1077.4200 2068.7600 ;
        RECT 1075.8200 2062.8400 1077.4200 2063.3200 ;
        RECT 1075.8200 2057.4000 1077.4200 2057.8800 ;
        RECT 1075.8200 2051.9600 1077.4200 2052.4400 ;
        RECT 1075.8200 2046.5200 1077.4200 2047.0000 ;
        RECT 1075.8200 2041.0800 1077.4200 2041.5600 ;
        RECT 1075.8200 2035.6400 1077.4200 2036.1200 ;
        RECT 1075.8200 2030.2000 1077.4200 2030.6800 ;
        RECT 1070.2600 2463.2000 1280.4800 2464.8000 ;
        RECT 1070.2600 2026.0100 1280.4800 2027.6100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 2020.5800 1077.4200 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 2468.8000 1077.4200 2470.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 2020.5800 1274.9200 2022.1800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 2468.8000 1274.9200 2470.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 2026.0100 1071.8600 2027.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 2026.0100 1280.4800 2027.6100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 2463.2000 1071.8600 2464.8000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 2463.2000 1280.4800 2464.8000 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1075.8200 1561.3000 1077.4200 2011.1200 ;
        RECT 1273.3200 1561.3000 1274.9200 2011.1200 ;
        RECT 1083.5800 1566.7300 1085.1800 2005.5200 ;
        RECT 1128.5800 1566.7300 1130.1800 2005.5200 ;
        RECT 1173.5800 1566.7300 1175.1800 2005.5200 ;
        RECT 1218.5800 1566.7300 1220.1800 2005.5200 ;
        RECT 1263.5800 1566.7300 1265.1800 2005.5200 ;
      LAYER met3 ;
        RECT 1273.3200 2000.6800 1274.9200 2001.1600 ;
        RECT 1273.3200 1995.2400 1274.9200 1995.7200 ;
        RECT 1273.3200 1989.8000 1274.9200 1990.2800 ;
        RECT 1273.3200 1984.3600 1274.9200 1984.8400 ;
        RECT 1273.3200 1978.9200 1274.9200 1979.4000 ;
        RECT 1273.3200 1973.4800 1274.9200 1973.9600 ;
        RECT 1273.3200 1968.0400 1274.9200 1968.5200 ;
        RECT 1273.3200 1962.6000 1274.9200 1963.0800 ;
        RECT 1273.3200 1957.1600 1274.9200 1957.6400 ;
        RECT 1273.3200 1951.7200 1274.9200 1952.2000 ;
        RECT 1273.3200 1946.2800 1274.9200 1946.7600 ;
        RECT 1273.3200 1940.8400 1274.9200 1941.3200 ;
        RECT 1273.3200 1935.4000 1274.9200 1935.8800 ;
        RECT 1273.3200 1929.9600 1274.9200 1930.4400 ;
        RECT 1273.3200 1924.5200 1274.9200 1925.0000 ;
        RECT 1273.3200 1919.0800 1274.9200 1919.5600 ;
        RECT 1273.3200 1913.6400 1274.9200 1914.1200 ;
        RECT 1273.3200 1908.2000 1274.9200 1908.6800 ;
        RECT 1273.3200 1902.7600 1274.9200 1903.2400 ;
        RECT 1273.3200 1897.3200 1274.9200 1897.8000 ;
        RECT 1273.3200 1891.8800 1274.9200 1892.3600 ;
        RECT 1273.3200 1886.4400 1274.9200 1886.9200 ;
        RECT 1273.3200 1881.0000 1274.9200 1881.4800 ;
        RECT 1273.3200 1875.5600 1274.9200 1876.0400 ;
        RECT 1273.3200 1864.6800 1274.9200 1865.1600 ;
        RECT 1273.3200 1859.2400 1274.9200 1859.7200 ;
        RECT 1273.3200 1853.8000 1274.9200 1854.2800 ;
        RECT 1273.3200 1848.3600 1274.9200 1848.8400 ;
        RECT 1273.3200 1842.9200 1274.9200 1843.4000 ;
        RECT 1273.3200 1870.1200 1274.9200 1870.6000 ;
        RECT 1273.3200 1837.4800 1274.9200 1837.9600 ;
        RECT 1273.3200 1832.0400 1274.9200 1832.5200 ;
        RECT 1273.3200 1826.6000 1274.9200 1827.0800 ;
        RECT 1273.3200 1821.1600 1274.9200 1821.6400 ;
        RECT 1273.3200 1815.7200 1274.9200 1816.2000 ;
        RECT 1273.3200 1810.2800 1274.9200 1810.7600 ;
        RECT 1273.3200 1804.8400 1274.9200 1805.3200 ;
        RECT 1273.3200 1799.4000 1274.9200 1799.8800 ;
        RECT 1273.3200 1793.9600 1274.9200 1794.4400 ;
        RECT 1273.3200 1788.5200 1274.9200 1789.0000 ;
        RECT 1075.8200 2000.6800 1077.4200 2001.1600 ;
        RECT 1075.8200 1995.2400 1077.4200 1995.7200 ;
        RECT 1075.8200 1989.8000 1077.4200 1990.2800 ;
        RECT 1075.8200 1984.3600 1077.4200 1984.8400 ;
        RECT 1075.8200 1978.9200 1077.4200 1979.4000 ;
        RECT 1075.8200 1973.4800 1077.4200 1973.9600 ;
        RECT 1075.8200 1968.0400 1077.4200 1968.5200 ;
        RECT 1075.8200 1962.6000 1077.4200 1963.0800 ;
        RECT 1075.8200 1957.1600 1077.4200 1957.6400 ;
        RECT 1075.8200 1951.7200 1077.4200 1952.2000 ;
        RECT 1075.8200 1946.2800 1077.4200 1946.7600 ;
        RECT 1075.8200 1940.8400 1077.4200 1941.3200 ;
        RECT 1075.8200 1935.4000 1077.4200 1935.8800 ;
        RECT 1075.8200 1929.9600 1077.4200 1930.4400 ;
        RECT 1075.8200 1924.5200 1077.4200 1925.0000 ;
        RECT 1075.8200 1919.0800 1077.4200 1919.5600 ;
        RECT 1075.8200 1913.6400 1077.4200 1914.1200 ;
        RECT 1075.8200 1908.2000 1077.4200 1908.6800 ;
        RECT 1075.8200 1902.7600 1077.4200 1903.2400 ;
        RECT 1075.8200 1897.3200 1077.4200 1897.8000 ;
        RECT 1075.8200 1891.8800 1077.4200 1892.3600 ;
        RECT 1075.8200 1886.4400 1077.4200 1886.9200 ;
        RECT 1075.8200 1881.0000 1077.4200 1881.4800 ;
        RECT 1075.8200 1875.5600 1077.4200 1876.0400 ;
        RECT 1075.8200 1864.6800 1077.4200 1865.1600 ;
        RECT 1075.8200 1859.2400 1077.4200 1859.7200 ;
        RECT 1075.8200 1853.8000 1077.4200 1854.2800 ;
        RECT 1075.8200 1848.3600 1077.4200 1848.8400 ;
        RECT 1075.8200 1842.9200 1077.4200 1843.4000 ;
        RECT 1075.8200 1870.1200 1077.4200 1870.6000 ;
        RECT 1075.8200 1837.4800 1077.4200 1837.9600 ;
        RECT 1075.8200 1832.0400 1077.4200 1832.5200 ;
        RECT 1075.8200 1826.6000 1077.4200 1827.0800 ;
        RECT 1075.8200 1821.1600 1077.4200 1821.6400 ;
        RECT 1075.8200 1815.7200 1077.4200 1816.2000 ;
        RECT 1075.8200 1810.2800 1077.4200 1810.7600 ;
        RECT 1075.8200 1804.8400 1077.4200 1805.3200 ;
        RECT 1075.8200 1799.4000 1077.4200 1799.8800 ;
        RECT 1075.8200 1793.9600 1077.4200 1794.4400 ;
        RECT 1075.8200 1788.5200 1077.4200 1789.0000 ;
        RECT 1273.3200 1783.0800 1274.9200 1783.5600 ;
        RECT 1273.3200 1777.6400 1274.9200 1778.1200 ;
        RECT 1273.3200 1772.2000 1274.9200 1772.6800 ;
        RECT 1273.3200 1766.7600 1274.9200 1767.2400 ;
        RECT 1273.3200 1761.3200 1274.9200 1761.8000 ;
        RECT 1273.3200 1755.8800 1274.9200 1756.3600 ;
        RECT 1273.3200 1750.4400 1274.9200 1750.9200 ;
        RECT 1273.3200 1745.0000 1274.9200 1745.4800 ;
        RECT 1273.3200 1739.5600 1274.9200 1740.0400 ;
        RECT 1273.3200 1734.1200 1274.9200 1734.6000 ;
        RECT 1273.3200 1728.6800 1274.9200 1729.1600 ;
        RECT 1273.3200 1723.2400 1274.9200 1723.7200 ;
        RECT 1273.3200 1717.8000 1274.9200 1718.2800 ;
        RECT 1273.3200 1712.3600 1274.9200 1712.8400 ;
        RECT 1273.3200 1706.9200 1274.9200 1707.4000 ;
        RECT 1273.3200 1696.0400 1274.9200 1696.5200 ;
        RECT 1273.3200 1690.6000 1274.9200 1691.0800 ;
        RECT 1273.3200 1685.1600 1274.9200 1685.6400 ;
        RECT 1273.3200 1679.7200 1274.9200 1680.2000 ;
        RECT 1273.3200 1674.2800 1274.9200 1674.7600 ;
        RECT 1273.3200 1701.4800 1274.9200 1701.9600 ;
        RECT 1273.3200 1668.8400 1274.9200 1669.3200 ;
        RECT 1273.3200 1663.4000 1274.9200 1663.8800 ;
        RECT 1273.3200 1657.9600 1274.9200 1658.4400 ;
        RECT 1273.3200 1652.5200 1274.9200 1653.0000 ;
        RECT 1273.3200 1647.0800 1274.9200 1647.5600 ;
        RECT 1273.3200 1641.6400 1274.9200 1642.1200 ;
        RECT 1273.3200 1636.2000 1274.9200 1636.6800 ;
        RECT 1273.3200 1630.7600 1274.9200 1631.2400 ;
        RECT 1273.3200 1625.3200 1274.9200 1625.8000 ;
        RECT 1273.3200 1619.8800 1274.9200 1620.3600 ;
        RECT 1273.3200 1614.4400 1274.9200 1614.9200 ;
        RECT 1273.3200 1609.0000 1274.9200 1609.4800 ;
        RECT 1273.3200 1603.5600 1274.9200 1604.0400 ;
        RECT 1273.3200 1598.1200 1274.9200 1598.6000 ;
        RECT 1273.3200 1592.6800 1274.9200 1593.1600 ;
        RECT 1273.3200 1587.2400 1274.9200 1587.7200 ;
        RECT 1273.3200 1581.8000 1274.9200 1582.2800 ;
        RECT 1273.3200 1576.3600 1274.9200 1576.8400 ;
        RECT 1273.3200 1570.9200 1274.9200 1571.4000 ;
        RECT 1075.8200 1783.0800 1077.4200 1783.5600 ;
        RECT 1075.8200 1777.6400 1077.4200 1778.1200 ;
        RECT 1075.8200 1772.2000 1077.4200 1772.6800 ;
        RECT 1075.8200 1766.7600 1077.4200 1767.2400 ;
        RECT 1075.8200 1761.3200 1077.4200 1761.8000 ;
        RECT 1075.8200 1755.8800 1077.4200 1756.3600 ;
        RECT 1075.8200 1750.4400 1077.4200 1750.9200 ;
        RECT 1075.8200 1745.0000 1077.4200 1745.4800 ;
        RECT 1075.8200 1739.5600 1077.4200 1740.0400 ;
        RECT 1075.8200 1734.1200 1077.4200 1734.6000 ;
        RECT 1075.8200 1728.6800 1077.4200 1729.1600 ;
        RECT 1075.8200 1723.2400 1077.4200 1723.7200 ;
        RECT 1075.8200 1717.8000 1077.4200 1718.2800 ;
        RECT 1075.8200 1712.3600 1077.4200 1712.8400 ;
        RECT 1075.8200 1706.9200 1077.4200 1707.4000 ;
        RECT 1075.8200 1696.0400 1077.4200 1696.5200 ;
        RECT 1075.8200 1690.6000 1077.4200 1691.0800 ;
        RECT 1075.8200 1685.1600 1077.4200 1685.6400 ;
        RECT 1075.8200 1679.7200 1077.4200 1680.2000 ;
        RECT 1075.8200 1674.2800 1077.4200 1674.7600 ;
        RECT 1075.8200 1701.4800 1077.4200 1701.9600 ;
        RECT 1075.8200 1668.8400 1077.4200 1669.3200 ;
        RECT 1075.8200 1663.4000 1077.4200 1663.8800 ;
        RECT 1075.8200 1657.9600 1077.4200 1658.4400 ;
        RECT 1075.8200 1652.5200 1077.4200 1653.0000 ;
        RECT 1075.8200 1647.0800 1077.4200 1647.5600 ;
        RECT 1075.8200 1641.6400 1077.4200 1642.1200 ;
        RECT 1075.8200 1636.2000 1077.4200 1636.6800 ;
        RECT 1075.8200 1630.7600 1077.4200 1631.2400 ;
        RECT 1075.8200 1625.3200 1077.4200 1625.8000 ;
        RECT 1075.8200 1619.8800 1077.4200 1620.3600 ;
        RECT 1075.8200 1614.4400 1077.4200 1614.9200 ;
        RECT 1075.8200 1609.0000 1077.4200 1609.4800 ;
        RECT 1075.8200 1603.5600 1077.4200 1604.0400 ;
        RECT 1075.8200 1598.1200 1077.4200 1598.6000 ;
        RECT 1075.8200 1592.6800 1077.4200 1593.1600 ;
        RECT 1075.8200 1587.2400 1077.4200 1587.7200 ;
        RECT 1075.8200 1581.8000 1077.4200 1582.2800 ;
        RECT 1075.8200 1576.3600 1077.4200 1576.8400 ;
        RECT 1075.8200 1570.9200 1077.4200 1571.4000 ;
        RECT 1070.2600 2003.9200 1280.4800 2005.5200 ;
        RECT 1070.2600 1566.7300 1280.4800 1568.3300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 1561.3000 1077.4200 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 2009.5200 1077.4200 2011.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 1561.3000 1274.9200 1562.9000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 2009.5200 1274.9200 2011.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1566.7300 1071.8600 1568.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1566.7300 1280.4800 1568.3300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 2003.9200 1071.8600 2005.5200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 2003.9200 1280.4800 2005.5200 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1075.8200 1102.0200 1077.4200 1551.8400 ;
        RECT 1273.3200 1102.0200 1274.9200 1551.8400 ;
        RECT 1083.5800 1107.4500 1085.1800 1546.2400 ;
        RECT 1128.5800 1107.4500 1130.1800 1546.2400 ;
        RECT 1173.5800 1107.4500 1175.1800 1546.2400 ;
        RECT 1218.5800 1107.4500 1220.1800 1546.2400 ;
        RECT 1263.5800 1107.4500 1265.1800 1546.2400 ;
      LAYER met3 ;
        RECT 1273.3200 1541.4000 1274.9200 1541.8800 ;
        RECT 1273.3200 1535.9600 1274.9200 1536.4400 ;
        RECT 1273.3200 1530.5200 1274.9200 1531.0000 ;
        RECT 1273.3200 1525.0800 1274.9200 1525.5600 ;
        RECT 1273.3200 1519.6400 1274.9200 1520.1200 ;
        RECT 1273.3200 1514.2000 1274.9200 1514.6800 ;
        RECT 1273.3200 1508.7600 1274.9200 1509.2400 ;
        RECT 1273.3200 1503.3200 1274.9200 1503.8000 ;
        RECT 1273.3200 1497.8800 1274.9200 1498.3600 ;
        RECT 1273.3200 1492.4400 1274.9200 1492.9200 ;
        RECT 1273.3200 1487.0000 1274.9200 1487.4800 ;
        RECT 1273.3200 1481.5600 1274.9200 1482.0400 ;
        RECT 1273.3200 1476.1200 1274.9200 1476.6000 ;
        RECT 1273.3200 1470.6800 1274.9200 1471.1600 ;
        RECT 1273.3200 1465.2400 1274.9200 1465.7200 ;
        RECT 1273.3200 1459.8000 1274.9200 1460.2800 ;
        RECT 1273.3200 1454.3600 1274.9200 1454.8400 ;
        RECT 1273.3200 1448.9200 1274.9200 1449.4000 ;
        RECT 1273.3200 1443.4800 1274.9200 1443.9600 ;
        RECT 1273.3200 1438.0400 1274.9200 1438.5200 ;
        RECT 1273.3200 1432.6000 1274.9200 1433.0800 ;
        RECT 1273.3200 1427.1600 1274.9200 1427.6400 ;
        RECT 1273.3200 1421.7200 1274.9200 1422.2000 ;
        RECT 1273.3200 1416.2800 1274.9200 1416.7600 ;
        RECT 1273.3200 1405.4000 1274.9200 1405.8800 ;
        RECT 1273.3200 1399.9600 1274.9200 1400.4400 ;
        RECT 1273.3200 1394.5200 1274.9200 1395.0000 ;
        RECT 1273.3200 1389.0800 1274.9200 1389.5600 ;
        RECT 1273.3200 1383.6400 1274.9200 1384.1200 ;
        RECT 1273.3200 1410.8400 1274.9200 1411.3200 ;
        RECT 1273.3200 1378.2000 1274.9200 1378.6800 ;
        RECT 1273.3200 1372.7600 1274.9200 1373.2400 ;
        RECT 1273.3200 1367.3200 1274.9200 1367.8000 ;
        RECT 1273.3200 1361.8800 1274.9200 1362.3600 ;
        RECT 1273.3200 1356.4400 1274.9200 1356.9200 ;
        RECT 1273.3200 1351.0000 1274.9200 1351.4800 ;
        RECT 1273.3200 1345.5600 1274.9200 1346.0400 ;
        RECT 1273.3200 1340.1200 1274.9200 1340.6000 ;
        RECT 1273.3200 1334.6800 1274.9200 1335.1600 ;
        RECT 1273.3200 1329.2400 1274.9200 1329.7200 ;
        RECT 1075.8200 1541.4000 1077.4200 1541.8800 ;
        RECT 1075.8200 1535.9600 1077.4200 1536.4400 ;
        RECT 1075.8200 1530.5200 1077.4200 1531.0000 ;
        RECT 1075.8200 1525.0800 1077.4200 1525.5600 ;
        RECT 1075.8200 1519.6400 1077.4200 1520.1200 ;
        RECT 1075.8200 1514.2000 1077.4200 1514.6800 ;
        RECT 1075.8200 1508.7600 1077.4200 1509.2400 ;
        RECT 1075.8200 1503.3200 1077.4200 1503.8000 ;
        RECT 1075.8200 1497.8800 1077.4200 1498.3600 ;
        RECT 1075.8200 1492.4400 1077.4200 1492.9200 ;
        RECT 1075.8200 1487.0000 1077.4200 1487.4800 ;
        RECT 1075.8200 1481.5600 1077.4200 1482.0400 ;
        RECT 1075.8200 1476.1200 1077.4200 1476.6000 ;
        RECT 1075.8200 1470.6800 1077.4200 1471.1600 ;
        RECT 1075.8200 1465.2400 1077.4200 1465.7200 ;
        RECT 1075.8200 1459.8000 1077.4200 1460.2800 ;
        RECT 1075.8200 1454.3600 1077.4200 1454.8400 ;
        RECT 1075.8200 1448.9200 1077.4200 1449.4000 ;
        RECT 1075.8200 1443.4800 1077.4200 1443.9600 ;
        RECT 1075.8200 1438.0400 1077.4200 1438.5200 ;
        RECT 1075.8200 1432.6000 1077.4200 1433.0800 ;
        RECT 1075.8200 1427.1600 1077.4200 1427.6400 ;
        RECT 1075.8200 1421.7200 1077.4200 1422.2000 ;
        RECT 1075.8200 1416.2800 1077.4200 1416.7600 ;
        RECT 1075.8200 1405.4000 1077.4200 1405.8800 ;
        RECT 1075.8200 1399.9600 1077.4200 1400.4400 ;
        RECT 1075.8200 1394.5200 1077.4200 1395.0000 ;
        RECT 1075.8200 1389.0800 1077.4200 1389.5600 ;
        RECT 1075.8200 1383.6400 1077.4200 1384.1200 ;
        RECT 1075.8200 1410.8400 1077.4200 1411.3200 ;
        RECT 1075.8200 1378.2000 1077.4200 1378.6800 ;
        RECT 1075.8200 1372.7600 1077.4200 1373.2400 ;
        RECT 1075.8200 1367.3200 1077.4200 1367.8000 ;
        RECT 1075.8200 1361.8800 1077.4200 1362.3600 ;
        RECT 1075.8200 1356.4400 1077.4200 1356.9200 ;
        RECT 1075.8200 1351.0000 1077.4200 1351.4800 ;
        RECT 1075.8200 1345.5600 1077.4200 1346.0400 ;
        RECT 1075.8200 1340.1200 1077.4200 1340.6000 ;
        RECT 1075.8200 1334.6800 1077.4200 1335.1600 ;
        RECT 1075.8200 1329.2400 1077.4200 1329.7200 ;
        RECT 1273.3200 1323.8000 1274.9200 1324.2800 ;
        RECT 1273.3200 1318.3600 1274.9200 1318.8400 ;
        RECT 1273.3200 1312.9200 1274.9200 1313.4000 ;
        RECT 1273.3200 1307.4800 1274.9200 1307.9600 ;
        RECT 1273.3200 1302.0400 1274.9200 1302.5200 ;
        RECT 1273.3200 1296.6000 1274.9200 1297.0800 ;
        RECT 1273.3200 1291.1600 1274.9200 1291.6400 ;
        RECT 1273.3200 1285.7200 1274.9200 1286.2000 ;
        RECT 1273.3200 1280.2800 1274.9200 1280.7600 ;
        RECT 1273.3200 1274.8400 1274.9200 1275.3200 ;
        RECT 1273.3200 1269.4000 1274.9200 1269.8800 ;
        RECT 1273.3200 1263.9600 1274.9200 1264.4400 ;
        RECT 1273.3200 1258.5200 1274.9200 1259.0000 ;
        RECT 1273.3200 1253.0800 1274.9200 1253.5600 ;
        RECT 1273.3200 1247.6400 1274.9200 1248.1200 ;
        RECT 1273.3200 1236.7600 1274.9200 1237.2400 ;
        RECT 1273.3200 1231.3200 1274.9200 1231.8000 ;
        RECT 1273.3200 1225.8800 1274.9200 1226.3600 ;
        RECT 1273.3200 1220.4400 1274.9200 1220.9200 ;
        RECT 1273.3200 1215.0000 1274.9200 1215.4800 ;
        RECT 1273.3200 1242.2000 1274.9200 1242.6800 ;
        RECT 1273.3200 1209.5600 1274.9200 1210.0400 ;
        RECT 1273.3200 1204.1200 1274.9200 1204.6000 ;
        RECT 1273.3200 1198.6800 1274.9200 1199.1600 ;
        RECT 1273.3200 1193.2400 1274.9200 1193.7200 ;
        RECT 1273.3200 1187.8000 1274.9200 1188.2800 ;
        RECT 1273.3200 1182.3600 1274.9200 1182.8400 ;
        RECT 1273.3200 1176.9200 1274.9200 1177.4000 ;
        RECT 1273.3200 1171.4800 1274.9200 1171.9600 ;
        RECT 1273.3200 1166.0400 1274.9200 1166.5200 ;
        RECT 1273.3200 1160.6000 1274.9200 1161.0800 ;
        RECT 1273.3200 1155.1600 1274.9200 1155.6400 ;
        RECT 1273.3200 1149.7200 1274.9200 1150.2000 ;
        RECT 1273.3200 1144.2800 1274.9200 1144.7600 ;
        RECT 1273.3200 1138.8400 1274.9200 1139.3200 ;
        RECT 1273.3200 1133.4000 1274.9200 1133.8800 ;
        RECT 1273.3200 1127.9600 1274.9200 1128.4400 ;
        RECT 1273.3200 1122.5200 1274.9200 1123.0000 ;
        RECT 1273.3200 1117.0800 1274.9200 1117.5600 ;
        RECT 1273.3200 1111.6400 1274.9200 1112.1200 ;
        RECT 1075.8200 1323.8000 1077.4200 1324.2800 ;
        RECT 1075.8200 1318.3600 1077.4200 1318.8400 ;
        RECT 1075.8200 1312.9200 1077.4200 1313.4000 ;
        RECT 1075.8200 1307.4800 1077.4200 1307.9600 ;
        RECT 1075.8200 1302.0400 1077.4200 1302.5200 ;
        RECT 1075.8200 1296.6000 1077.4200 1297.0800 ;
        RECT 1075.8200 1291.1600 1077.4200 1291.6400 ;
        RECT 1075.8200 1285.7200 1077.4200 1286.2000 ;
        RECT 1075.8200 1280.2800 1077.4200 1280.7600 ;
        RECT 1075.8200 1274.8400 1077.4200 1275.3200 ;
        RECT 1075.8200 1269.4000 1077.4200 1269.8800 ;
        RECT 1075.8200 1263.9600 1077.4200 1264.4400 ;
        RECT 1075.8200 1258.5200 1077.4200 1259.0000 ;
        RECT 1075.8200 1253.0800 1077.4200 1253.5600 ;
        RECT 1075.8200 1247.6400 1077.4200 1248.1200 ;
        RECT 1075.8200 1236.7600 1077.4200 1237.2400 ;
        RECT 1075.8200 1231.3200 1077.4200 1231.8000 ;
        RECT 1075.8200 1225.8800 1077.4200 1226.3600 ;
        RECT 1075.8200 1220.4400 1077.4200 1220.9200 ;
        RECT 1075.8200 1215.0000 1077.4200 1215.4800 ;
        RECT 1075.8200 1242.2000 1077.4200 1242.6800 ;
        RECT 1075.8200 1209.5600 1077.4200 1210.0400 ;
        RECT 1075.8200 1204.1200 1077.4200 1204.6000 ;
        RECT 1075.8200 1198.6800 1077.4200 1199.1600 ;
        RECT 1075.8200 1193.2400 1077.4200 1193.7200 ;
        RECT 1075.8200 1187.8000 1077.4200 1188.2800 ;
        RECT 1075.8200 1182.3600 1077.4200 1182.8400 ;
        RECT 1075.8200 1176.9200 1077.4200 1177.4000 ;
        RECT 1075.8200 1171.4800 1077.4200 1171.9600 ;
        RECT 1075.8200 1166.0400 1077.4200 1166.5200 ;
        RECT 1075.8200 1160.6000 1077.4200 1161.0800 ;
        RECT 1075.8200 1155.1600 1077.4200 1155.6400 ;
        RECT 1075.8200 1149.7200 1077.4200 1150.2000 ;
        RECT 1075.8200 1144.2800 1077.4200 1144.7600 ;
        RECT 1075.8200 1138.8400 1077.4200 1139.3200 ;
        RECT 1075.8200 1133.4000 1077.4200 1133.8800 ;
        RECT 1075.8200 1127.9600 1077.4200 1128.4400 ;
        RECT 1075.8200 1122.5200 1077.4200 1123.0000 ;
        RECT 1075.8200 1117.0800 1077.4200 1117.5600 ;
        RECT 1075.8200 1111.6400 1077.4200 1112.1200 ;
        RECT 1070.2600 1544.6400 1280.4800 1546.2400 ;
        RECT 1070.2600 1107.4500 1280.4800 1109.0500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 1102.0200 1077.4200 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 1550.2400 1077.4200 1551.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 1102.0200 1274.9200 1103.6200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 1550.2400 1274.9200 1551.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1107.4500 1071.8600 1109.0500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1107.4500 1280.4800 1109.0500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1544.6400 1071.8600 1546.2400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1544.6400 1280.4800 1546.2400 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1075.8200 642.7400 1077.4200 1092.5600 ;
        RECT 1273.3200 642.7400 1274.9200 1092.5600 ;
        RECT 1083.5800 648.1700 1085.1800 1086.9600 ;
        RECT 1128.5800 648.1700 1130.1800 1086.9600 ;
        RECT 1173.5800 648.1700 1175.1800 1086.9600 ;
        RECT 1218.5800 648.1700 1220.1800 1086.9600 ;
        RECT 1263.5800 648.1700 1265.1800 1086.9600 ;
      LAYER met3 ;
        RECT 1273.3200 1082.1200 1274.9200 1082.6000 ;
        RECT 1273.3200 1076.6800 1274.9200 1077.1600 ;
        RECT 1273.3200 1071.2400 1274.9200 1071.7200 ;
        RECT 1273.3200 1065.8000 1274.9200 1066.2800 ;
        RECT 1273.3200 1060.3600 1274.9200 1060.8400 ;
        RECT 1273.3200 1054.9200 1274.9200 1055.4000 ;
        RECT 1273.3200 1049.4800 1274.9200 1049.9600 ;
        RECT 1273.3200 1044.0400 1274.9200 1044.5200 ;
        RECT 1273.3200 1038.6000 1274.9200 1039.0800 ;
        RECT 1273.3200 1033.1600 1274.9200 1033.6400 ;
        RECT 1273.3200 1027.7200 1274.9200 1028.2000 ;
        RECT 1273.3200 1022.2800 1274.9200 1022.7600 ;
        RECT 1273.3200 1016.8400 1274.9200 1017.3200 ;
        RECT 1273.3200 1011.4000 1274.9200 1011.8800 ;
        RECT 1273.3200 1005.9600 1274.9200 1006.4400 ;
        RECT 1273.3200 1000.5200 1274.9200 1001.0000 ;
        RECT 1273.3200 995.0800 1274.9200 995.5600 ;
        RECT 1273.3200 989.6400 1274.9200 990.1200 ;
        RECT 1273.3200 984.2000 1274.9200 984.6800 ;
        RECT 1273.3200 978.7600 1274.9200 979.2400 ;
        RECT 1273.3200 973.3200 1274.9200 973.8000 ;
        RECT 1273.3200 967.8800 1274.9200 968.3600 ;
        RECT 1273.3200 962.4400 1274.9200 962.9200 ;
        RECT 1273.3200 957.0000 1274.9200 957.4800 ;
        RECT 1273.3200 946.1200 1274.9200 946.6000 ;
        RECT 1273.3200 940.6800 1274.9200 941.1600 ;
        RECT 1273.3200 935.2400 1274.9200 935.7200 ;
        RECT 1273.3200 929.8000 1274.9200 930.2800 ;
        RECT 1273.3200 924.3600 1274.9200 924.8400 ;
        RECT 1273.3200 951.5600 1274.9200 952.0400 ;
        RECT 1273.3200 918.9200 1274.9200 919.4000 ;
        RECT 1273.3200 913.4800 1274.9200 913.9600 ;
        RECT 1273.3200 908.0400 1274.9200 908.5200 ;
        RECT 1273.3200 902.6000 1274.9200 903.0800 ;
        RECT 1273.3200 897.1600 1274.9200 897.6400 ;
        RECT 1273.3200 891.7200 1274.9200 892.2000 ;
        RECT 1273.3200 886.2800 1274.9200 886.7600 ;
        RECT 1273.3200 880.8400 1274.9200 881.3200 ;
        RECT 1273.3200 875.4000 1274.9200 875.8800 ;
        RECT 1273.3200 869.9600 1274.9200 870.4400 ;
        RECT 1075.8200 1082.1200 1077.4200 1082.6000 ;
        RECT 1075.8200 1076.6800 1077.4200 1077.1600 ;
        RECT 1075.8200 1071.2400 1077.4200 1071.7200 ;
        RECT 1075.8200 1065.8000 1077.4200 1066.2800 ;
        RECT 1075.8200 1060.3600 1077.4200 1060.8400 ;
        RECT 1075.8200 1054.9200 1077.4200 1055.4000 ;
        RECT 1075.8200 1049.4800 1077.4200 1049.9600 ;
        RECT 1075.8200 1044.0400 1077.4200 1044.5200 ;
        RECT 1075.8200 1038.6000 1077.4200 1039.0800 ;
        RECT 1075.8200 1033.1600 1077.4200 1033.6400 ;
        RECT 1075.8200 1027.7200 1077.4200 1028.2000 ;
        RECT 1075.8200 1022.2800 1077.4200 1022.7600 ;
        RECT 1075.8200 1016.8400 1077.4200 1017.3200 ;
        RECT 1075.8200 1011.4000 1077.4200 1011.8800 ;
        RECT 1075.8200 1005.9600 1077.4200 1006.4400 ;
        RECT 1075.8200 1000.5200 1077.4200 1001.0000 ;
        RECT 1075.8200 995.0800 1077.4200 995.5600 ;
        RECT 1075.8200 989.6400 1077.4200 990.1200 ;
        RECT 1075.8200 984.2000 1077.4200 984.6800 ;
        RECT 1075.8200 978.7600 1077.4200 979.2400 ;
        RECT 1075.8200 973.3200 1077.4200 973.8000 ;
        RECT 1075.8200 967.8800 1077.4200 968.3600 ;
        RECT 1075.8200 962.4400 1077.4200 962.9200 ;
        RECT 1075.8200 957.0000 1077.4200 957.4800 ;
        RECT 1075.8200 946.1200 1077.4200 946.6000 ;
        RECT 1075.8200 940.6800 1077.4200 941.1600 ;
        RECT 1075.8200 935.2400 1077.4200 935.7200 ;
        RECT 1075.8200 929.8000 1077.4200 930.2800 ;
        RECT 1075.8200 924.3600 1077.4200 924.8400 ;
        RECT 1075.8200 951.5600 1077.4200 952.0400 ;
        RECT 1075.8200 918.9200 1077.4200 919.4000 ;
        RECT 1075.8200 913.4800 1077.4200 913.9600 ;
        RECT 1075.8200 908.0400 1077.4200 908.5200 ;
        RECT 1075.8200 902.6000 1077.4200 903.0800 ;
        RECT 1075.8200 897.1600 1077.4200 897.6400 ;
        RECT 1075.8200 891.7200 1077.4200 892.2000 ;
        RECT 1075.8200 886.2800 1077.4200 886.7600 ;
        RECT 1075.8200 880.8400 1077.4200 881.3200 ;
        RECT 1075.8200 875.4000 1077.4200 875.8800 ;
        RECT 1075.8200 869.9600 1077.4200 870.4400 ;
        RECT 1273.3200 864.5200 1274.9200 865.0000 ;
        RECT 1273.3200 859.0800 1274.9200 859.5600 ;
        RECT 1273.3200 853.6400 1274.9200 854.1200 ;
        RECT 1273.3200 848.2000 1274.9200 848.6800 ;
        RECT 1273.3200 842.7600 1274.9200 843.2400 ;
        RECT 1273.3200 837.3200 1274.9200 837.8000 ;
        RECT 1273.3200 831.8800 1274.9200 832.3600 ;
        RECT 1273.3200 826.4400 1274.9200 826.9200 ;
        RECT 1273.3200 821.0000 1274.9200 821.4800 ;
        RECT 1273.3200 815.5600 1274.9200 816.0400 ;
        RECT 1273.3200 810.1200 1274.9200 810.6000 ;
        RECT 1273.3200 804.6800 1274.9200 805.1600 ;
        RECT 1273.3200 799.2400 1274.9200 799.7200 ;
        RECT 1273.3200 793.8000 1274.9200 794.2800 ;
        RECT 1273.3200 788.3600 1274.9200 788.8400 ;
        RECT 1273.3200 777.4800 1274.9200 777.9600 ;
        RECT 1273.3200 772.0400 1274.9200 772.5200 ;
        RECT 1273.3200 766.6000 1274.9200 767.0800 ;
        RECT 1273.3200 761.1600 1274.9200 761.6400 ;
        RECT 1273.3200 755.7200 1274.9200 756.2000 ;
        RECT 1273.3200 782.9200 1274.9200 783.4000 ;
        RECT 1273.3200 750.2800 1274.9200 750.7600 ;
        RECT 1273.3200 744.8400 1274.9200 745.3200 ;
        RECT 1273.3200 739.4000 1274.9200 739.8800 ;
        RECT 1273.3200 733.9600 1274.9200 734.4400 ;
        RECT 1273.3200 728.5200 1274.9200 729.0000 ;
        RECT 1273.3200 723.0800 1274.9200 723.5600 ;
        RECT 1273.3200 717.6400 1274.9200 718.1200 ;
        RECT 1273.3200 712.2000 1274.9200 712.6800 ;
        RECT 1273.3200 706.7600 1274.9200 707.2400 ;
        RECT 1273.3200 701.3200 1274.9200 701.8000 ;
        RECT 1273.3200 695.8800 1274.9200 696.3600 ;
        RECT 1273.3200 690.4400 1274.9200 690.9200 ;
        RECT 1273.3200 685.0000 1274.9200 685.4800 ;
        RECT 1273.3200 679.5600 1274.9200 680.0400 ;
        RECT 1273.3200 674.1200 1274.9200 674.6000 ;
        RECT 1273.3200 668.6800 1274.9200 669.1600 ;
        RECT 1273.3200 663.2400 1274.9200 663.7200 ;
        RECT 1273.3200 657.8000 1274.9200 658.2800 ;
        RECT 1273.3200 652.3600 1274.9200 652.8400 ;
        RECT 1075.8200 864.5200 1077.4200 865.0000 ;
        RECT 1075.8200 859.0800 1077.4200 859.5600 ;
        RECT 1075.8200 853.6400 1077.4200 854.1200 ;
        RECT 1075.8200 848.2000 1077.4200 848.6800 ;
        RECT 1075.8200 842.7600 1077.4200 843.2400 ;
        RECT 1075.8200 837.3200 1077.4200 837.8000 ;
        RECT 1075.8200 831.8800 1077.4200 832.3600 ;
        RECT 1075.8200 826.4400 1077.4200 826.9200 ;
        RECT 1075.8200 821.0000 1077.4200 821.4800 ;
        RECT 1075.8200 815.5600 1077.4200 816.0400 ;
        RECT 1075.8200 810.1200 1077.4200 810.6000 ;
        RECT 1075.8200 804.6800 1077.4200 805.1600 ;
        RECT 1075.8200 799.2400 1077.4200 799.7200 ;
        RECT 1075.8200 793.8000 1077.4200 794.2800 ;
        RECT 1075.8200 788.3600 1077.4200 788.8400 ;
        RECT 1075.8200 777.4800 1077.4200 777.9600 ;
        RECT 1075.8200 772.0400 1077.4200 772.5200 ;
        RECT 1075.8200 766.6000 1077.4200 767.0800 ;
        RECT 1075.8200 761.1600 1077.4200 761.6400 ;
        RECT 1075.8200 755.7200 1077.4200 756.2000 ;
        RECT 1075.8200 782.9200 1077.4200 783.4000 ;
        RECT 1075.8200 750.2800 1077.4200 750.7600 ;
        RECT 1075.8200 744.8400 1077.4200 745.3200 ;
        RECT 1075.8200 739.4000 1077.4200 739.8800 ;
        RECT 1075.8200 733.9600 1077.4200 734.4400 ;
        RECT 1075.8200 728.5200 1077.4200 729.0000 ;
        RECT 1075.8200 723.0800 1077.4200 723.5600 ;
        RECT 1075.8200 717.6400 1077.4200 718.1200 ;
        RECT 1075.8200 712.2000 1077.4200 712.6800 ;
        RECT 1075.8200 706.7600 1077.4200 707.2400 ;
        RECT 1075.8200 701.3200 1077.4200 701.8000 ;
        RECT 1075.8200 695.8800 1077.4200 696.3600 ;
        RECT 1075.8200 690.4400 1077.4200 690.9200 ;
        RECT 1075.8200 685.0000 1077.4200 685.4800 ;
        RECT 1075.8200 679.5600 1077.4200 680.0400 ;
        RECT 1075.8200 674.1200 1077.4200 674.6000 ;
        RECT 1075.8200 668.6800 1077.4200 669.1600 ;
        RECT 1075.8200 663.2400 1077.4200 663.7200 ;
        RECT 1075.8200 657.8000 1077.4200 658.2800 ;
        RECT 1075.8200 652.3600 1077.4200 652.8400 ;
        RECT 1070.2600 1085.3600 1280.4800 1086.9600 ;
        RECT 1070.2600 648.1700 1280.4800 649.7700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 642.7400 1077.4200 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 1090.9600 1077.4200 1092.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 642.7400 1274.9200 644.3400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 1090.9600 1274.9200 1092.5600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 648.1700 1071.8600 649.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 648.1700 1280.4800 649.7700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 1085.3600 1071.8600 1086.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 1085.3600 1280.4800 1086.9600 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1075.8200 183.4600 1077.4200 633.2800 ;
        RECT 1273.3200 183.4600 1274.9200 633.2800 ;
        RECT 1083.5800 188.8900 1085.1800 627.6800 ;
        RECT 1128.5800 188.8900 1130.1800 627.6800 ;
        RECT 1173.5800 188.8900 1175.1800 627.6800 ;
        RECT 1218.5800 188.8900 1220.1800 627.6800 ;
        RECT 1263.5800 188.8900 1265.1800 627.6800 ;
      LAYER met3 ;
        RECT 1273.3200 622.8400 1274.9200 623.3200 ;
        RECT 1273.3200 617.4000 1274.9200 617.8800 ;
        RECT 1273.3200 611.9600 1274.9200 612.4400 ;
        RECT 1273.3200 606.5200 1274.9200 607.0000 ;
        RECT 1273.3200 601.0800 1274.9200 601.5600 ;
        RECT 1273.3200 595.6400 1274.9200 596.1200 ;
        RECT 1273.3200 590.2000 1274.9200 590.6800 ;
        RECT 1273.3200 584.7600 1274.9200 585.2400 ;
        RECT 1273.3200 579.3200 1274.9200 579.8000 ;
        RECT 1273.3200 573.8800 1274.9200 574.3600 ;
        RECT 1273.3200 568.4400 1274.9200 568.9200 ;
        RECT 1273.3200 563.0000 1274.9200 563.4800 ;
        RECT 1273.3200 557.5600 1274.9200 558.0400 ;
        RECT 1273.3200 552.1200 1274.9200 552.6000 ;
        RECT 1273.3200 546.6800 1274.9200 547.1600 ;
        RECT 1273.3200 541.2400 1274.9200 541.7200 ;
        RECT 1273.3200 535.8000 1274.9200 536.2800 ;
        RECT 1273.3200 530.3600 1274.9200 530.8400 ;
        RECT 1273.3200 524.9200 1274.9200 525.4000 ;
        RECT 1273.3200 519.4800 1274.9200 519.9600 ;
        RECT 1273.3200 514.0400 1274.9200 514.5200 ;
        RECT 1273.3200 508.6000 1274.9200 509.0800 ;
        RECT 1273.3200 503.1600 1274.9200 503.6400 ;
        RECT 1273.3200 497.7200 1274.9200 498.2000 ;
        RECT 1273.3200 486.8400 1274.9200 487.3200 ;
        RECT 1273.3200 481.4000 1274.9200 481.8800 ;
        RECT 1273.3200 475.9600 1274.9200 476.4400 ;
        RECT 1273.3200 470.5200 1274.9200 471.0000 ;
        RECT 1273.3200 465.0800 1274.9200 465.5600 ;
        RECT 1273.3200 492.2800 1274.9200 492.7600 ;
        RECT 1273.3200 459.6400 1274.9200 460.1200 ;
        RECT 1273.3200 454.2000 1274.9200 454.6800 ;
        RECT 1273.3200 448.7600 1274.9200 449.2400 ;
        RECT 1273.3200 443.3200 1274.9200 443.8000 ;
        RECT 1273.3200 437.8800 1274.9200 438.3600 ;
        RECT 1273.3200 432.4400 1274.9200 432.9200 ;
        RECT 1273.3200 427.0000 1274.9200 427.4800 ;
        RECT 1273.3200 421.5600 1274.9200 422.0400 ;
        RECT 1273.3200 416.1200 1274.9200 416.6000 ;
        RECT 1273.3200 410.6800 1274.9200 411.1600 ;
        RECT 1075.8200 622.8400 1077.4200 623.3200 ;
        RECT 1075.8200 617.4000 1077.4200 617.8800 ;
        RECT 1075.8200 611.9600 1077.4200 612.4400 ;
        RECT 1075.8200 606.5200 1077.4200 607.0000 ;
        RECT 1075.8200 601.0800 1077.4200 601.5600 ;
        RECT 1075.8200 595.6400 1077.4200 596.1200 ;
        RECT 1075.8200 590.2000 1077.4200 590.6800 ;
        RECT 1075.8200 584.7600 1077.4200 585.2400 ;
        RECT 1075.8200 579.3200 1077.4200 579.8000 ;
        RECT 1075.8200 573.8800 1077.4200 574.3600 ;
        RECT 1075.8200 568.4400 1077.4200 568.9200 ;
        RECT 1075.8200 563.0000 1077.4200 563.4800 ;
        RECT 1075.8200 557.5600 1077.4200 558.0400 ;
        RECT 1075.8200 552.1200 1077.4200 552.6000 ;
        RECT 1075.8200 546.6800 1077.4200 547.1600 ;
        RECT 1075.8200 541.2400 1077.4200 541.7200 ;
        RECT 1075.8200 535.8000 1077.4200 536.2800 ;
        RECT 1075.8200 530.3600 1077.4200 530.8400 ;
        RECT 1075.8200 524.9200 1077.4200 525.4000 ;
        RECT 1075.8200 519.4800 1077.4200 519.9600 ;
        RECT 1075.8200 514.0400 1077.4200 514.5200 ;
        RECT 1075.8200 508.6000 1077.4200 509.0800 ;
        RECT 1075.8200 503.1600 1077.4200 503.6400 ;
        RECT 1075.8200 497.7200 1077.4200 498.2000 ;
        RECT 1075.8200 486.8400 1077.4200 487.3200 ;
        RECT 1075.8200 481.4000 1077.4200 481.8800 ;
        RECT 1075.8200 475.9600 1077.4200 476.4400 ;
        RECT 1075.8200 470.5200 1077.4200 471.0000 ;
        RECT 1075.8200 465.0800 1077.4200 465.5600 ;
        RECT 1075.8200 492.2800 1077.4200 492.7600 ;
        RECT 1075.8200 459.6400 1077.4200 460.1200 ;
        RECT 1075.8200 454.2000 1077.4200 454.6800 ;
        RECT 1075.8200 448.7600 1077.4200 449.2400 ;
        RECT 1075.8200 443.3200 1077.4200 443.8000 ;
        RECT 1075.8200 437.8800 1077.4200 438.3600 ;
        RECT 1075.8200 432.4400 1077.4200 432.9200 ;
        RECT 1075.8200 427.0000 1077.4200 427.4800 ;
        RECT 1075.8200 421.5600 1077.4200 422.0400 ;
        RECT 1075.8200 416.1200 1077.4200 416.6000 ;
        RECT 1075.8200 410.6800 1077.4200 411.1600 ;
        RECT 1273.3200 405.2400 1274.9200 405.7200 ;
        RECT 1273.3200 399.8000 1274.9200 400.2800 ;
        RECT 1273.3200 394.3600 1274.9200 394.8400 ;
        RECT 1273.3200 388.9200 1274.9200 389.4000 ;
        RECT 1273.3200 383.4800 1274.9200 383.9600 ;
        RECT 1273.3200 378.0400 1274.9200 378.5200 ;
        RECT 1273.3200 372.6000 1274.9200 373.0800 ;
        RECT 1273.3200 367.1600 1274.9200 367.6400 ;
        RECT 1273.3200 361.7200 1274.9200 362.2000 ;
        RECT 1273.3200 356.2800 1274.9200 356.7600 ;
        RECT 1273.3200 350.8400 1274.9200 351.3200 ;
        RECT 1273.3200 345.4000 1274.9200 345.8800 ;
        RECT 1273.3200 339.9600 1274.9200 340.4400 ;
        RECT 1273.3200 334.5200 1274.9200 335.0000 ;
        RECT 1273.3200 329.0800 1274.9200 329.5600 ;
        RECT 1273.3200 318.2000 1274.9200 318.6800 ;
        RECT 1273.3200 312.7600 1274.9200 313.2400 ;
        RECT 1273.3200 307.3200 1274.9200 307.8000 ;
        RECT 1273.3200 301.8800 1274.9200 302.3600 ;
        RECT 1273.3200 296.4400 1274.9200 296.9200 ;
        RECT 1273.3200 323.6400 1274.9200 324.1200 ;
        RECT 1273.3200 291.0000 1274.9200 291.4800 ;
        RECT 1273.3200 285.5600 1274.9200 286.0400 ;
        RECT 1273.3200 280.1200 1274.9200 280.6000 ;
        RECT 1273.3200 274.6800 1274.9200 275.1600 ;
        RECT 1273.3200 269.2400 1274.9200 269.7200 ;
        RECT 1273.3200 263.8000 1274.9200 264.2800 ;
        RECT 1273.3200 258.3600 1274.9200 258.8400 ;
        RECT 1273.3200 252.9200 1274.9200 253.4000 ;
        RECT 1273.3200 247.4800 1274.9200 247.9600 ;
        RECT 1273.3200 242.0400 1274.9200 242.5200 ;
        RECT 1273.3200 236.6000 1274.9200 237.0800 ;
        RECT 1273.3200 231.1600 1274.9200 231.6400 ;
        RECT 1273.3200 225.7200 1274.9200 226.2000 ;
        RECT 1273.3200 220.2800 1274.9200 220.7600 ;
        RECT 1273.3200 214.8400 1274.9200 215.3200 ;
        RECT 1273.3200 209.4000 1274.9200 209.8800 ;
        RECT 1273.3200 203.9600 1274.9200 204.4400 ;
        RECT 1273.3200 198.5200 1274.9200 199.0000 ;
        RECT 1273.3200 193.0800 1274.9200 193.5600 ;
        RECT 1075.8200 405.2400 1077.4200 405.7200 ;
        RECT 1075.8200 399.8000 1077.4200 400.2800 ;
        RECT 1075.8200 394.3600 1077.4200 394.8400 ;
        RECT 1075.8200 388.9200 1077.4200 389.4000 ;
        RECT 1075.8200 383.4800 1077.4200 383.9600 ;
        RECT 1075.8200 378.0400 1077.4200 378.5200 ;
        RECT 1075.8200 372.6000 1077.4200 373.0800 ;
        RECT 1075.8200 367.1600 1077.4200 367.6400 ;
        RECT 1075.8200 361.7200 1077.4200 362.2000 ;
        RECT 1075.8200 356.2800 1077.4200 356.7600 ;
        RECT 1075.8200 350.8400 1077.4200 351.3200 ;
        RECT 1075.8200 345.4000 1077.4200 345.8800 ;
        RECT 1075.8200 339.9600 1077.4200 340.4400 ;
        RECT 1075.8200 334.5200 1077.4200 335.0000 ;
        RECT 1075.8200 329.0800 1077.4200 329.5600 ;
        RECT 1075.8200 318.2000 1077.4200 318.6800 ;
        RECT 1075.8200 312.7600 1077.4200 313.2400 ;
        RECT 1075.8200 307.3200 1077.4200 307.8000 ;
        RECT 1075.8200 301.8800 1077.4200 302.3600 ;
        RECT 1075.8200 296.4400 1077.4200 296.9200 ;
        RECT 1075.8200 323.6400 1077.4200 324.1200 ;
        RECT 1075.8200 291.0000 1077.4200 291.4800 ;
        RECT 1075.8200 285.5600 1077.4200 286.0400 ;
        RECT 1075.8200 280.1200 1077.4200 280.6000 ;
        RECT 1075.8200 274.6800 1077.4200 275.1600 ;
        RECT 1075.8200 269.2400 1077.4200 269.7200 ;
        RECT 1075.8200 263.8000 1077.4200 264.2800 ;
        RECT 1075.8200 258.3600 1077.4200 258.8400 ;
        RECT 1075.8200 252.9200 1077.4200 253.4000 ;
        RECT 1075.8200 247.4800 1077.4200 247.9600 ;
        RECT 1075.8200 242.0400 1077.4200 242.5200 ;
        RECT 1075.8200 236.6000 1077.4200 237.0800 ;
        RECT 1075.8200 231.1600 1077.4200 231.6400 ;
        RECT 1075.8200 225.7200 1077.4200 226.2000 ;
        RECT 1075.8200 220.2800 1077.4200 220.7600 ;
        RECT 1075.8200 214.8400 1077.4200 215.3200 ;
        RECT 1075.8200 209.4000 1077.4200 209.8800 ;
        RECT 1075.8200 203.9600 1077.4200 204.4400 ;
        RECT 1075.8200 198.5200 1077.4200 199.0000 ;
        RECT 1075.8200 193.0800 1077.4200 193.5600 ;
        RECT 1070.2600 626.0800 1280.4800 627.6800 ;
        RECT 1070.2600 188.8900 1280.4800 190.4900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 183.4600 1077.4200 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.8200 631.6800 1077.4200 633.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 183.4600 1274.9200 185.0600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1273.3200 631.6800 1274.9200 633.2800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 188.8900 1071.8600 190.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 188.8900 1280.4800 190.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1070.2600 626.0800 1071.8600 627.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1278.8800 626.0800 1280.4800 627.6800 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1295.8000 2479.6000 1297.4000 2509.8600 ;
        RECT 1493.5000 2479.6000 1495.1000 2509.8600 ;
      LAYER met3 ;
        RECT 1493.5000 2497.3800 1495.1000 2497.8600 ;
        RECT 1295.8000 2497.3800 1297.4000 2497.8600 ;
        RECT 1493.5000 2491.9400 1495.1000 2492.4200 ;
        RECT 1493.5000 2486.5000 1495.1000 2486.9800 ;
        RECT 1295.8000 2491.9400 1297.4000 2492.4200 ;
        RECT 1295.8000 2486.5000 1297.4000 2486.9800 ;
        RECT 1290.3400 2503.1000 1500.5600 2504.7000 ;
        RECT 1290.3400 2483.5700 1500.5600 2485.1700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.8000 2479.6000 1297.4000 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.8000 2508.2600 1297.4000 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.5000 2479.6000 1495.1000 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.5000 2508.2600 1495.1000 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2483.5700 1291.9400 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2483.5700 1500.5600 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2503.1000 1291.9400 2504.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2503.1000 1500.5600 2504.7000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 188.6300 1485.2600 396.7300 ;
        RECT 1438.6600 188.6300 1440.2600 396.7300 ;
        RECT 1393.6600 188.6300 1395.2600 396.7300 ;
        RECT 1348.6600 188.6300 1350.2600 396.7300 ;
        RECT 1303.6600 188.6300 1305.2600 396.7300 ;
        RECT 1493.4000 183.2000 1495.0000 402.8400 ;
        RECT 1295.9000 183.2000 1297.5000 402.8400 ;
      LAYER met3 ;
        RECT 1493.4000 377.7800 1495.0000 378.2600 ;
        RECT 1493.4000 383.2200 1495.0000 383.7000 ;
        RECT 1483.6600 377.7800 1485.2600 378.2600 ;
        RECT 1483.6600 383.2200 1485.2600 383.7000 ;
        RECT 1483.6600 388.6600 1485.2600 389.1400 ;
        RECT 1493.4000 388.6600 1495.0000 389.1400 ;
        RECT 1493.4000 366.9000 1495.0000 367.3800 ;
        RECT 1493.4000 372.3400 1495.0000 372.8200 ;
        RECT 1483.6600 366.9000 1485.2600 367.3800 ;
        RECT 1483.6600 372.3400 1485.2600 372.8200 ;
        RECT 1493.4000 350.5800 1495.0000 351.0600 ;
        RECT 1493.4000 356.0200 1495.0000 356.5000 ;
        RECT 1483.6600 350.5800 1485.2600 351.0600 ;
        RECT 1483.6600 356.0200 1485.2600 356.5000 ;
        RECT 1483.6600 361.4600 1485.2600 361.9400 ;
        RECT 1493.4000 361.4600 1495.0000 361.9400 ;
        RECT 1438.6600 377.7800 1440.2600 378.2600 ;
        RECT 1438.6600 383.2200 1440.2600 383.7000 ;
        RECT 1438.6600 388.6600 1440.2600 389.1400 ;
        RECT 1438.6600 366.9000 1440.2600 367.3800 ;
        RECT 1438.6600 372.3400 1440.2600 372.8200 ;
        RECT 1438.6600 350.5800 1440.2600 351.0600 ;
        RECT 1438.6600 356.0200 1440.2600 356.5000 ;
        RECT 1438.6600 361.4600 1440.2600 361.9400 ;
        RECT 1493.4000 334.2600 1495.0000 334.7400 ;
        RECT 1493.4000 339.7000 1495.0000 340.1800 ;
        RECT 1493.4000 345.1400 1495.0000 345.6200 ;
        RECT 1483.6600 334.2600 1485.2600 334.7400 ;
        RECT 1483.6600 339.7000 1485.2600 340.1800 ;
        RECT 1483.6600 345.1400 1485.2600 345.6200 ;
        RECT 1493.4000 323.3800 1495.0000 323.8600 ;
        RECT 1493.4000 328.8200 1495.0000 329.3000 ;
        RECT 1483.6600 323.3800 1485.2600 323.8600 ;
        RECT 1483.6600 328.8200 1485.2600 329.3000 ;
        RECT 1493.4000 307.0600 1495.0000 307.5400 ;
        RECT 1493.4000 312.5000 1495.0000 312.9800 ;
        RECT 1493.4000 317.9400 1495.0000 318.4200 ;
        RECT 1483.6600 307.0600 1485.2600 307.5400 ;
        RECT 1483.6600 312.5000 1485.2600 312.9800 ;
        RECT 1483.6600 317.9400 1485.2600 318.4200 ;
        RECT 1493.4000 296.1800 1495.0000 296.6600 ;
        RECT 1493.4000 301.6200 1495.0000 302.1000 ;
        RECT 1483.6600 296.1800 1485.2600 296.6600 ;
        RECT 1483.6600 301.6200 1485.2600 302.1000 ;
        RECT 1438.6600 334.2600 1440.2600 334.7400 ;
        RECT 1438.6600 339.7000 1440.2600 340.1800 ;
        RECT 1438.6600 345.1400 1440.2600 345.6200 ;
        RECT 1438.6600 323.3800 1440.2600 323.8600 ;
        RECT 1438.6600 328.8200 1440.2600 329.3000 ;
        RECT 1438.6600 307.0600 1440.2600 307.5400 ;
        RECT 1438.6600 312.5000 1440.2600 312.9800 ;
        RECT 1438.6600 317.9400 1440.2600 318.4200 ;
        RECT 1438.6600 296.1800 1440.2600 296.6600 ;
        RECT 1438.6600 301.6200 1440.2600 302.1000 ;
        RECT 1393.6600 377.7800 1395.2600 378.2600 ;
        RECT 1393.6600 383.2200 1395.2600 383.7000 ;
        RECT 1393.6600 388.6600 1395.2600 389.1400 ;
        RECT 1348.6600 377.7800 1350.2600 378.2600 ;
        RECT 1348.6600 383.2200 1350.2600 383.7000 ;
        RECT 1348.6600 388.6600 1350.2600 389.1400 ;
        RECT 1393.6600 366.9000 1395.2600 367.3800 ;
        RECT 1393.6600 372.3400 1395.2600 372.8200 ;
        RECT 1393.6600 350.5800 1395.2600 351.0600 ;
        RECT 1393.6600 356.0200 1395.2600 356.5000 ;
        RECT 1393.6600 361.4600 1395.2600 361.9400 ;
        RECT 1348.6600 366.9000 1350.2600 367.3800 ;
        RECT 1348.6600 372.3400 1350.2600 372.8200 ;
        RECT 1348.6600 350.5800 1350.2600 351.0600 ;
        RECT 1348.6600 356.0200 1350.2600 356.5000 ;
        RECT 1348.6600 361.4600 1350.2600 361.9400 ;
        RECT 1303.6600 377.7800 1305.2600 378.2600 ;
        RECT 1303.6600 383.2200 1305.2600 383.7000 ;
        RECT 1295.9000 377.7800 1297.5000 378.2600 ;
        RECT 1295.9000 383.2200 1297.5000 383.7000 ;
        RECT 1295.9000 388.6600 1297.5000 389.1400 ;
        RECT 1303.6600 388.6600 1305.2600 389.1400 ;
        RECT 1303.6600 366.9000 1305.2600 367.3800 ;
        RECT 1303.6600 372.3400 1305.2600 372.8200 ;
        RECT 1295.9000 366.9000 1297.5000 367.3800 ;
        RECT 1295.9000 372.3400 1297.5000 372.8200 ;
        RECT 1303.6600 350.5800 1305.2600 351.0600 ;
        RECT 1303.6600 356.0200 1305.2600 356.5000 ;
        RECT 1295.9000 350.5800 1297.5000 351.0600 ;
        RECT 1295.9000 356.0200 1297.5000 356.5000 ;
        RECT 1295.9000 361.4600 1297.5000 361.9400 ;
        RECT 1303.6600 361.4600 1305.2600 361.9400 ;
        RECT 1393.6600 334.2600 1395.2600 334.7400 ;
        RECT 1393.6600 339.7000 1395.2600 340.1800 ;
        RECT 1393.6600 345.1400 1395.2600 345.6200 ;
        RECT 1393.6600 323.3800 1395.2600 323.8600 ;
        RECT 1393.6600 328.8200 1395.2600 329.3000 ;
        RECT 1348.6600 334.2600 1350.2600 334.7400 ;
        RECT 1348.6600 339.7000 1350.2600 340.1800 ;
        RECT 1348.6600 345.1400 1350.2600 345.6200 ;
        RECT 1348.6600 323.3800 1350.2600 323.8600 ;
        RECT 1348.6600 328.8200 1350.2600 329.3000 ;
        RECT 1393.6600 307.0600 1395.2600 307.5400 ;
        RECT 1393.6600 312.5000 1395.2600 312.9800 ;
        RECT 1393.6600 317.9400 1395.2600 318.4200 ;
        RECT 1393.6600 296.1800 1395.2600 296.6600 ;
        RECT 1393.6600 301.6200 1395.2600 302.1000 ;
        RECT 1348.6600 307.0600 1350.2600 307.5400 ;
        RECT 1348.6600 312.5000 1350.2600 312.9800 ;
        RECT 1348.6600 317.9400 1350.2600 318.4200 ;
        RECT 1348.6600 296.1800 1350.2600 296.6600 ;
        RECT 1348.6600 301.6200 1350.2600 302.1000 ;
        RECT 1303.6600 334.2600 1305.2600 334.7400 ;
        RECT 1303.6600 339.7000 1305.2600 340.1800 ;
        RECT 1303.6600 345.1400 1305.2600 345.6200 ;
        RECT 1295.9000 334.2600 1297.5000 334.7400 ;
        RECT 1295.9000 339.7000 1297.5000 340.1800 ;
        RECT 1295.9000 345.1400 1297.5000 345.6200 ;
        RECT 1303.6600 323.3800 1305.2600 323.8600 ;
        RECT 1303.6600 328.8200 1305.2600 329.3000 ;
        RECT 1295.9000 323.3800 1297.5000 323.8600 ;
        RECT 1295.9000 328.8200 1297.5000 329.3000 ;
        RECT 1303.6600 307.0600 1305.2600 307.5400 ;
        RECT 1303.6600 312.5000 1305.2600 312.9800 ;
        RECT 1303.6600 317.9400 1305.2600 318.4200 ;
        RECT 1295.9000 307.0600 1297.5000 307.5400 ;
        RECT 1295.9000 312.5000 1297.5000 312.9800 ;
        RECT 1295.9000 317.9400 1297.5000 318.4200 ;
        RECT 1303.6600 296.1800 1305.2600 296.6600 ;
        RECT 1303.6600 301.6200 1305.2600 302.1000 ;
        RECT 1295.9000 296.1800 1297.5000 296.6600 ;
        RECT 1295.9000 301.6200 1297.5000 302.1000 ;
        RECT 1493.4000 279.8600 1495.0000 280.3400 ;
        RECT 1493.4000 285.3000 1495.0000 285.7800 ;
        RECT 1493.4000 290.7400 1495.0000 291.2200 ;
        RECT 1483.6600 279.8600 1485.2600 280.3400 ;
        RECT 1483.6600 285.3000 1485.2600 285.7800 ;
        RECT 1483.6600 290.7400 1485.2600 291.2200 ;
        RECT 1493.4000 268.9800 1495.0000 269.4600 ;
        RECT 1493.4000 274.4200 1495.0000 274.9000 ;
        RECT 1483.6600 268.9800 1485.2600 269.4600 ;
        RECT 1483.6600 274.4200 1485.2600 274.9000 ;
        RECT 1493.4000 252.6600 1495.0000 253.1400 ;
        RECT 1493.4000 258.1000 1495.0000 258.5800 ;
        RECT 1493.4000 263.5400 1495.0000 264.0200 ;
        RECT 1483.6600 252.6600 1485.2600 253.1400 ;
        RECT 1483.6600 258.1000 1485.2600 258.5800 ;
        RECT 1483.6600 263.5400 1485.2600 264.0200 ;
        RECT 1493.4000 241.7800 1495.0000 242.2600 ;
        RECT 1493.4000 247.2200 1495.0000 247.7000 ;
        RECT 1483.6600 241.7800 1485.2600 242.2600 ;
        RECT 1483.6600 247.2200 1485.2600 247.7000 ;
        RECT 1438.6600 279.8600 1440.2600 280.3400 ;
        RECT 1438.6600 285.3000 1440.2600 285.7800 ;
        RECT 1438.6600 290.7400 1440.2600 291.2200 ;
        RECT 1438.6600 268.9800 1440.2600 269.4600 ;
        RECT 1438.6600 274.4200 1440.2600 274.9000 ;
        RECT 1438.6600 252.6600 1440.2600 253.1400 ;
        RECT 1438.6600 258.1000 1440.2600 258.5800 ;
        RECT 1438.6600 263.5400 1440.2600 264.0200 ;
        RECT 1438.6600 241.7800 1440.2600 242.2600 ;
        RECT 1438.6600 247.2200 1440.2600 247.7000 ;
        RECT 1493.4000 225.4600 1495.0000 225.9400 ;
        RECT 1493.4000 230.9000 1495.0000 231.3800 ;
        RECT 1493.4000 236.3400 1495.0000 236.8200 ;
        RECT 1483.6600 225.4600 1485.2600 225.9400 ;
        RECT 1483.6600 230.9000 1485.2600 231.3800 ;
        RECT 1483.6600 236.3400 1485.2600 236.8200 ;
        RECT 1493.4000 214.5800 1495.0000 215.0600 ;
        RECT 1493.4000 220.0200 1495.0000 220.5000 ;
        RECT 1483.6600 214.5800 1485.2600 215.0600 ;
        RECT 1483.6600 220.0200 1485.2600 220.5000 ;
        RECT 1493.4000 198.2600 1495.0000 198.7400 ;
        RECT 1493.4000 203.7000 1495.0000 204.1800 ;
        RECT 1493.4000 209.1400 1495.0000 209.6200 ;
        RECT 1483.6600 198.2600 1485.2600 198.7400 ;
        RECT 1483.6600 203.7000 1485.2600 204.1800 ;
        RECT 1483.6600 209.1400 1485.2600 209.6200 ;
        RECT 1483.6600 192.8200 1485.2600 193.3000 ;
        RECT 1493.4000 192.8200 1495.0000 193.3000 ;
        RECT 1438.6600 225.4600 1440.2600 225.9400 ;
        RECT 1438.6600 230.9000 1440.2600 231.3800 ;
        RECT 1438.6600 236.3400 1440.2600 236.8200 ;
        RECT 1438.6600 214.5800 1440.2600 215.0600 ;
        RECT 1438.6600 220.0200 1440.2600 220.5000 ;
        RECT 1438.6600 198.2600 1440.2600 198.7400 ;
        RECT 1438.6600 203.7000 1440.2600 204.1800 ;
        RECT 1438.6600 209.1400 1440.2600 209.6200 ;
        RECT 1438.6600 192.8200 1440.2600 193.3000 ;
        RECT 1393.6600 279.8600 1395.2600 280.3400 ;
        RECT 1393.6600 285.3000 1395.2600 285.7800 ;
        RECT 1393.6600 290.7400 1395.2600 291.2200 ;
        RECT 1393.6600 268.9800 1395.2600 269.4600 ;
        RECT 1393.6600 274.4200 1395.2600 274.9000 ;
        RECT 1348.6600 279.8600 1350.2600 280.3400 ;
        RECT 1348.6600 285.3000 1350.2600 285.7800 ;
        RECT 1348.6600 290.7400 1350.2600 291.2200 ;
        RECT 1348.6600 268.9800 1350.2600 269.4600 ;
        RECT 1348.6600 274.4200 1350.2600 274.9000 ;
        RECT 1393.6600 252.6600 1395.2600 253.1400 ;
        RECT 1393.6600 258.1000 1395.2600 258.5800 ;
        RECT 1393.6600 263.5400 1395.2600 264.0200 ;
        RECT 1393.6600 241.7800 1395.2600 242.2600 ;
        RECT 1393.6600 247.2200 1395.2600 247.7000 ;
        RECT 1348.6600 252.6600 1350.2600 253.1400 ;
        RECT 1348.6600 258.1000 1350.2600 258.5800 ;
        RECT 1348.6600 263.5400 1350.2600 264.0200 ;
        RECT 1348.6600 241.7800 1350.2600 242.2600 ;
        RECT 1348.6600 247.2200 1350.2600 247.7000 ;
        RECT 1303.6600 279.8600 1305.2600 280.3400 ;
        RECT 1303.6600 285.3000 1305.2600 285.7800 ;
        RECT 1303.6600 290.7400 1305.2600 291.2200 ;
        RECT 1295.9000 279.8600 1297.5000 280.3400 ;
        RECT 1295.9000 285.3000 1297.5000 285.7800 ;
        RECT 1295.9000 290.7400 1297.5000 291.2200 ;
        RECT 1303.6600 268.9800 1305.2600 269.4600 ;
        RECT 1303.6600 274.4200 1305.2600 274.9000 ;
        RECT 1295.9000 268.9800 1297.5000 269.4600 ;
        RECT 1295.9000 274.4200 1297.5000 274.9000 ;
        RECT 1303.6600 252.6600 1305.2600 253.1400 ;
        RECT 1303.6600 258.1000 1305.2600 258.5800 ;
        RECT 1303.6600 263.5400 1305.2600 264.0200 ;
        RECT 1295.9000 252.6600 1297.5000 253.1400 ;
        RECT 1295.9000 258.1000 1297.5000 258.5800 ;
        RECT 1295.9000 263.5400 1297.5000 264.0200 ;
        RECT 1303.6600 241.7800 1305.2600 242.2600 ;
        RECT 1303.6600 247.2200 1305.2600 247.7000 ;
        RECT 1295.9000 241.7800 1297.5000 242.2600 ;
        RECT 1295.9000 247.2200 1297.5000 247.7000 ;
        RECT 1393.6600 225.4600 1395.2600 225.9400 ;
        RECT 1393.6600 230.9000 1395.2600 231.3800 ;
        RECT 1393.6600 236.3400 1395.2600 236.8200 ;
        RECT 1393.6600 214.5800 1395.2600 215.0600 ;
        RECT 1393.6600 220.0200 1395.2600 220.5000 ;
        RECT 1348.6600 225.4600 1350.2600 225.9400 ;
        RECT 1348.6600 230.9000 1350.2600 231.3800 ;
        RECT 1348.6600 236.3400 1350.2600 236.8200 ;
        RECT 1348.6600 214.5800 1350.2600 215.0600 ;
        RECT 1348.6600 220.0200 1350.2600 220.5000 ;
        RECT 1393.6600 198.2600 1395.2600 198.7400 ;
        RECT 1393.6600 203.7000 1395.2600 204.1800 ;
        RECT 1393.6600 209.1400 1395.2600 209.6200 ;
        RECT 1393.6600 192.8200 1395.2600 193.3000 ;
        RECT 1348.6600 198.2600 1350.2600 198.7400 ;
        RECT 1348.6600 203.7000 1350.2600 204.1800 ;
        RECT 1348.6600 209.1400 1350.2600 209.6200 ;
        RECT 1348.6600 192.8200 1350.2600 193.3000 ;
        RECT 1303.6600 225.4600 1305.2600 225.9400 ;
        RECT 1303.6600 230.9000 1305.2600 231.3800 ;
        RECT 1303.6600 236.3400 1305.2600 236.8200 ;
        RECT 1295.9000 225.4600 1297.5000 225.9400 ;
        RECT 1295.9000 230.9000 1297.5000 231.3800 ;
        RECT 1295.9000 236.3400 1297.5000 236.8200 ;
        RECT 1303.6600 214.5800 1305.2600 215.0600 ;
        RECT 1303.6600 220.0200 1305.2600 220.5000 ;
        RECT 1295.9000 214.5800 1297.5000 215.0600 ;
        RECT 1295.9000 220.0200 1297.5000 220.5000 ;
        RECT 1303.6600 198.2600 1305.2600 198.7400 ;
        RECT 1303.6600 203.7000 1305.2600 204.1800 ;
        RECT 1303.6600 209.1400 1305.2600 209.6200 ;
        RECT 1295.9000 198.2600 1297.5000 198.7400 ;
        RECT 1295.9000 203.7000 1297.5000 204.1800 ;
        RECT 1295.9000 209.1400 1297.5000 209.6200 ;
        RECT 1295.9000 192.8200 1297.5000 193.3000 ;
        RECT 1303.6600 192.8200 1305.2600 193.3000 ;
        RECT 1290.3400 395.1300 1500.5600 396.7300 ;
        RECT 1290.3400 188.6300 1500.5600 190.2300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 183.2000 1297.5000 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 401.2400 1297.5000 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 183.2000 1495.0000 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 401.2400 1495.0000 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 188.6300 1291.9400 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 188.6300 1500.5600 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 395.1300 1291.9400 396.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 395.1300 1500.5600 396.7300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1295.8000 142.9400 1297.4000 173.2000 ;
        RECT 1493.5000 142.9400 1495.1000 173.2000 ;
      LAYER met3 ;
        RECT 1493.5000 160.7200 1495.1000 161.2000 ;
        RECT 1295.8000 160.7200 1297.4000 161.2000 ;
        RECT 1493.5000 155.2800 1495.1000 155.7600 ;
        RECT 1493.5000 149.8400 1495.1000 150.3200 ;
        RECT 1295.8000 155.2800 1297.4000 155.7600 ;
        RECT 1295.8000 149.8400 1297.4000 150.3200 ;
        RECT 1290.3400 166.4400 1500.5600 168.0400 ;
        RECT 1290.3400 146.9100 1500.5600 148.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.8000 142.9400 1297.4000 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.8000 171.6000 1297.4000 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.5000 142.9400 1495.1000 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.5000 171.6000 1495.1000 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 146.9100 1291.9400 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 146.9100 1500.5600 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 166.4400 1291.9400 168.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 166.4400 1500.5600 168.0400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 2255.3900 1485.2600 2463.4900 ;
        RECT 1438.6600 2255.3900 1440.2600 2463.4900 ;
        RECT 1393.6600 2255.3900 1395.2600 2463.4900 ;
        RECT 1348.6600 2255.3900 1350.2600 2463.4900 ;
        RECT 1303.6600 2255.3900 1305.2600 2463.4900 ;
        RECT 1493.4000 2249.9600 1495.0000 2469.6000 ;
        RECT 1295.9000 2249.9600 1297.5000 2469.6000 ;
      LAYER met3 ;
        RECT 1493.4000 2444.5400 1495.0000 2445.0200 ;
        RECT 1493.4000 2449.9800 1495.0000 2450.4600 ;
        RECT 1483.6600 2444.5400 1485.2600 2445.0200 ;
        RECT 1483.6600 2449.9800 1485.2600 2450.4600 ;
        RECT 1483.6600 2455.4200 1485.2600 2455.9000 ;
        RECT 1493.4000 2455.4200 1495.0000 2455.9000 ;
        RECT 1493.4000 2433.6600 1495.0000 2434.1400 ;
        RECT 1493.4000 2439.1000 1495.0000 2439.5800 ;
        RECT 1483.6600 2433.6600 1485.2600 2434.1400 ;
        RECT 1483.6600 2439.1000 1485.2600 2439.5800 ;
        RECT 1493.4000 2417.3400 1495.0000 2417.8200 ;
        RECT 1493.4000 2422.7800 1495.0000 2423.2600 ;
        RECT 1483.6600 2417.3400 1485.2600 2417.8200 ;
        RECT 1483.6600 2422.7800 1485.2600 2423.2600 ;
        RECT 1483.6600 2428.2200 1485.2600 2428.7000 ;
        RECT 1493.4000 2428.2200 1495.0000 2428.7000 ;
        RECT 1438.6600 2444.5400 1440.2600 2445.0200 ;
        RECT 1438.6600 2449.9800 1440.2600 2450.4600 ;
        RECT 1438.6600 2455.4200 1440.2600 2455.9000 ;
        RECT 1438.6600 2433.6600 1440.2600 2434.1400 ;
        RECT 1438.6600 2439.1000 1440.2600 2439.5800 ;
        RECT 1438.6600 2417.3400 1440.2600 2417.8200 ;
        RECT 1438.6600 2422.7800 1440.2600 2423.2600 ;
        RECT 1438.6600 2428.2200 1440.2600 2428.7000 ;
        RECT 1493.4000 2401.0200 1495.0000 2401.5000 ;
        RECT 1493.4000 2406.4600 1495.0000 2406.9400 ;
        RECT 1493.4000 2411.9000 1495.0000 2412.3800 ;
        RECT 1483.6600 2401.0200 1485.2600 2401.5000 ;
        RECT 1483.6600 2406.4600 1485.2600 2406.9400 ;
        RECT 1483.6600 2411.9000 1485.2600 2412.3800 ;
        RECT 1493.4000 2390.1400 1495.0000 2390.6200 ;
        RECT 1493.4000 2395.5800 1495.0000 2396.0600 ;
        RECT 1483.6600 2390.1400 1485.2600 2390.6200 ;
        RECT 1483.6600 2395.5800 1485.2600 2396.0600 ;
        RECT 1493.4000 2373.8200 1495.0000 2374.3000 ;
        RECT 1493.4000 2379.2600 1495.0000 2379.7400 ;
        RECT 1493.4000 2384.7000 1495.0000 2385.1800 ;
        RECT 1483.6600 2373.8200 1485.2600 2374.3000 ;
        RECT 1483.6600 2379.2600 1485.2600 2379.7400 ;
        RECT 1483.6600 2384.7000 1485.2600 2385.1800 ;
        RECT 1493.4000 2362.9400 1495.0000 2363.4200 ;
        RECT 1493.4000 2368.3800 1495.0000 2368.8600 ;
        RECT 1483.6600 2362.9400 1485.2600 2363.4200 ;
        RECT 1483.6600 2368.3800 1485.2600 2368.8600 ;
        RECT 1438.6600 2401.0200 1440.2600 2401.5000 ;
        RECT 1438.6600 2406.4600 1440.2600 2406.9400 ;
        RECT 1438.6600 2411.9000 1440.2600 2412.3800 ;
        RECT 1438.6600 2390.1400 1440.2600 2390.6200 ;
        RECT 1438.6600 2395.5800 1440.2600 2396.0600 ;
        RECT 1438.6600 2373.8200 1440.2600 2374.3000 ;
        RECT 1438.6600 2379.2600 1440.2600 2379.7400 ;
        RECT 1438.6600 2384.7000 1440.2600 2385.1800 ;
        RECT 1438.6600 2362.9400 1440.2600 2363.4200 ;
        RECT 1438.6600 2368.3800 1440.2600 2368.8600 ;
        RECT 1393.6600 2444.5400 1395.2600 2445.0200 ;
        RECT 1393.6600 2449.9800 1395.2600 2450.4600 ;
        RECT 1393.6600 2455.4200 1395.2600 2455.9000 ;
        RECT 1348.6600 2444.5400 1350.2600 2445.0200 ;
        RECT 1348.6600 2449.9800 1350.2600 2450.4600 ;
        RECT 1348.6600 2455.4200 1350.2600 2455.9000 ;
        RECT 1393.6600 2433.6600 1395.2600 2434.1400 ;
        RECT 1393.6600 2439.1000 1395.2600 2439.5800 ;
        RECT 1393.6600 2417.3400 1395.2600 2417.8200 ;
        RECT 1393.6600 2422.7800 1395.2600 2423.2600 ;
        RECT 1393.6600 2428.2200 1395.2600 2428.7000 ;
        RECT 1348.6600 2433.6600 1350.2600 2434.1400 ;
        RECT 1348.6600 2439.1000 1350.2600 2439.5800 ;
        RECT 1348.6600 2417.3400 1350.2600 2417.8200 ;
        RECT 1348.6600 2422.7800 1350.2600 2423.2600 ;
        RECT 1348.6600 2428.2200 1350.2600 2428.7000 ;
        RECT 1303.6600 2444.5400 1305.2600 2445.0200 ;
        RECT 1303.6600 2449.9800 1305.2600 2450.4600 ;
        RECT 1295.9000 2444.5400 1297.5000 2445.0200 ;
        RECT 1295.9000 2449.9800 1297.5000 2450.4600 ;
        RECT 1295.9000 2455.4200 1297.5000 2455.9000 ;
        RECT 1303.6600 2455.4200 1305.2600 2455.9000 ;
        RECT 1303.6600 2433.6600 1305.2600 2434.1400 ;
        RECT 1303.6600 2439.1000 1305.2600 2439.5800 ;
        RECT 1295.9000 2433.6600 1297.5000 2434.1400 ;
        RECT 1295.9000 2439.1000 1297.5000 2439.5800 ;
        RECT 1303.6600 2417.3400 1305.2600 2417.8200 ;
        RECT 1303.6600 2422.7800 1305.2600 2423.2600 ;
        RECT 1295.9000 2417.3400 1297.5000 2417.8200 ;
        RECT 1295.9000 2422.7800 1297.5000 2423.2600 ;
        RECT 1295.9000 2428.2200 1297.5000 2428.7000 ;
        RECT 1303.6600 2428.2200 1305.2600 2428.7000 ;
        RECT 1393.6600 2401.0200 1395.2600 2401.5000 ;
        RECT 1393.6600 2406.4600 1395.2600 2406.9400 ;
        RECT 1393.6600 2411.9000 1395.2600 2412.3800 ;
        RECT 1393.6600 2390.1400 1395.2600 2390.6200 ;
        RECT 1393.6600 2395.5800 1395.2600 2396.0600 ;
        RECT 1348.6600 2401.0200 1350.2600 2401.5000 ;
        RECT 1348.6600 2406.4600 1350.2600 2406.9400 ;
        RECT 1348.6600 2411.9000 1350.2600 2412.3800 ;
        RECT 1348.6600 2390.1400 1350.2600 2390.6200 ;
        RECT 1348.6600 2395.5800 1350.2600 2396.0600 ;
        RECT 1393.6600 2373.8200 1395.2600 2374.3000 ;
        RECT 1393.6600 2379.2600 1395.2600 2379.7400 ;
        RECT 1393.6600 2384.7000 1395.2600 2385.1800 ;
        RECT 1393.6600 2362.9400 1395.2600 2363.4200 ;
        RECT 1393.6600 2368.3800 1395.2600 2368.8600 ;
        RECT 1348.6600 2373.8200 1350.2600 2374.3000 ;
        RECT 1348.6600 2379.2600 1350.2600 2379.7400 ;
        RECT 1348.6600 2384.7000 1350.2600 2385.1800 ;
        RECT 1348.6600 2362.9400 1350.2600 2363.4200 ;
        RECT 1348.6600 2368.3800 1350.2600 2368.8600 ;
        RECT 1303.6600 2401.0200 1305.2600 2401.5000 ;
        RECT 1303.6600 2406.4600 1305.2600 2406.9400 ;
        RECT 1303.6600 2411.9000 1305.2600 2412.3800 ;
        RECT 1295.9000 2401.0200 1297.5000 2401.5000 ;
        RECT 1295.9000 2406.4600 1297.5000 2406.9400 ;
        RECT 1295.9000 2411.9000 1297.5000 2412.3800 ;
        RECT 1303.6600 2390.1400 1305.2600 2390.6200 ;
        RECT 1303.6600 2395.5800 1305.2600 2396.0600 ;
        RECT 1295.9000 2390.1400 1297.5000 2390.6200 ;
        RECT 1295.9000 2395.5800 1297.5000 2396.0600 ;
        RECT 1303.6600 2373.8200 1305.2600 2374.3000 ;
        RECT 1303.6600 2379.2600 1305.2600 2379.7400 ;
        RECT 1303.6600 2384.7000 1305.2600 2385.1800 ;
        RECT 1295.9000 2373.8200 1297.5000 2374.3000 ;
        RECT 1295.9000 2379.2600 1297.5000 2379.7400 ;
        RECT 1295.9000 2384.7000 1297.5000 2385.1800 ;
        RECT 1303.6600 2362.9400 1305.2600 2363.4200 ;
        RECT 1303.6600 2368.3800 1305.2600 2368.8600 ;
        RECT 1295.9000 2362.9400 1297.5000 2363.4200 ;
        RECT 1295.9000 2368.3800 1297.5000 2368.8600 ;
        RECT 1493.4000 2346.6200 1495.0000 2347.1000 ;
        RECT 1493.4000 2352.0600 1495.0000 2352.5400 ;
        RECT 1493.4000 2357.5000 1495.0000 2357.9800 ;
        RECT 1483.6600 2346.6200 1485.2600 2347.1000 ;
        RECT 1483.6600 2352.0600 1485.2600 2352.5400 ;
        RECT 1483.6600 2357.5000 1485.2600 2357.9800 ;
        RECT 1493.4000 2335.7400 1495.0000 2336.2200 ;
        RECT 1493.4000 2341.1800 1495.0000 2341.6600 ;
        RECT 1483.6600 2335.7400 1485.2600 2336.2200 ;
        RECT 1483.6600 2341.1800 1485.2600 2341.6600 ;
        RECT 1493.4000 2319.4200 1495.0000 2319.9000 ;
        RECT 1493.4000 2324.8600 1495.0000 2325.3400 ;
        RECT 1493.4000 2330.3000 1495.0000 2330.7800 ;
        RECT 1483.6600 2319.4200 1485.2600 2319.9000 ;
        RECT 1483.6600 2324.8600 1485.2600 2325.3400 ;
        RECT 1483.6600 2330.3000 1485.2600 2330.7800 ;
        RECT 1493.4000 2308.5400 1495.0000 2309.0200 ;
        RECT 1493.4000 2313.9800 1495.0000 2314.4600 ;
        RECT 1483.6600 2308.5400 1485.2600 2309.0200 ;
        RECT 1483.6600 2313.9800 1485.2600 2314.4600 ;
        RECT 1438.6600 2346.6200 1440.2600 2347.1000 ;
        RECT 1438.6600 2352.0600 1440.2600 2352.5400 ;
        RECT 1438.6600 2357.5000 1440.2600 2357.9800 ;
        RECT 1438.6600 2335.7400 1440.2600 2336.2200 ;
        RECT 1438.6600 2341.1800 1440.2600 2341.6600 ;
        RECT 1438.6600 2319.4200 1440.2600 2319.9000 ;
        RECT 1438.6600 2324.8600 1440.2600 2325.3400 ;
        RECT 1438.6600 2330.3000 1440.2600 2330.7800 ;
        RECT 1438.6600 2308.5400 1440.2600 2309.0200 ;
        RECT 1438.6600 2313.9800 1440.2600 2314.4600 ;
        RECT 1493.4000 2292.2200 1495.0000 2292.7000 ;
        RECT 1493.4000 2297.6600 1495.0000 2298.1400 ;
        RECT 1493.4000 2303.1000 1495.0000 2303.5800 ;
        RECT 1483.6600 2292.2200 1485.2600 2292.7000 ;
        RECT 1483.6600 2297.6600 1485.2600 2298.1400 ;
        RECT 1483.6600 2303.1000 1485.2600 2303.5800 ;
        RECT 1493.4000 2281.3400 1495.0000 2281.8200 ;
        RECT 1493.4000 2286.7800 1495.0000 2287.2600 ;
        RECT 1483.6600 2281.3400 1485.2600 2281.8200 ;
        RECT 1483.6600 2286.7800 1485.2600 2287.2600 ;
        RECT 1493.4000 2265.0200 1495.0000 2265.5000 ;
        RECT 1493.4000 2270.4600 1495.0000 2270.9400 ;
        RECT 1493.4000 2275.9000 1495.0000 2276.3800 ;
        RECT 1483.6600 2265.0200 1485.2600 2265.5000 ;
        RECT 1483.6600 2270.4600 1485.2600 2270.9400 ;
        RECT 1483.6600 2275.9000 1485.2600 2276.3800 ;
        RECT 1483.6600 2259.5800 1485.2600 2260.0600 ;
        RECT 1493.4000 2259.5800 1495.0000 2260.0600 ;
        RECT 1438.6600 2292.2200 1440.2600 2292.7000 ;
        RECT 1438.6600 2297.6600 1440.2600 2298.1400 ;
        RECT 1438.6600 2303.1000 1440.2600 2303.5800 ;
        RECT 1438.6600 2281.3400 1440.2600 2281.8200 ;
        RECT 1438.6600 2286.7800 1440.2600 2287.2600 ;
        RECT 1438.6600 2265.0200 1440.2600 2265.5000 ;
        RECT 1438.6600 2270.4600 1440.2600 2270.9400 ;
        RECT 1438.6600 2275.9000 1440.2600 2276.3800 ;
        RECT 1438.6600 2259.5800 1440.2600 2260.0600 ;
        RECT 1393.6600 2346.6200 1395.2600 2347.1000 ;
        RECT 1393.6600 2352.0600 1395.2600 2352.5400 ;
        RECT 1393.6600 2357.5000 1395.2600 2357.9800 ;
        RECT 1393.6600 2335.7400 1395.2600 2336.2200 ;
        RECT 1393.6600 2341.1800 1395.2600 2341.6600 ;
        RECT 1348.6600 2346.6200 1350.2600 2347.1000 ;
        RECT 1348.6600 2352.0600 1350.2600 2352.5400 ;
        RECT 1348.6600 2357.5000 1350.2600 2357.9800 ;
        RECT 1348.6600 2335.7400 1350.2600 2336.2200 ;
        RECT 1348.6600 2341.1800 1350.2600 2341.6600 ;
        RECT 1393.6600 2319.4200 1395.2600 2319.9000 ;
        RECT 1393.6600 2324.8600 1395.2600 2325.3400 ;
        RECT 1393.6600 2330.3000 1395.2600 2330.7800 ;
        RECT 1393.6600 2308.5400 1395.2600 2309.0200 ;
        RECT 1393.6600 2313.9800 1395.2600 2314.4600 ;
        RECT 1348.6600 2319.4200 1350.2600 2319.9000 ;
        RECT 1348.6600 2324.8600 1350.2600 2325.3400 ;
        RECT 1348.6600 2330.3000 1350.2600 2330.7800 ;
        RECT 1348.6600 2308.5400 1350.2600 2309.0200 ;
        RECT 1348.6600 2313.9800 1350.2600 2314.4600 ;
        RECT 1303.6600 2346.6200 1305.2600 2347.1000 ;
        RECT 1303.6600 2352.0600 1305.2600 2352.5400 ;
        RECT 1303.6600 2357.5000 1305.2600 2357.9800 ;
        RECT 1295.9000 2346.6200 1297.5000 2347.1000 ;
        RECT 1295.9000 2352.0600 1297.5000 2352.5400 ;
        RECT 1295.9000 2357.5000 1297.5000 2357.9800 ;
        RECT 1303.6600 2335.7400 1305.2600 2336.2200 ;
        RECT 1303.6600 2341.1800 1305.2600 2341.6600 ;
        RECT 1295.9000 2335.7400 1297.5000 2336.2200 ;
        RECT 1295.9000 2341.1800 1297.5000 2341.6600 ;
        RECT 1303.6600 2319.4200 1305.2600 2319.9000 ;
        RECT 1303.6600 2324.8600 1305.2600 2325.3400 ;
        RECT 1303.6600 2330.3000 1305.2600 2330.7800 ;
        RECT 1295.9000 2319.4200 1297.5000 2319.9000 ;
        RECT 1295.9000 2324.8600 1297.5000 2325.3400 ;
        RECT 1295.9000 2330.3000 1297.5000 2330.7800 ;
        RECT 1303.6600 2308.5400 1305.2600 2309.0200 ;
        RECT 1303.6600 2313.9800 1305.2600 2314.4600 ;
        RECT 1295.9000 2308.5400 1297.5000 2309.0200 ;
        RECT 1295.9000 2313.9800 1297.5000 2314.4600 ;
        RECT 1393.6600 2292.2200 1395.2600 2292.7000 ;
        RECT 1393.6600 2297.6600 1395.2600 2298.1400 ;
        RECT 1393.6600 2303.1000 1395.2600 2303.5800 ;
        RECT 1393.6600 2281.3400 1395.2600 2281.8200 ;
        RECT 1393.6600 2286.7800 1395.2600 2287.2600 ;
        RECT 1348.6600 2292.2200 1350.2600 2292.7000 ;
        RECT 1348.6600 2297.6600 1350.2600 2298.1400 ;
        RECT 1348.6600 2303.1000 1350.2600 2303.5800 ;
        RECT 1348.6600 2281.3400 1350.2600 2281.8200 ;
        RECT 1348.6600 2286.7800 1350.2600 2287.2600 ;
        RECT 1393.6600 2265.0200 1395.2600 2265.5000 ;
        RECT 1393.6600 2270.4600 1395.2600 2270.9400 ;
        RECT 1393.6600 2275.9000 1395.2600 2276.3800 ;
        RECT 1393.6600 2259.5800 1395.2600 2260.0600 ;
        RECT 1348.6600 2265.0200 1350.2600 2265.5000 ;
        RECT 1348.6600 2270.4600 1350.2600 2270.9400 ;
        RECT 1348.6600 2275.9000 1350.2600 2276.3800 ;
        RECT 1348.6600 2259.5800 1350.2600 2260.0600 ;
        RECT 1303.6600 2292.2200 1305.2600 2292.7000 ;
        RECT 1303.6600 2297.6600 1305.2600 2298.1400 ;
        RECT 1303.6600 2303.1000 1305.2600 2303.5800 ;
        RECT 1295.9000 2292.2200 1297.5000 2292.7000 ;
        RECT 1295.9000 2297.6600 1297.5000 2298.1400 ;
        RECT 1295.9000 2303.1000 1297.5000 2303.5800 ;
        RECT 1303.6600 2281.3400 1305.2600 2281.8200 ;
        RECT 1303.6600 2286.7800 1305.2600 2287.2600 ;
        RECT 1295.9000 2281.3400 1297.5000 2281.8200 ;
        RECT 1295.9000 2286.7800 1297.5000 2287.2600 ;
        RECT 1303.6600 2265.0200 1305.2600 2265.5000 ;
        RECT 1303.6600 2270.4600 1305.2600 2270.9400 ;
        RECT 1303.6600 2275.9000 1305.2600 2276.3800 ;
        RECT 1295.9000 2265.0200 1297.5000 2265.5000 ;
        RECT 1295.9000 2270.4600 1297.5000 2270.9400 ;
        RECT 1295.9000 2275.9000 1297.5000 2276.3800 ;
        RECT 1295.9000 2259.5800 1297.5000 2260.0600 ;
        RECT 1303.6600 2259.5800 1305.2600 2260.0600 ;
        RECT 1290.3400 2461.8900 1500.5600 2463.4900 ;
        RECT 1290.3400 2255.3900 1500.5600 2256.9900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 2249.9600 1297.5000 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 2468.0000 1297.5000 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 2249.9600 1495.0000 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 2468.0000 1495.0000 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2255.3900 1291.9400 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2255.3900 1500.5600 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2461.8900 1291.9400 2463.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2461.8900 1500.5600 2463.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 2025.7500 1485.2600 2233.8500 ;
        RECT 1438.6600 2025.7500 1440.2600 2233.8500 ;
        RECT 1393.6600 2025.7500 1395.2600 2233.8500 ;
        RECT 1348.6600 2025.7500 1350.2600 2233.8500 ;
        RECT 1303.6600 2025.7500 1305.2600 2233.8500 ;
        RECT 1493.4000 2020.3200 1495.0000 2239.9600 ;
        RECT 1295.9000 2020.3200 1297.5000 2239.9600 ;
      LAYER met3 ;
        RECT 1493.4000 2214.9000 1495.0000 2215.3800 ;
        RECT 1493.4000 2220.3400 1495.0000 2220.8200 ;
        RECT 1483.6600 2214.9000 1485.2600 2215.3800 ;
        RECT 1483.6600 2220.3400 1485.2600 2220.8200 ;
        RECT 1483.6600 2225.7800 1485.2600 2226.2600 ;
        RECT 1493.4000 2225.7800 1495.0000 2226.2600 ;
        RECT 1493.4000 2204.0200 1495.0000 2204.5000 ;
        RECT 1493.4000 2209.4600 1495.0000 2209.9400 ;
        RECT 1483.6600 2204.0200 1485.2600 2204.5000 ;
        RECT 1483.6600 2209.4600 1485.2600 2209.9400 ;
        RECT 1493.4000 2187.7000 1495.0000 2188.1800 ;
        RECT 1493.4000 2193.1400 1495.0000 2193.6200 ;
        RECT 1483.6600 2187.7000 1485.2600 2188.1800 ;
        RECT 1483.6600 2193.1400 1485.2600 2193.6200 ;
        RECT 1483.6600 2198.5800 1485.2600 2199.0600 ;
        RECT 1493.4000 2198.5800 1495.0000 2199.0600 ;
        RECT 1438.6600 2214.9000 1440.2600 2215.3800 ;
        RECT 1438.6600 2220.3400 1440.2600 2220.8200 ;
        RECT 1438.6600 2225.7800 1440.2600 2226.2600 ;
        RECT 1438.6600 2204.0200 1440.2600 2204.5000 ;
        RECT 1438.6600 2209.4600 1440.2600 2209.9400 ;
        RECT 1438.6600 2187.7000 1440.2600 2188.1800 ;
        RECT 1438.6600 2193.1400 1440.2600 2193.6200 ;
        RECT 1438.6600 2198.5800 1440.2600 2199.0600 ;
        RECT 1493.4000 2171.3800 1495.0000 2171.8600 ;
        RECT 1493.4000 2176.8200 1495.0000 2177.3000 ;
        RECT 1493.4000 2182.2600 1495.0000 2182.7400 ;
        RECT 1483.6600 2171.3800 1485.2600 2171.8600 ;
        RECT 1483.6600 2176.8200 1485.2600 2177.3000 ;
        RECT 1483.6600 2182.2600 1485.2600 2182.7400 ;
        RECT 1493.4000 2160.5000 1495.0000 2160.9800 ;
        RECT 1493.4000 2165.9400 1495.0000 2166.4200 ;
        RECT 1483.6600 2160.5000 1485.2600 2160.9800 ;
        RECT 1483.6600 2165.9400 1485.2600 2166.4200 ;
        RECT 1493.4000 2144.1800 1495.0000 2144.6600 ;
        RECT 1493.4000 2149.6200 1495.0000 2150.1000 ;
        RECT 1493.4000 2155.0600 1495.0000 2155.5400 ;
        RECT 1483.6600 2144.1800 1485.2600 2144.6600 ;
        RECT 1483.6600 2149.6200 1485.2600 2150.1000 ;
        RECT 1483.6600 2155.0600 1485.2600 2155.5400 ;
        RECT 1493.4000 2133.3000 1495.0000 2133.7800 ;
        RECT 1493.4000 2138.7400 1495.0000 2139.2200 ;
        RECT 1483.6600 2133.3000 1485.2600 2133.7800 ;
        RECT 1483.6600 2138.7400 1485.2600 2139.2200 ;
        RECT 1438.6600 2171.3800 1440.2600 2171.8600 ;
        RECT 1438.6600 2176.8200 1440.2600 2177.3000 ;
        RECT 1438.6600 2182.2600 1440.2600 2182.7400 ;
        RECT 1438.6600 2160.5000 1440.2600 2160.9800 ;
        RECT 1438.6600 2165.9400 1440.2600 2166.4200 ;
        RECT 1438.6600 2144.1800 1440.2600 2144.6600 ;
        RECT 1438.6600 2149.6200 1440.2600 2150.1000 ;
        RECT 1438.6600 2155.0600 1440.2600 2155.5400 ;
        RECT 1438.6600 2133.3000 1440.2600 2133.7800 ;
        RECT 1438.6600 2138.7400 1440.2600 2139.2200 ;
        RECT 1393.6600 2214.9000 1395.2600 2215.3800 ;
        RECT 1393.6600 2220.3400 1395.2600 2220.8200 ;
        RECT 1393.6600 2225.7800 1395.2600 2226.2600 ;
        RECT 1348.6600 2214.9000 1350.2600 2215.3800 ;
        RECT 1348.6600 2220.3400 1350.2600 2220.8200 ;
        RECT 1348.6600 2225.7800 1350.2600 2226.2600 ;
        RECT 1393.6600 2204.0200 1395.2600 2204.5000 ;
        RECT 1393.6600 2209.4600 1395.2600 2209.9400 ;
        RECT 1393.6600 2187.7000 1395.2600 2188.1800 ;
        RECT 1393.6600 2193.1400 1395.2600 2193.6200 ;
        RECT 1393.6600 2198.5800 1395.2600 2199.0600 ;
        RECT 1348.6600 2204.0200 1350.2600 2204.5000 ;
        RECT 1348.6600 2209.4600 1350.2600 2209.9400 ;
        RECT 1348.6600 2187.7000 1350.2600 2188.1800 ;
        RECT 1348.6600 2193.1400 1350.2600 2193.6200 ;
        RECT 1348.6600 2198.5800 1350.2600 2199.0600 ;
        RECT 1303.6600 2214.9000 1305.2600 2215.3800 ;
        RECT 1303.6600 2220.3400 1305.2600 2220.8200 ;
        RECT 1295.9000 2214.9000 1297.5000 2215.3800 ;
        RECT 1295.9000 2220.3400 1297.5000 2220.8200 ;
        RECT 1295.9000 2225.7800 1297.5000 2226.2600 ;
        RECT 1303.6600 2225.7800 1305.2600 2226.2600 ;
        RECT 1303.6600 2204.0200 1305.2600 2204.5000 ;
        RECT 1303.6600 2209.4600 1305.2600 2209.9400 ;
        RECT 1295.9000 2204.0200 1297.5000 2204.5000 ;
        RECT 1295.9000 2209.4600 1297.5000 2209.9400 ;
        RECT 1303.6600 2187.7000 1305.2600 2188.1800 ;
        RECT 1303.6600 2193.1400 1305.2600 2193.6200 ;
        RECT 1295.9000 2187.7000 1297.5000 2188.1800 ;
        RECT 1295.9000 2193.1400 1297.5000 2193.6200 ;
        RECT 1295.9000 2198.5800 1297.5000 2199.0600 ;
        RECT 1303.6600 2198.5800 1305.2600 2199.0600 ;
        RECT 1393.6600 2171.3800 1395.2600 2171.8600 ;
        RECT 1393.6600 2176.8200 1395.2600 2177.3000 ;
        RECT 1393.6600 2182.2600 1395.2600 2182.7400 ;
        RECT 1393.6600 2160.5000 1395.2600 2160.9800 ;
        RECT 1393.6600 2165.9400 1395.2600 2166.4200 ;
        RECT 1348.6600 2171.3800 1350.2600 2171.8600 ;
        RECT 1348.6600 2176.8200 1350.2600 2177.3000 ;
        RECT 1348.6600 2182.2600 1350.2600 2182.7400 ;
        RECT 1348.6600 2160.5000 1350.2600 2160.9800 ;
        RECT 1348.6600 2165.9400 1350.2600 2166.4200 ;
        RECT 1393.6600 2144.1800 1395.2600 2144.6600 ;
        RECT 1393.6600 2149.6200 1395.2600 2150.1000 ;
        RECT 1393.6600 2155.0600 1395.2600 2155.5400 ;
        RECT 1393.6600 2133.3000 1395.2600 2133.7800 ;
        RECT 1393.6600 2138.7400 1395.2600 2139.2200 ;
        RECT 1348.6600 2144.1800 1350.2600 2144.6600 ;
        RECT 1348.6600 2149.6200 1350.2600 2150.1000 ;
        RECT 1348.6600 2155.0600 1350.2600 2155.5400 ;
        RECT 1348.6600 2133.3000 1350.2600 2133.7800 ;
        RECT 1348.6600 2138.7400 1350.2600 2139.2200 ;
        RECT 1303.6600 2171.3800 1305.2600 2171.8600 ;
        RECT 1303.6600 2176.8200 1305.2600 2177.3000 ;
        RECT 1303.6600 2182.2600 1305.2600 2182.7400 ;
        RECT 1295.9000 2171.3800 1297.5000 2171.8600 ;
        RECT 1295.9000 2176.8200 1297.5000 2177.3000 ;
        RECT 1295.9000 2182.2600 1297.5000 2182.7400 ;
        RECT 1303.6600 2160.5000 1305.2600 2160.9800 ;
        RECT 1303.6600 2165.9400 1305.2600 2166.4200 ;
        RECT 1295.9000 2160.5000 1297.5000 2160.9800 ;
        RECT 1295.9000 2165.9400 1297.5000 2166.4200 ;
        RECT 1303.6600 2144.1800 1305.2600 2144.6600 ;
        RECT 1303.6600 2149.6200 1305.2600 2150.1000 ;
        RECT 1303.6600 2155.0600 1305.2600 2155.5400 ;
        RECT 1295.9000 2144.1800 1297.5000 2144.6600 ;
        RECT 1295.9000 2149.6200 1297.5000 2150.1000 ;
        RECT 1295.9000 2155.0600 1297.5000 2155.5400 ;
        RECT 1303.6600 2133.3000 1305.2600 2133.7800 ;
        RECT 1303.6600 2138.7400 1305.2600 2139.2200 ;
        RECT 1295.9000 2133.3000 1297.5000 2133.7800 ;
        RECT 1295.9000 2138.7400 1297.5000 2139.2200 ;
        RECT 1493.4000 2116.9800 1495.0000 2117.4600 ;
        RECT 1493.4000 2122.4200 1495.0000 2122.9000 ;
        RECT 1493.4000 2127.8600 1495.0000 2128.3400 ;
        RECT 1483.6600 2116.9800 1485.2600 2117.4600 ;
        RECT 1483.6600 2122.4200 1485.2600 2122.9000 ;
        RECT 1483.6600 2127.8600 1485.2600 2128.3400 ;
        RECT 1493.4000 2106.1000 1495.0000 2106.5800 ;
        RECT 1493.4000 2111.5400 1495.0000 2112.0200 ;
        RECT 1483.6600 2106.1000 1485.2600 2106.5800 ;
        RECT 1483.6600 2111.5400 1485.2600 2112.0200 ;
        RECT 1493.4000 2089.7800 1495.0000 2090.2600 ;
        RECT 1493.4000 2095.2200 1495.0000 2095.7000 ;
        RECT 1493.4000 2100.6600 1495.0000 2101.1400 ;
        RECT 1483.6600 2089.7800 1485.2600 2090.2600 ;
        RECT 1483.6600 2095.2200 1485.2600 2095.7000 ;
        RECT 1483.6600 2100.6600 1485.2600 2101.1400 ;
        RECT 1493.4000 2078.9000 1495.0000 2079.3800 ;
        RECT 1493.4000 2084.3400 1495.0000 2084.8200 ;
        RECT 1483.6600 2078.9000 1485.2600 2079.3800 ;
        RECT 1483.6600 2084.3400 1485.2600 2084.8200 ;
        RECT 1438.6600 2116.9800 1440.2600 2117.4600 ;
        RECT 1438.6600 2122.4200 1440.2600 2122.9000 ;
        RECT 1438.6600 2127.8600 1440.2600 2128.3400 ;
        RECT 1438.6600 2106.1000 1440.2600 2106.5800 ;
        RECT 1438.6600 2111.5400 1440.2600 2112.0200 ;
        RECT 1438.6600 2089.7800 1440.2600 2090.2600 ;
        RECT 1438.6600 2095.2200 1440.2600 2095.7000 ;
        RECT 1438.6600 2100.6600 1440.2600 2101.1400 ;
        RECT 1438.6600 2078.9000 1440.2600 2079.3800 ;
        RECT 1438.6600 2084.3400 1440.2600 2084.8200 ;
        RECT 1493.4000 2062.5800 1495.0000 2063.0600 ;
        RECT 1493.4000 2068.0200 1495.0000 2068.5000 ;
        RECT 1493.4000 2073.4600 1495.0000 2073.9400 ;
        RECT 1483.6600 2062.5800 1485.2600 2063.0600 ;
        RECT 1483.6600 2068.0200 1485.2600 2068.5000 ;
        RECT 1483.6600 2073.4600 1485.2600 2073.9400 ;
        RECT 1493.4000 2051.7000 1495.0000 2052.1800 ;
        RECT 1493.4000 2057.1400 1495.0000 2057.6200 ;
        RECT 1483.6600 2051.7000 1485.2600 2052.1800 ;
        RECT 1483.6600 2057.1400 1485.2600 2057.6200 ;
        RECT 1493.4000 2035.3800 1495.0000 2035.8600 ;
        RECT 1493.4000 2040.8200 1495.0000 2041.3000 ;
        RECT 1493.4000 2046.2600 1495.0000 2046.7400 ;
        RECT 1483.6600 2035.3800 1485.2600 2035.8600 ;
        RECT 1483.6600 2040.8200 1485.2600 2041.3000 ;
        RECT 1483.6600 2046.2600 1485.2600 2046.7400 ;
        RECT 1483.6600 2029.9400 1485.2600 2030.4200 ;
        RECT 1493.4000 2029.9400 1495.0000 2030.4200 ;
        RECT 1438.6600 2062.5800 1440.2600 2063.0600 ;
        RECT 1438.6600 2068.0200 1440.2600 2068.5000 ;
        RECT 1438.6600 2073.4600 1440.2600 2073.9400 ;
        RECT 1438.6600 2051.7000 1440.2600 2052.1800 ;
        RECT 1438.6600 2057.1400 1440.2600 2057.6200 ;
        RECT 1438.6600 2035.3800 1440.2600 2035.8600 ;
        RECT 1438.6600 2040.8200 1440.2600 2041.3000 ;
        RECT 1438.6600 2046.2600 1440.2600 2046.7400 ;
        RECT 1438.6600 2029.9400 1440.2600 2030.4200 ;
        RECT 1393.6600 2116.9800 1395.2600 2117.4600 ;
        RECT 1393.6600 2122.4200 1395.2600 2122.9000 ;
        RECT 1393.6600 2127.8600 1395.2600 2128.3400 ;
        RECT 1393.6600 2106.1000 1395.2600 2106.5800 ;
        RECT 1393.6600 2111.5400 1395.2600 2112.0200 ;
        RECT 1348.6600 2116.9800 1350.2600 2117.4600 ;
        RECT 1348.6600 2122.4200 1350.2600 2122.9000 ;
        RECT 1348.6600 2127.8600 1350.2600 2128.3400 ;
        RECT 1348.6600 2106.1000 1350.2600 2106.5800 ;
        RECT 1348.6600 2111.5400 1350.2600 2112.0200 ;
        RECT 1393.6600 2089.7800 1395.2600 2090.2600 ;
        RECT 1393.6600 2095.2200 1395.2600 2095.7000 ;
        RECT 1393.6600 2100.6600 1395.2600 2101.1400 ;
        RECT 1393.6600 2078.9000 1395.2600 2079.3800 ;
        RECT 1393.6600 2084.3400 1395.2600 2084.8200 ;
        RECT 1348.6600 2089.7800 1350.2600 2090.2600 ;
        RECT 1348.6600 2095.2200 1350.2600 2095.7000 ;
        RECT 1348.6600 2100.6600 1350.2600 2101.1400 ;
        RECT 1348.6600 2078.9000 1350.2600 2079.3800 ;
        RECT 1348.6600 2084.3400 1350.2600 2084.8200 ;
        RECT 1303.6600 2116.9800 1305.2600 2117.4600 ;
        RECT 1303.6600 2122.4200 1305.2600 2122.9000 ;
        RECT 1303.6600 2127.8600 1305.2600 2128.3400 ;
        RECT 1295.9000 2116.9800 1297.5000 2117.4600 ;
        RECT 1295.9000 2122.4200 1297.5000 2122.9000 ;
        RECT 1295.9000 2127.8600 1297.5000 2128.3400 ;
        RECT 1303.6600 2106.1000 1305.2600 2106.5800 ;
        RECT 1303.6600 2111.5400 1305.2600 2112.0200 ;
        RECT 1295.9000 2106.1000 1297.5000 2106.5800 ;
        RECT 1295.9000 2111.5400 1297.5000 2112.0200 ;
        RECT 1303.6600 2089.7800 1305.2600 2090.2600 ;
        RECT 1303.6600 2095.2200 1305.2600 2095.7000 ;
        RECT 1303.6600 2100.6600 1305.2600 2101.1400 ;
        RECT 1295.9000 2089.7800 1297.5000 2090.2600 ;
        RECT 1295.9000 2095.2200 1297.5000 2095.7000 ;
        RECT 1295.9000 2100.6600 1297.5000 2101.1400 ;
        RECT 1303.6600 2078.9000 1305.2600 2079.3800 ;
        RECT 1303.6600 2084.3400 1305.2600 2084.8200 ;
        RECT 1295.9000 2078.9000 1297.5000 2079.3800 ;
        RECT 1295.9000 2084.3400 1297.5000 2084.8200 ;
        RECT 1393.6600 2062.5800 1395.2600 2063.0600 ;
        RECT 1393.6600 2068.0200 1395.2600 2068.5000 ;
        RECT 1393.6600 2073.4600 1395.2600 2073.9400 ;
        RECT 1393.6600 2051.7000 1395.2600 2052.1800 ;
        RECT 1393.6600 2057.1400 1395.2600 2057.6200 ;
        RECT 1348.6600 2062.5800 1350.2600 2063.0600 ;
        RECT 1348.6600 2068.0200 1350.2600 2068.5000 ;
        RECT 1348.6600 2073.4600 1350.2600 2073.9400 ;
        RECT 1348.6600 2051.7000 1350.2600 2052.1800 ;
        RECT 1348.6600 2057.1400 1350.2600 2057.6200 ;
        RECT 1393.6600 2035.3800 1395.2600 2035.8600 ;
        RECT 1393.6600 2040.8200 1395.2600 2041.3000 ;
        RECT 1393.6600 2046.2600 1395.2600 2046.7400 ;
        RECT 1393.6600 2029.9400 1395.2600 2030.4200 ;
        RECT 1348.6600 2035.3800 1350.2600 2035.8600 ;
        RECT 1348.6600 2040.8200 1350.2600 2041.3000 ;
        RECT 1348.6600 2046.2600 1350.2600 2046.7400 ;
        RECT 1348.6600 2029.9400 1350.2600 2030.4200 ;
        RECT 1303.6600 2062.5800 1305.2600 2063.0600 ;
        RECT 1303.6600 2068.0200 1305.2600 2068.5000 ;
        RECT 1303.6600 2073.4600 1305.2600 2073.9400 ;
        RECT 1295.9000 2062.5800 1297.5000 2063.0600 ;
        RECT 1295.9000 2068.0200 1297.5000 2068.5000 ;
        RECT 1295.9000 2073.4600 1297.5000 2073.9400 ;
        RECT 1303.6600 2051.7000 1305.2600 2052.1800 ;
        RECT 1303.6600 2057.1400 1305.2600 2057.6200 ;
        RECT 1295.9000 2051.7000 1297.5000 2052.1800 ;
        RECT 1295.9000 2057.1400 1297.5000 2057.6200 ;
        RECT 1303.6600 2035.3800 1305.2600 2035.8600 ;
        RECT 1303.6600 2040.8200 1305.2600 2041.3000 ;
        RECT 1303.6600 2046.2600 1305.2600 2046.7400 ;
        RECT 1295.9000 2035.3800 1297.5000 2035.8600 ;
        RECT 1295.9000 2040.8200 1297.5000 2041.3000 ;
        RECT 1295.9000 2046.2600 1297.5000 2046.7400 ;
        RECT 1295.9000 2029.9400 1297.5000 2030.4200 ;
        RECT 1303.6600 2029.9400 1305.2600 2030.4200 ;
        RECT 1290.3400 2232.2500 1500.5600 2233.8500 ;
        RECT 1290.3400 2025.7500 1500.5600 2027.3500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 2020.3200 1297.5000 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 2238.3600 1297.5000 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 2020.3200 1495.0000 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 2238.3600 1495.0000 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2025.7500 1291.9400 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2025.7500 1500.5600 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2232.2500 1291.9400 2233.8500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2232.2500 1500.5600 2233.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 1796.1100 1485.2600 2004.2100 ;
        RECT 1438.6600 1796.1100 1440.2600 2004.2100 ;
        RECT 1393.6600 1796.1100 1395.2600 2004.2100 ;
        RECT 1348.6600 1796.1100 1350.2600 2004.2100 ;
        RECT 1303.6600 1796.1100 1305.2600 2004.2100 ;
        RECT 1493.4000 1790.6800 1495.0000 2010.3200 ;
        RECT 1295.9000 1790.6800 1297.5000 2010.3200 ;
      LAYER met3 ;
        RECT 1493.4000 1985.2600 1495.0000 1985.7400 ;
        RECT 1493.4000 1990.7000 1495.0000 1991.1800 ;
        RECT 1483.6600 1985.2600 1485.2600 1985.7400 ;
        RECT 1483.6600 1990.7000 1485.2600 1991.1800 ;
        RECT 1483.6600 1996.1400 1485.2600 1996.6200 ;
        RECT 1493.4000 1996.1400 1495.0000 1996.6200 ;
        RECT 1493.4000 1974.3800 1495.0000 1974.8600 ;
        RECT 1493.4000 1979.8200 1495.0000 1980.3000 ;
        RECT 1483.6600 1974.3800 1485.2600 1974.8600 ;
        RECT 1483.6600 1979.8200 1485.2600 1980.3000 ;
        RECT 1493.4000 1958.0600 1495.0000 1958.5400 ;
        RECT 1493.4000 1963.5000 1495.0000 1963.9800 ;
        RECT 1483.6600 1958.0600 1485.2600 1958.5400 ;
        RECT 1483.6600 1963.5000 1485.2600 1963.9800 ;
        RECT 1483.6600 1968.9400 1485.2600 1969.4200 ;
        RECT 1493.4000 1968.9400 1495.0000 1969.4200 ;
        RECT 1438.6600 1985.2600 1440.2600 1985.7400 ;
        RECT 1438.6600 1990.7000 1440.2600 1991.1800 ;
        RECT 1438.6600 1996.1400 1440.2600 1996.6200 ;
        RECT 1438.6600 1974.3800 1440.2600 1974.8600 ;
        RECT 1438.6600 1979.8200 1440.2600 1980.3000 ;
        RECT 1438.6600 1958.0600 1440.2600 1958.5400 ;
        RECT 1438.6600 1963.5000 1440.2600 1963.9800 ;
        RECT 1438.6600 1968.9400 1440.2600 1969.4200 ;
        RECT 1493.4000 1941.7400 1495.0000 1942.2200 ;
        RECT 1493.4000 1947.1800 1495.0000 1947.6600 ;
        RECT 1493.4000 1952.6200 1495.0000 1953.1000 ;
        RECT 1483.6600 1941.7400 1485.2600 1942.2200 ;
        RECT 1483.6600 1947.1800 1485.2600 1947.6600 ;
        RECT 1483.6600 1952.6200 1485.2600 1953.1000 ;
        RECT 1493.4000 1930.8600 1495.0000 1931.3400 ;
        RECT 1493.4000 1936.3000 1495.0000 1936.7800 ;
        RECT 1483.6600 1930.8600 1485.2600 1931.3400 ;
        RECT 1483.6600 1936.3000 1485.2600 1936.7800 ;
        RECT 1493.4000 1914.5400 1495.0000 1915.0200 ;
        RECT 1493.4000 1919.9800 1495.0000 1920.4600 ;
        RECT 1493.4000 1925.4200 1495.0000 1925.9000 ;
        RECT 1483.6600 1914.5400 1485.2600 1915.0200 ;
        RECT 1483.6600 1919.9800 1485.2600 1920.4600 ;
        RECT 1483.6600 1925.4200 1485.2600 1925.9000 ;
        RECT 1493.4000 1903.6600 1495.0000 1904.1400 ;
        RECT 1493.4000 1909.1000 1495.0000 1909.5800 ;
        RECT 1483.6600 1903.6600 1485.2600 1904.1400 ;
        RECT 1483.6600 1909.1000 1485.2600 1909.5800 ;
        RECT 1438.6600 1941.7400 1440.2600 1942.2200 ;
        RECT 1438.6600 1947.1800 1440.2600 1947.6600 ;
        RECT 1438.6600 1952.6200 1440.2600 1953.1000 ;
        RECT 1438.6600 1930.8600 1440.2600 1931.3400 ;
        RECT 1438.6600 1936.3000 1440.2600 1936.7800 ;
        RECT 1438.6600 1914.5400 1440.2600 1915.0200 ;
        RECT 1438.6600 1919.9800 1440.2600 1920.4600 ;
        RECT 1438.6600 1925.4200 1440.2600 1925.9000 ;
        RECT 1438.6600 1903.6600 1440.2600 1904.1400 ;
        RECT 1438.6600 1909.1000 1440.2600 1909.5800 ;
        RECT 1393.6600 1985.2600 1395.2600 1985.7400 ;
        RECT 1393.6600 1990.7000 1395.2600 1991.1800 ;
        RECT 1393.6600 1996.1400 1395.2600 1996.6200 ;
        RECT 1348.6600 1985.2600 1350.2600 1985.7400 ;
        RECT 1348.6600 1990.7000 1350.2600 1991.1800 ;
        RECT 1348.6600 1996.1400 1350.2600 1996.6200 ;
        RECT 1393.6600 1974.3800 1395.2600 1974.8600 ;
        RECT 1393.6600 1979.8200 1395.2600 1980.3000 ;
        RECT 1393.6600 1958.0600 1395.2600 1958.5400 ;
        RECT 1393.6600 1963.5000 1395.2600 1963.9800 ;
        RECT 1393.6600 1968.9400 1395.2600 1969.4200 ;
        RECT 1348.6600 1974.3800 1350.2600 1974.8600 ;
        RECT 1348.6600 1979.8200 1350.2600 1980.3000 ;
        RECT 1348.6600 1958.0600 1350.2600 1958.5400 ;
        RECT 1348.6600 1963.5000 1350.2600 1963.9800 ;
        RECT 1348.6600 1968.9400 1350.2600 1969.4200 ;
        RECT 1303.6600 1985.2600 1305.2600 1985.7400 ;
        RECT 1303.6600 1990.7000 1305.2600 1991.1800 ;
        RECT 1295.9000 1985.2600 1297.5000 1985.7400 ;
        RECT 1295.9000 1990.7000 1297.5000 1991.1800 ;
        RECT 1295.9000 1996.1400 1297.5000 1996.6200 ;
        RECT 1303.6600 1996.1400 1305.2600 1996.6200 ;
        RECT 1303.6600 1974.3800 1305.2600 1974.8600 ;
        RECT 1303.6600 1979.8200 1305.2600 1980.3000 ;
        RECT 1295.9000 1974.3800 1297.5000 1974.8600 ;
        RECT 1295.9000 1979.8200 1297.5000 1980.3000 ;
        RECT 1303.6600 1958.0600 1305.2600 1958.5400 ;
        RECT 1303.6600 1963.5000 1305.2600 1963.9800 ;
        RECT 1295.9000 1958.0600 1297.5000 1958.5400 ;
        RECT 1295.9000 1963.5000 1297.5000 1963.9800 ;
        RECT 1295.9000 1968.9400 1297.5000 1969.4200 ;
        RECT 1303.6600 1968.9400 1305.2600 1969.4200 ;
        RECT 1393.6600 1941.7400 1395.2600 1942.2200 ;
        RECT 1393.6600 1947.1800 1395.2600 1947.6600 ;
        RECT 1393.6600 1952.6200 1395.2600 1953.1000 ;
        RECT 1393.6600 1930.8600 1395.2600 1931.3400 ;
        RECT 1393.6600 1936.3000 1395.2600 1936.7800 ;
        RECT 1348.6600 1941.7400 1350.2600 1942.2200 ;
        RECT 1348.6600 1947.1800 1350.2600 1947.6600 ;
        RECT 1348.6600 1952.6200 1350.2600 1953.1000 ;
        RECT 1348.6600 1930.8600 1350.2600 1931.3400 ;
        RECT 1348.6600 1936.3000 1350.2600 1936.7800 ;
        RECT 1393.6600 1914.5400 1395.2600 1915.0200 ;
        RECT 1393.6600 1919.9800 1395.2600 1920.4600 ;
        RECT 1393.6600 1925.4200 1395.2600 1925.9000 ;
        RECT 1393.6600 1903.6600 1395.2600 1904.1400 ;
        RECT 1393.6600 1909.1000 1395.2600 1909.5800 ;
        RECT 1348.6600 1914.5400 1350.2600 1915.0200 ;
        RECT 1348.6600 1919.9800 1350.2600 1920.4600 ;
        RECT 1348.6600 1925.4200 1350.2600 1925.9000 ;
        RECT 1348.6600 1903.6600 1350.2600 1904.1400 ;
        RECT 1348.6600 1909.1000 1350.2600 1909.5800 ;
        RECT 1303.6600 1941.7400 1305.2600 1942.2200 ;
        RECT 1303.6600 1947.1800 1305.2600 1947.6600 ;
        RECT 1303.6600 1952.6200 1305.2600 1953.1000 ;
        RECT 1295.9000 1941.7400 1297.5000 1942.2200 ;
        RECT 1295.9000 1947.1800 1297.5000 1947.6600 ;
        RECT 1295.9000 1952.6200 1297.5000 1953.1000 ;
        RECT 1303.6600 1930.8600 1305.2600 1931.3400 ;
        RECT 1303.6600 1936.3000 1305.2600 1936.7800 ;
        RECT 1295.9000 1930.8600 1297.5000 1931.3400 ;
        RECT 1295.9000 1936.3000 1297.5000 1936.7800 ;
        RECT 1303.6600 1914.5400 1305.2600 1915.0200 ;
        RECT 1303.6600 1919.9800 1305.2600 1920.4600 ;
        RECT 1303.6600 1925.4200 1305.2600 1925.9000 ;
        RECT 1295.9000 1914.5400 1297.5000 1915.0200 ;
        RECT 1295.9000 1919.9800 1297.5000 1920.4600 ;
        RECT 1295.9000 1925.4200 1297.5000 1925.9000 ;
        RECT 1303.6600 1903.6600 1305.2600 1904.1400 ;
        RECT 1303.6600 1909.1000 1305.2600 1909.5800 ;
        RECT 1295.9000 1903.6600 1297.5000 1904.1400 ;
        RECT 1295.9000 1909.1000 1297.5000 1909.5800 ;
        RECT 1493.4000 1887.3400 1495.0000 1887.8200 ;
        RECT 1493.4000 1892.7800 1495.0000 1893.2600 ;
        RECT 1493.4000 1898.2200 1495.0000 1898.7000 ;
        RECT 1483.6600 1887.3400 1485.2600 1887.8200 ;
        RECT 1483.6600 1892.7800 1485.2600 1893.2600 ;
        RECT 1483.6600 1898.2200 1485.2600 1898.7000 ;
        RECT 1493.4000 1876.4600 1495.0000 1876.9400 ;
        RECT 1493.4000 1881.9000 1495.0000 1882.3800 ;
        RECT 1483.6600 1876.4600 1485.2600 1876.9400 ;
        RECT 1483.6600 1881.9000 1485.2600 1882.3800 ;
        RECT 1493.4000 1860.1400 1495.0000 1860.6200 ;
        RECT 1493.4000 1865.5800 1495.0000 1866.0600 ;
        RECT 1493.4000 1871.0200 1495.0000 1871.5000 ;
        RECT 1483.6600 1860.1400 1485.2600 1860.6200 ;
        RECT 1483.6600 1865.5800 1485.2600 1866.0600 ;
        RECT 1483.6600 1871.0200 1485.2600 1871.5000 ;
        RECT 1493.4000 1849.2600 1495.0000 1849.7400 ;
        RECT 1493.4000 1854.7000 1495.0000 1855.1800 ;
        RECT 1483.6600 1849.2600 1485.2600 1849.7400 ;
        RECT 1483.6600 1854.7000 1485.2600 1855.1800 ;
        RECT 1438.6600 1887.3400 1440.2600 1887.8200 ;
        RECT 1438.6600 1892.7800 1440.2600 1893.2600 ;
        RECT 1438.6600 1898.2200 1440.2600 1898.7000 ;
        RECT 1438.6600 1876.4600 1440.2600 1876.9400 ;
        RECT 1438.6600 1881.9000 1440.2600 1882.3800 ;
        RECT 1438.6600 1860.1400 1440.2600 1860.6200 ;
        RECT 1438.6600 1865.5800 1440.2600 1866.0600 ;
        RECT 1438.6600 1871.0200 1440.2600 1871.5000 ;
        RECT 1438.6600 1849.2600 1440.2600 1849.7400 ;
        RECT 1438.6600 1854.7000 1440.2600 1855.1800 ;
        RECT 1493.4000 1832.9400 1495.0000 1833.4200 ;
        RECT 1493.4000 1838.3800 1495.0000 1838.8600 ;
        RECT 1493.4000 1843.8200 1495.0000 1844.3000 ;
        RECT 1483.6600 1832.9400 1485.2600 1833.4200 ;
        RECT 1483.6600 1838.3800 1485.2600 1838.8600 ;
        RECT 1483.6600 1843.8200 1485.2600 1844.3000 ;
        RECT 1493.4000 1822.0600 1495.0000 1822.5400 ;
        RECT 1493.4000 1827.5000 1495.0000 1827.9800 ;
        RECT 1483.6600 1822.0600 1485.2600 1822.5400 ;
        RECT 1483.6600 1827.5000 1485.2600 1827.9800 ;
        RECT 1493.4000 1805.7400 1495.0000 1806.2200 ;
        RECT 1493.4000 1811.1800 1495.0000 1811.6600 ;
        RECT 1493.4000 1816.6200 1495.0000 1817.1000 ;
        RECT 1483.6600 1805.7400 1485.2600 1806.2200 ;
        RECT 1483.6600 1811.1800 1485.2600 1811.6600 ;
        RECT 1483.6600 1816.6200 1485.2600 1817.1000 ;
        RECT 1483.6600 1800.3000 1485.2600 1800.7800 ;
        RECT 1493.4000 1800.3000 1495.0000 1800.7800 ;
        RECT 1438.6600 1832.9400 1440.2600 1833.4200 ;
        RECT 1438.6600 1838.3800 1440.2600 1838.8600 ;
        RECT 1438.6600 1843.8200 1440.2600 1844.3000 ;
        RECT 1438.6600 1822.0600 1440.2600 1822.5400 ;
        RECT 1438.6600 1827.5000 1440.2600 1827.9800 ;
        RECT 1438.6600 1805.7400 1440.2600 1806.2200 ;
        RECT 1438.6600 1811.1800 1440.2600 1811.6600 ;
        RECT 1438.6600 1816.6200 1440.2600 1817.1000 ;
        RECT 1438.6600 1800.3000 1440.2600 1800.7800 ;
        RECT 1393.6600 1887.3400 1395.2600 1887.8200 ;
        RECT 1393.6600 1892.7800 1395.2600 1893.2600 ;
        RECT 1393.6600 1898.2200 1395.2600 1898.7000 ;
        RECT 1393.6600 1876.4600 1395.2600 1876.9400 ;
        RECT 1393.6600 1881.9000 1395.2600 1882.3800 ;
        RECT 1348.6600 1887.3400 1350.2600 1887.8200 ;
        RECT 1348.6600 1892.7800 1350.2600 1893.2600 ;
        RECT 1348.6600 1898.2200 1350.2600 1898.7000 ;
        RECT 1348.6600 1876.4600 1350.2600 1876.9400 ;
        RECT 1348.6600 1881.9000 1350.2600 1882.3800 ;
        RECT 1393.6600 1860.1400 1395.2600 1860.6200 ;
        RECT 1393.6600 1865.5800 1395.2600 1866.0600 ;
        RECT 1393.6600 1871.0200 1395.2600 1871.5000 ;
        RECT 1393.6600 1849.2600 1395.2600 1849.7400 ;
        RECT 1393.6600 1854.7000 1395.2600 1855.1800 ;
        RECT 1348.6600 1860.1400 1350.2600 1860.6200 ;
        RECT 1348.6600 1865.5800 1350.2600 1866.0600 ;
        RECT 1348.6600 1871.0200 1350.2600 1871.5000 ;
        RECT 1348.6600 1849.2600 1350.2600 1849.7400 ;
        RECT 1348.6600 1854.7000 1350.2600 1855.1800 ;
        RECT 1303.6600 1887.3400 1305.2600 1887.8200 ;
        RECT 1303.6600 1892.7800 1305.2600 1893.2600 ;
        RECT 1303.6600 1898.2200 1305.2600 1898.7000 ;
        RECT 1295.9000 1887.3400 1297.5000 1887.8200 ;
        RECT 1295.9000 1892.7800 1297.5000 1893.2600 ;
        RECT 1295.9000 1898.2200 1297.5000 1898.7000 ;
        RECT 1303.6600 1876.4600 1305.2600 1876.9400 ;
        RECT 1303.6600 1881.9000 1305.2600 1882.3800 ;
        RECT 1295.9000 1876.4600 1297.5000 1876.9400 ;
        RECT 1295.9000 1881.9000 1297.5000 1882.3800 ;
        RECT 1303.6600 1860.1400 1305.2600 1860.6200 ;
        RECT 1303.6600 1865.5800 1305.2600 1866.0600 ;
        RECT 1303.6600 1871.0200 1305.2600 1871.5000 ;
        RECT 1295.9000 1860.1400 1297.5000 1860.6200 ;
        RECT 1295.9000 1865.5800 1297.5000 1866.0600 ;
        RECT 1295.9000 1871.0200 1297.5000 1871.5000 ;
        RECT 1303.6600 1849.2600 1305.2600 1849.7400 ;
        RECT 1303.6600 1854.7000 1305.2600 1855.1800 ;
        RECT 1295.9000 1849.2600 1297.5000 1849.7400 ;
        RECT 1295.9000 1854.7000 1297.5000 1855.1800 ;
        RECT 1393.6600 1832.9400 1395.2600 1833.4200 ;
        RECT 1393.6600 1838.3800 1395.2600 1838.8600 ;
        RECT 1393.6600 1843.8200 1395.2600 1844.3000 ;
        RECT 1393.6600 1822.0600 1395.2600 1822.5400 ;
        RECT 1393.6600 1827.5000 1395.2600 1827.9800 ;
        RECT 1348.6600 1832.9400 1350.2600 1833.4200 ;
        RECT 1348.6600 1838.3800 1350.2600 1838.8600 ;
        RECT 1348.6600 1843.8200 1350.2600 1844.3000 ;
        RECT 1348.6600 1822.0600 1350.2600 1822.5400 ;
        RECT 1348.6600 1827.5000 1350.2600 1827.9800 ;
        RECT 1393.6600 1805.7400 1395.2600 1806.2200 ;
        RECT 1393.6600 1811.1800 1395.2600 1811.6600 ;
        RECT 1393.6600 1816.6200 1395.2600 1817.1000 ;
        RECT 1393.6600 1800.3000 1395.2600 1800.7800 ;
        RECT 1348.6600 1805.7400 1350.2600 1806.2200 ;
        RECT 1348.6600 1811.1800 1350.2600 1811.6600 ;
        RECT 1348.6600 1816.6200 1350.2600 1817.1000 ;
        RECT 1348.6600 1800.3000 1350.2600 1800.7800 ;
        RECT 1303.6600 1832.9400 1305.2600 1833.4200 ;
        RECT 1303.6600 1838.3800 1305.2600 1838.8600 ;
        RECT 1303.6600 1843.8200 1305.2600 1844.3000 ;
        RECT 1295.9000 1832.9400 1297.5000 1833.4200 ;
        RECT 1295.9000 1838.3800 1297.5000 1838.8600 ;
        RECT 1295.9000 1843.8200 1297.5000 1844.3000 ;
        RECT 1303.6600 1822.0600 1305.2600 1822.5400 ;
        RECT 1303.6600 1827.5000 1305.2600 1827.9800 ;
        RECT 1295.9000 1822.0600 1297.5000 1822.5400 ;
        RECT 1295.9000 1827.5000 1297.5000 1827.9800 ;
        RECT 1303.6600 1805.7400 1305.2600 1806.2200 ;
        RECT 1303.6600 1811.1800 1305.2600 1811.6600 ;
        RECT 1303.6600 1816.6200 1305.2600 1817.1000 ;
        RECT 1295.9000 1805.7400 1297.5000 1806.2200 ;
        RECT 1295.9000 1811.1800 1297.5000 1811.6600 ;
        RECT 1295.9000 1816.6200 1297.5000 1817.1000 ;
        RECT 1295.9000 1800.3000 1297.5000 1800.7800 ;
        RECT 1303.6600 1800.3000 1305.2600 1800.7800 ;
        RECT 1290.3400 2002.6100 1500.5600 2004.2100 ;
        RECT 1290.3400 1796.1100 1500.5600 1797.7100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1790.6800 1297.5000 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 2008.7200 1297.5000 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1790.6800 1495.0000 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 2008.7200 1495.0000 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1796.1100 1291.9400 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1796.1100 1500.5600 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 2002.6100 1291.9400 2004.2100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 2002.6100 1500.5600 2004.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 1566.4700 1485.2600 1774.5700 ;
        RECT 1438.6600 1566.4700 1440.2600 1774.5700 ;
        RECT 1393.6600 1566.4700 1395.2600 1774.5700 ;
        RECT 1348.6600 1566.4700 1350.2600 1774.5700 ;
        RECT 1303.6600 1566.4700 1305.2600 1774.5700 ;
        RECT 1493.4000 1561.0400 1495.0000 1780.6800 ;
        RECT 1295.9000 1561.0400 1297.5000 1780.6800 ;
      LAYER met3 ;
        RECT 1493.4000 1755.6200 1495.0000 1756.1000 ;
        RECT 1493.4000 1761.0600 1495.0000 1761.5400 ;
        RECT 1483.6600 1755.6200 1485.2600 1756.1000 ;
        RECT 1483.6600 1761.0600 1485.2600 1761.5400 ;
        RECT 1483.6600 1766.5000 1485.2600 1766.9800 ;
        RECT 1493.4000 1766.5000 1495.0000 1766.9800 ;
        RECT 1493.4000 1744.7400 1495.0000 1745.2200 ;
        RECT 1493.4000 1750.1800 1495.0000 1750.6600 ;
        RECT 1483.6600 1744.7400 1485.2600 1745.2200 ;
        RECT 1483.6600 1750.1800 1485.2600 1750.6600 ;
        RECT 1493.4000 1728.4200 1495.0000 1728.9000 ;
        RECT 1493.4000 1733.8600 1495.0000 1734.3400 ;
        RECT 1483.6600 1728.4200 1485.2600 1728.9000 ;
        RECT 1483.6600 1733.8600 1485.2600 1734.3400 ;
        RECT 1483.6600 1739.3000 1485.2600 1739.7800 ;
        RECT 1493.4000 1739.3000 1495.0000 1739.7800 ;
        RECT 1438.6600 1755.6200 1440.2600 1756.1000 ;
        RECT 1438.6600 1761.0600 1440.2600 1761.5400 ;
        RECT 1438.6600 1766.5000 1440.2600 1766.9800 ;
        RECT 1438.6600 1744.7400 1440.2600 1745.2200 ;
        RECT 1438.6600 1750.1800 1440.2600 1750.6600 ;
        RECT 1438.6600 1728.4200 1440.2600 1728.9000 ;
        RECT 1438.6600 1733.8600 1440.2600 1734.3400 ;
        RECT 1438.6600 1739.3000 1440.2600 1739.7800 ;
        RECT 1493.4000 1712.1000 1495.0000 1712.5800 ;
        RECT 1493.4000 1717.5400 1495.0000 1718.0200 ;
        RECT 1493.4000 1722.9800 1495.0000 1723.4600 ;
        RECT 1483.6600 1712.1000 1485.2600 1712.5800 ;
        RECT 1483.6600 1717.5400 1485.2600 1718.0200 ;
        RECT 1483.6600 1722.9800 1485.2600 1723.4600 ;
        RECT 1493.4000 1701.2200 1495.0000 1701.7000 ;
        RECT 1493.4000 1706.6600 1495.0000 1707.1400 ;
        RECT 1483.6600 1701.2200 1485.2600 1701.7000 ;
        RECT 1483.6600 1706.6600 1485.2600 1707.1400 ;
        RECT 1493.4000 1684.9000 1495.0000 1685.3800 ;
        RECT 1493.4000 1690.3400 1495.0000 1690.8200 ;
        RECT 1493.4000 1695.7800 1495.0000 1696.2600 ;
        RECT 1483.6600 1684.9000 1485.2600 1685.3800 ;
        RECT 1483.6600 1690.3400 1485.2600 1690.8200 ;
        RECT 1483.6600 1695.7800 1485.2600 1696.2600 ;
        RECT 1493.4000 1674.0200 1495.0000 1674.5000 ;
        RECT 1493.4000 1679.4600 1495.0000 1679.9400 ;
        RECT 1483.6600 1674.0200 1485.2600 1674.5000 ;
        RECT 1483.6600 1679.4600 1485.2600 1679.9400 ;
        RECT 1438.6600 1712.1000 1440.2600 1712.5800 ;
        RECT 1438.6600 1717.5400 1440.2600 1718.0200 ;
        RECT 1438.6600 1722.9800 1440.2600 1723.4600 ;
        RECT 1438.6600 1701.2200 1440.2600 1701.7000 ;
        RECT 1438.6600 1706.6600 1440.2600 1707.1400 ;
        RECT 1438.6600 1684.9000 1440.2600 1685.3800 ;
        RECT 1438.6600 1690.3400 1440.2600 1690.8200 ;
        RECT 1438.6600 1695.7800 1440.2600 1696.2600 ;
        RECT 1438.6600 1674.0200 1440.2600 1674.5000 ;
        RECT 1438.6600 1679.4600 1440.2600 1679.9400 ;
        RECT 1393.6600 1755.6200 1395.2600 1756.1000 ;
        RECT 1393.6600 1761.0600 1395.2600 1761.5400 ;
        RECT 1393.6600 1766.5000 1395.2600 1766.9800 ;
        RECT 1348.6600 1755.6200 1350.2600 1756.1000 ;
        RECT 1348.6600 1761.0600 1350.2600 1761.5400 ;
        RECT 1348.6600 1766.5000 1350.2600 1766.9800 ;
        RECT 1393.6600 1744.7400 1395.2600 1745.2200 ;
        RECT 1393.6600 1750.1800 1395.2600 1750.6600 ;
        RECT 1393.6600 1728.4200 1395.2600 1728.9000 ;
        RECT 1393.6600 1733.8600 1395.2600 1734.3400 ;
        RECT 1393.6600 1739.3000 1395.2600 1739.7800 ;
        RECT 1348.6600 1744.7400 1350.2600 1745.2200 ;
        RECT 1348.6600 1750.1800 1350.2600 1750.6600 ;
        RECT 1348.6600 1728.4200 1350.2600 1728.9000 ;
        RECT 1348.6600 1733.8600 1350.2600 1734.3400 ;
        RECT 1348.6600 1739.3000 1350.2600 1739.7800 ;
        RECT 1303.6600 1755.6200 1305.2600 1756.1000 ;
        RECT 1303.6600 1761.0600 1305.2600 1761.5400 ;
        RECT 1295.9000 1755.6200 1297.5000 1756.1000 ;
        RECT 1295.9000 1761.0600 1297.5000 1761.5400 ;
        RECT 1295.9000 1766.5000 1297.5000 1766.9800 ;
        RECT 1303.6600 1766.5000 1305.2600 1766.9800 ;
        RECT 1303.6600 1744.7400 1305.2600 1745.2200 ;
        RECT 1303.6600 1750.1800 1305.2600 1750.6600 ;
        RECT 1295.9000 1744.7400 1297.5000 1745.2200 ;
        RECT 1295.9000 1750.1800 1297.5000 1750.6600 ;
        RECT 1303.6600 1728.4200 1305.2600 1728.9000 ;
        RECT 1303.6600 1733.8600 1305.2600 1734.3400 ;
        RECT 1295.9000 1728.4200 1297.5000 1728.9000 ;
        RECT 1295.9000 1733.8600 1297.5000 1734.3400 ;
        RECT 1295.9000 1739.3000 1297.5000 1739.7800 ;
        RECT 1303.6600 1739.3000 1305.2600 1739.7800 ;
        RECT 1393.6600 1712.1000 1395.2600 1712.5800 ;
        RECT 1393.6600 1717.5400 1395.2600 1718.0200 ;
        RECT 1393.6600 1722.9800 1395.2600 1723.4600 ;
        RECT 1393.6600 1701.2200 1395.2600 1701.7000 ;
        RECT 1393.6600 1706.6600 1395.2600 1707.1400 ;
        RECT 1348.6600 1712.1000 1350.2600 1712.5800 ;
        RECT 1348.6600 1717.5400 1350.2600 1718.0200 ;
        RECT 1348.6600 1722.9800 1350.2600 1723.4600 ;
        RECT 1348.6600 1701.2200 1350.2600 1701.7000 ;
        RECT 1348.6600 1706.6600 1350.2600 1707.1400 ;
        RECT 1393.6600 1684.9000 1395.2600 1685.3800 ;
        RECT 1393.6600 1690.3400 1395.2600 1690.8200 ;
        RECT 1393.6600 1695.7800 1395.2600 1696.2600 ;
        RECT 1393.6600 1674.0200 1395.2600 1674.5000 ;
        RECT 1393.6600 1679.4600 1395.2600 1679.9400 ;
        RECT 1348.6600 1684.9000 1350.2600 1685.3800 ;
        RECT 1348.6600 1690.3400 1350.2600 1690.8200 ;
        RECT 1348.6600 1695.7800 1350.2600 1696.2600 ;
        RECT 1348.6600 1674.0200 1350.2600 1674.5000 ;
        RECT 1348.6600 1679.4600 1350.2600 1679.9400 ;
        RECT 1303.6600 1712.1000 1305.2600 1712.5800 ;
        RECT 1303.6600 1717.5400 1305.2600 1718.0200 ;
        RECT 1303.6600 1722.9800 1305.2600 1723.4600 ;
        RECT 1295.9000 1712.1000 1297.5000 1712.5800 ;
        RECT 1295.9000 1717.5400 1297.5000 1718.0200 ;
        RECT 1295.9000 1722.9800 1297.5000 1723.4600 ;
        RECT 1303.6600 1701.2200 1305.2600 1701.7000 ;
        RECT 1303.6600 1706.6600 1305.2600 1707.1400 ;
        RECT 1295.9000 1701.2200 1297.5000 1701.7000 ;
        RECT 1295.9000 1706.6600 1297.5000 1707.1400 ;
        RECT 1303.6600 1684.9000 1305.2600 1685.3800 ;
        RECT 1303.6600 1690.3400 1305.2600 1690.8200 ;
        RECT 1303.6600 1695.7800 1305.2600 1696.2600 ;
        RECT 1295.9000 1684.9000 1297.5000 1685.3800 ;
        RECT 1295.9000 1690.3400 1297.5000 1690.8200 ;
        RECT 1295.9000 1695.7800 1297.5000 1696.2600 ;
        RECT 1303.6600 1674.0200 1305.2600 1674.5000 ;
        RECT 1303.6600 1679.4600 1305.2600 1679.9400 ;
        RECT 1295.9000 1674.0200 1297.5000 1674.5000 ;
        RECT 1295.9000 1679.4600 1297.5000 1679.9400 ;
        RECT 1493.4000 1657.7000 1495.0000 1658.1800 ;
        RECT 1493.4000 1663.1400 1495.0000 1663.6200 ;
        RECT 1493.4000 1668.5800 1495.0000 1669.0600 ;
        RECT 1483.6600 1657.7000 1485.2600 1658.1800 ;
        RECT 1483.6600 1663.1400 1485.2600 1663.6200 ;
        RECT 1483.6600 1668.5800 1485.2600 1669.0600 ;
        RECT 1493.4000 1646.8200 1495.0000 1647.3000 ;
        RECT 1493.4000 1652.2600 1495.0000 1652.7400 ;
        RECT 1483.6600 1646.8200 1485.2600 1647.3000 ;
        RECT 1483.6600 1652.2600 1485.2600 1652.7400 ;
        RECT 1493.4000 1630.5000 1495.0000 1630.9800 ;
        RECT 1493.4000 1635.9400 1495.0000 1636.4200 ;
        RECT 1493.4000 1641.3800 1495.0000 1641.8600 ;
        RECT 1483.6600 1630.5000 1485.2600 1630.9800 ;
        RECT 1483.6600 1635.9400 1485.2600 1636.4200 ;
        RECT 1483.6600 1641.3800 1485.2600 1641.8600 ;
        RECT 1493.4000 1619.6200 1495.0000 1620.1000 ;
        RECT 1493.4000 1625.0600 1495.0000 1625.5400 ;
        RECT 1483.6600 1619.6200 1485.2600 1620.1000 ;
        RECT 1483.6600 1625.0600 1485.2600 1625.5400 ;
        RECT 1438.6600 1657.7000 1440.2600 1658.1800 ;
        RECT 1438.6600 1663.1400 1440.2600 1663.6200 ;
        RECT 1438.6600 1668.5800 1440.2600 1669.0600 ;
        RECT 1438.6600 1646.8200 1440.2600 1647.3000 ;
        RECT 1438.6600 1652.2600 1440.2600 1652.7400 ;
        RECT 1438.6600 1630.5000 1440.2600 1630.9800 ;
        RECT 1438.6600 1635.9400 1440.2600 1636.4200 ;
        RECT 1438.6600 1641.3800 1440.2600 1641.8600 ;
        RECT 1438.6600 1619.6200 1440.2600 1620.1000 ;
        RECT 1438.6600 1625.0600 1440.2600 1625.5400 ;
        RECT 1493.4000 1603.3000 1495.0000 1603.7800 ;
        RECT 1493.4000 1608.7400 1495.0000 1609.2200 ;
        RECT 1493.4000 1614.1800 1495.0000 1614.6600 ;
        RECT 1483.6600 1603.3000 1485.2600 1603.7800 ;
        RECT 1483.6600 1608.7400 1485.2600 1609.2200 ;
        RECT 1483.6600 1614.1800 1485.2600 1614.6600 ;
        RECT 1493.4000 1592.4200 1495.0000 1592.9000 ;
        RECT 1493.4000 1597.8600 1495.0000 1598.3400 ;
        RECT 1483.6600 1592.4200 1485.2600 1592.9000 ;
        RECT 1483.6600 1597.8600 1485.2600 1598.3400 ;
        RECT 1493.4000 1576.1000 1495.0000 1576.5800 ;
        RECT 1493.4000 1581.5400 1495.0000 1582.0200 ;
        RECT 1493.4000 1586.9800 1495.0000 1587.4600 ;
        RECT 1483.6600 1576.1000 1485.2600 1576.5800 ;
        RECT 1483.6600 1581.5400 1485.2600 1582.0200 ;
        RECT 1483.6600 1586.9800 1485.2600 1587.4600 ;
        RECT 1483.6600 1570.6600 1485.2600 1571.1400 ;
        RECT 1493.4000 1570.6600 1495.0000 1571.1400 ;
        RECT 1438.6600 1603.3000 1440.2600 1603.7800 ;
        RECT 1438.6600 1608.7400 1440.2600 1609.2200 ;
        RECT 1438.6600 1614.1800 1440.2600 1614.6600 ;
        RECT 1438.6600 1592.4200 1440.2600 1592.9000 ;
        RECT 1438.6600 1597.8600 1440.2600 1598.3400 ;
        RECT 1438.6600 1576.1000 1440.2600 1576.5800 ;
        RECT 1438.6600 1581.5400 1440.2600 1582.0200 ;
        RECT 1438.6600 1586.9800 1440.2600 1587.4600 ;
        RECT 1438.6600 1570.6600 1440.2600 1571.1400 ;
        RECT 1393.6600 1657.7000 1395.2600 1658.1800 ;
        RECT 1393.6600 1663.1400 1395.2600 1663.6200 ;
        RECT 1393.6600 1668.5800 1395.2600 1669.0600 ;
        RECT 1393.6600 1646.8200 1395.2600 1647.3000 ;
        RECT 1393.6600 1652.2600 1395.2600 1652.7400 ;
        RECT 1348.6600 1657.7000 1350.2600 1658.1800 ;
        RECT 1348.6600 1663.1400 1350.2600 1663.6200 ;
        RECT 1348.6600 1668.5800 1350.2600 1669.0600 ;
        RECT 1348.6600 1646.8200 1350.2600 1647.3000 ;
        RECT 1348.6600 1652.2600 1350.2600 1652.7400 ;
        RECT 1393.6600 1630.5000 1395.2600 1630.9800 ;
        RECT 1393.6600 1635.9400 1395.2600 1636.4200 ;
        RECT 1393.6600 1641.3800 1395.2600 1641.8600 ;
        RECT 1393.6600 1619.6200 1395.2600 1620.1000 ;
        RECT 1393.6600 1625.0600 1395.2600 1625.5400 ;
        RECT 1348.6600 1630.5000 1350.2600 1630.9800 ;
        RECT 1348.6600 1635.9400 1350.2600 1636.4200 ;
        RECT 1348.6600 1641.3800 1350.2600 1641.8600 ;
        RECT 1348.6600 1619.6200 1350.2600 1620.1000 ;
        RECT 1348.6600 1625.0600 1350.2600 1625.5400 ;
        RECT 1303.6600 1657.7000 1305.2600 1658.1800 ;
        RECT 1303.6600 1663.1400 1305.2600 1663.6200 ;
        RECT 1303.6600 1668.5800 1305.2600 1669.0600 ;
        RECT 1295.9000 1657.7000 1297.5000 1658.1800 ;
        RECT 1295.9000 1663.1400 1297.5000 1663.6200 ;
        RECT 1295.9000 1668.5800 1297.5000 1669.0600 ;
        RECT 1303.6600 1646.8200 1305.2600 1647.3000 ;
        RECT 1303.6600 1652.2600 1305.2600 1652.7400 ;
        RECT 1295.9000 1646.8200 1297.5000 1647.3000 ;
        RECT 1295.9000 1652.2600 1297.5000 1652.7400 ;
        RECT 1303.6600 1630.5000 1305.2600 1630.9800 ;
        RECT 1303.6600 1635.9400 1305.2600 1636.4200 ;
        RECT 1303.6600 1641.3800 1305.2600 1641.8600 ;
        RECT 1295.9000 1630.5000 1297.5000 1630.9800 ;
        RECT 1295.9000 1635.9400 1297.5000 1636.4200 ;
        RECT 1295.9000 1641.3800 1297.5000 1641.8600 ;
        RECT 1303.6600 1619.6200 1305.2600 1620.1000 ;
        RECT 1303.6600 1625.0600 1305.2600 1625.5400 ;
        RECT 1295.9000 1619.6200 1297.5000 1620.1000 ;
        RECT 1295.9000 1625.0600 1297.5000 1625.5400 ;
        RECT 1393.6600 1603.3000 1395.2600 1603.7800 ;
        RECT 1393.6600 1608.7400 1395.2600 1609.2200 ;
        RECT 1393.6600 1614.1800 1395.2600 1614.6600 ;
        RECT 1393.6600 1592.4200 1395.2600 1592.9000 ;
        RECT 1393.6600 1597.8600 1395.2600 1598.3400 ;
        RECT 1348.6600 1603.3000 1350.2600 1603.7800 ;
        RECT 1348.6600 1608.7400 1350.2600 1609.2200 ;
        RECT 1348.6600 1614.1800 1350.2600 1614.6600 ;
        RECT 1348.6600 1592.4200 1350.2600 1592.9000 ;
        RECT 1348.6600 1597.8600 1350.2600 1598.3400 ;
        RECT 1393.6600 1576.1000 1395.2600 1576.5800 ;
        RECT 1393.6600 1581.5400 1395.2600 1582.0200 ;
        RECT 1393.6600 1586.9800 1395.2600 1587.4600 ;
        RECT 1393.6600 1570.6600 1395.2600 1571.1400 ;
        RECT 1348.6600 1576.1000 1350.2600 1576.5800 ;
        RECT 1348.6600 1581.5400 1350.2600 1582.0200 ;
        RECT 1348.6600 1586.9800 1350.2600 1587.4600 ;
        RECT 1348.6600 1570.6600 1350.2600 1571.1400 ;
        RECT 1303.6600 1603.3000 1305.2600 1603.7800 ;
        RECT 1303.6600 1608.7400 1305.2600 1609.2200 ;
        RECT 1303.6600 1614.1800 1305.2600 1614.6600 ;
        RECT 1295.9000 1603.3000 1297.5000 1603.7800 ;
        RECT 1295.9000 1608.7400 1297.5000 1609.2200 ;
        RECT 1295.9000 1614.1800 1297.5000 1614.6600 ;
        RECT 1303.6600 1592.4200 1305.2600 1592.9000 ;
        RECT 1303.6600 1597.8600 1305.2600 1598.3400 ;
        RECT 1295.9000 1592.4200 1297.5000 1592.9000 ;
        RECT 1295.9000 1597.8600 1297.5000 1598.3400 ;
        RECT 1303.6600 1576.1000 1305.2600 1576.5800 ;
        RECT 1303.6600 1581.5400 1305.2600 1582.0200 ;
        RECT 1303.6600 1586.9800 1305.2600 1587.4600 ;
        RECT 1295.9000 1576.1000 1297.5000 1576.5800 ;
        RECT 1295.9000 1581.5400 1297.5000 1582.0200 ;
        RECT 1295.9000 1586.9800 1297.5000 1587.4600 ;
        RECT 1295.9000 1570.6600 1297.5000 1571.1400 ;
        RECT 1303.6600 1570.6600 1305.2600 1571.1400 ;
        RECT 1290.3400 1772.9700 1500.5600 1774.5700 ;
        RECT 1290.3400 1566.4700 1500.5600 1568.0700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1561.0400 1297.5000 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1779.0800 1297.5000 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1561.0400 1495.0000 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1779.0800 1495.0000 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1566.4700 1291.9400 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1566.4700 1500.5600 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1772.9700 1291.9400 1774.5700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1772.9700 1500.5600 1774.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 1336.8300 1485.2600 1544.9300 ;
        RECT 1438.6600 1336.8300 1440.2600 1544.9300 ;
        RECT 1393.6600 1336.8300 1395.2600 1544.9300 ;
        RECT 1348.6600 1336.8300 1350.2600 1544.9300 ;
        RECT 1303.6600 1336.8300 1305.2600 1544.9300 ;
        RECT 1493.4000 1331.4000 1495.0000 1551.0400 ;
        RECT 1295.9000 1331.4000 1297.5000 1551.0400 ;
      LAYER met3 ;
        RECT 1493.4000 1525.9800 1495.0000 1526.4600 ;
        RECT 1493.4000 1531.4200 1495.0000 1531.9000 ;
        RECT 1483.6600 1525.9800 1485.2600 1526.4600 ;
        RECT 1483.6600 1531.4200 1485.2600 1531.9000 ;
        RECT 1483.6600 1536.8600 1485.2600 1537.3400 ;
        RECT 1493.4000 1536.8600 1495.0000 1537.3400 ;
        RECT 1493.4000 1515.1000 1495.0000 1515.5800 ;
        RECT 1493.4000 1520.5400 1495.0000 1521.0200 ;
        RECT 1483.6600 1515.1000 1485.2600 1515.5800 ;
        RECT 1483.6600 1520.5400 1485.2600 1521.0200 ;
        RECT 1493.4000 1498.7800 1495.0000 1499.2600 ;
        RECT 1493.4000 1504.2200 1495.0000 1504.7000 ;
        RECT 1483.6600 1498.7800 1485.2600 1499.2600 ;
        RECT 1483.6600 1504.2200 1485.2600 1504.7000 ;
        RECT 1483.6600 1509.6600 1485.2600 1510.1400 ;
        RECT 1493.4000 1509.6600 1495.0000 1510.1400 ;
        RECT 1438.6600 1525.9800 1440.2600 1526.4600 ;
        RECT 1438.6600 1531.4200 1440.2600 1531.9000 ;
        RECT 1438.6600 1536.8600 1440.2600 1537.3400 ;
        RECT 1438.6600 1515.1000 1440.2600 1515.5800 ;
        RECT 1438.6600 1520.5400 1440.2600 1521.0200 ;
        RECT 1438.6600 1498.7800 1440.2600 1499.2600 ;
        RECT 1438.6600 1504.2200 1440.2600 1504.7000 ;
        RECT 1438.6600 1509.6600 1440.2600 1510.1400 ;
        RECT 1493.4000 1482.4600 1495.0000 1482.9400 ;
        RECT 1493.4000 1487.9000 1495.0000 1488.3800 ;
        RECT 1493.4000 1493.3400 1495.0000 1493.8200 ;
        RECT 1483.6600 1482.4600 1485.2600 1482.9400 ;
        RECT 1483.6600 1487.9000 1485.2600 1488.3800 ;
        RECT 1483.6600 1493.3400 1485.2600 1493.8200 ;
        RECT 1493.4000 1471.5800 1495.0000 1472.0600 ;
        RECT 1493.4000 1477.0200 1495.0000 1477.5000 ;
        RECT 1483.6600 1471.5800 1485.2600 1472.0600 ;
        RECT 1483.6600 1477.0200 1485.2600 1477.5000 ;
        RECT 1493.4000 1455.2600 1495.0000 1455.7400 ;
        RECT 1493.4000 1460.7000 1495.0000 1461.1800 ;
        RECT 1493.4000 1466.1400 1495.0000 1466.6200 ;
        RECT 1483.6600 1455.2600 1485.2600 1455.7400 ;
        RECT 1483.6600 1460.7000 1485.2600 1461.1800 ;
        RECT 1483.6600 1466.1400 1485.2600 1466.6200 ;
        RECT 1493.4000 1444.3800 1495.0000 1444.8600 ;
        RECT 1493.4000 1449.8200 1495.0000 1450.3000 ;
        RECT 1483.6600 1444.3800 1485.2600 1444.8600 ;
        RECT 1483.6600 1449.8200 1485.2600 1450.3000 ;
        RECT 1438.6600 1482.4600 1440.2600 1482.9400 ;
        RECT 1438.6600 1487.9000 1440.2600 1488.3800 ;
        RECT 1438.6600 1493.3400 1440.2600 1493.8200 ;
        RECT 1438.6600 1471.5800 1440.2600 1472.0600 ;
        RECT 1438.6600 1477.0200 1440.2600 1477.5000 ;
        RECT 1438.6600 1455.2600 1440.2600 1455.7400 ;
        RECT 1438.6600 1460.7000 1440.2600 1461.1800 ;
        RECT 1438.6600 1466.1400 1440.2600 1466.6200 ;
        RECT 1438.6600 1444.3800 1440.2600 1444.8600 ;
        RECT 1438.6600 1449.8200 1440.2600 1450.3000 ;
        RECT 1393.6600 1525.9800 1395.2600 1526.4600 ;
        RECT 1393.6600 1531.4200 1395.2600 1531.9000 ;
        RECT 1393.6600 1536.8600 1395.2600 1537.3400 ;
        RECT 1348.6600 1525.9800 1350.2600 1526.4600 ;
        RECT 1348.6600 1531.4200 1350.2600 1531.9000 ;
        RECT 1348.6600 1536.8600 1350.2600 1537.3400 ;
        RECT 1393.6600 1515.1000 1395.2600 1515.5800 ;
        RECT 1393.6600 1520.5400 1395.2600 1521.0200 ;
        RECT 1393.6600 1498.7800 1395.2600 1499.2600 ;
        RECT 1393.6600 1504.2200 1395.2600 1504.7000 ;
        RECT 1393.6600 1509.6600 1395.2600 1510.1400 ;
        RECT 1348.6600 1515.1000 1350.2600 1515.5800 ;
        RECT 1348.6600 1520.5400 1350.2600 1521.0200 ;
        RECT 1348.6600 1498.7800 1350.2600 1499.2600 ;
        RECT 1348.6600 1504.2200 1350.2600 1504.7000 ;
        RECT 1348.6600 1509.6600 1350.2600 1510.1400 ;
        RECT 1303.6600 1525.9800 1305.2600 1526.4600 ;
        RECT 1303.6600 1531.4200 1305.2600 1531.9000 ;
        RECT 1295.9000 1525.9800 1297.5000 1526.4600 ;
        RECT 1295.9000 1531.4200 1297.5000 1531.9000 ;
        RECT 1295.9000 1536.8600 1297.5000 1537.3400 ;
        RECT 1303.6600 1536.8600 1305.2600 1537.3400 ;
        RECT 1303.6600 1515.1000 1305.2600 1515.5800 ;
        RECT 1303.6600 1520.5400 1305.2600 1521.0200 ;
        RECT 1295.9000 1515.1000 1297.5000 1515.5800 ;
        RECT 1295.9000 1520.5400 1297.5000 1521.0200 ;
        RECT 1303.6600 1498.7800 1305.2600 1499.2600 ;
        RECT 1303.6600 1504.2200 1305.2600 1504.7000 ;
        RECT 1295.9000 1498.7800 1297.5000 1499.2600 ;
        RECT 1295.9000 1504.2200 1297.5000 1504.7000 ;
        RECT 1295.9000 1509.6600 1297.5000 1510.1400 ;
        RECT 1303.6600 1509.6600 1305.2600 1510.1400 ;
        RECT 1393.6600 1482.4600 1395.2600 1482.9400 ;
        RECT 1393.6600 1487.9000 1395.2600 1488.3800 ;
        RECT 1393.6600 1493.3400 1395.2600 1493.8200 ;
        RECT 1393.6600 1471.5800 1395.2600 1472.0600 ;
        RECT 1393.6600 1477.0200 1395.2600 1477.5000 ;
        RECT 1348.6600 1482.4600 1350.2600 1482.9400 ;
        RECT 1348.6600 1487.9000 1350.2600 1488.3800 ;
        RECT 1348.6600 1493.3400 1350.2600 1493.8200 ;
        RECT 1348.6600 1471.5800 1350.2600 1472.0600 ;
        RECT 1348.6600 1477.0200 1350.2600 1477.5000 ;
        RECT 1393.6600 1455.2600 1395.2600 1455.7400 ;
        RECT 1393.6600 1460.7000 1395.2600 1461.1800 ;
        RECT 1393.6600 1466.1400 1395.2600 1466.6200 ;
        RECT 1393.6600 1444.3800 1395.2600 1444.8600 ;
        RECT 1393.6600 1449.8200 1395.2600 1450.3000 ;
        RECT 1348.6600 1455.2600 1350.2600 1455.7400 ;
        RECT 1348.6600 1460.7000 1350.2600 1461.1800 ;
        RECT 1348.6600 1466.1400 1350.2600 1466.6200 ;
        RECT 1348.6600 1444.3800 1350.2600 1444.8600 ;
        RECT 1348.6600 1449.8200 1350.2600 1450.3000 ;
        RECT 1303.6600 1482.4600 1305.2600 1482.9400 ;
        RECT 1303.6600 1487.9000 1305.2600 1488.3800 ;
        RECT 1303.6600 1493.3400 1305.2600 1493.8200 ;
        RECT 1295.9000 1482.4600 1297.5000 1482.9400 ;
        RECT 1295.9000 1487.9000 1297.5000 1488.3800 ;
        RECT 1295.9000 1493.3400 1297.5000 1493.8200 ;
        RECT 1303.6600 1471.5800 1305.2600 1472.0600 ;
        RECT 1303.6600 1477.0200 1305.2600 1477.5000 ;
        RECT 1295.9000 1471.5800 1297.5000 1472.0600 ;
        RECT 1295.9000 1477.0200 1297.5000 1477.5000 ;
        RECT 1303.6600 1455.2600 1305.2600 1455.7400 ;
        RECT 1303.6600 1460.7000 1305.2600 1461.1800 ;
        RECT 1303.6600 1466.1400 1305.2600 1466.6200 ;
        RECT 1295.9000 1455.2600 1297.5000 1455.7400 ;
        RECT 1295.9000 1460.7000 1297.5000 1461.1800 ;
        RECT 1295.9000 1466.1400 1297.5000 1466.6200 ;
        RECT 1303.6600 1444.3800 1305.2600 1444.8600 ;
        RECT 1303.6600 1449.8200 1305.2600 1450.3000 ;
        RECT 1295.9000 1444.3800 1297.5000 1444.8600 ;
        RECT 1295.9000 1449.8200 1297.5000 1450.3000 ;
        RECT 1493.4000 1428.0600 1495.0000 1428.5400 ;
        RECT 1493.4000 1433.5000 1495.0000 1433.9800 ;
        RECT 1493.4000 1438.9400 1495.0000 1439.4200 ;
        RECT 1483.6600 1428.0600 1485.2600 1428.5400 ;
        RECT 1483.6600 1433.5000 1485.2600 1433.9800 ;
        RECT 1483.6600 1438.9400 1485.2600 1439.4200 ;
        RECT 1493.4000 1417.1800 1495.0000 1417.6600 ;
        RECT 1493.4000 1422.6200 1495.0000 1423.1000 ;
        RECT 1483.6600 1417.1800 1485.2600 1417.6600 ;
        RECT 1483.6600 1422.6200 1485.2600 1423.1000 ;
        RECT 1493.4000 1400.8600 1495.0000 1401.3400 ;
        RECT 1493.4000 1406.3000 1495.0000 1406.7800 ;
        RECT 1493.4000 1411.7400 1495.0000 1412.2200 ;
        RECT 1483.6600 1400.8600 1485.2600 1401.3400 ;
        RECT 1483.6600 1406.3000 1485.2600 1406.7800 ;
        RECT 1483.6600 1411.7400 1485.2600 1412.2200 ;
        RECT 1493.4000 1389.9800 1495.0000 1390.4600 ;
        RECT 1493.4000 1395.4200 1495.0000 1395.9000 ;
        RECT 1483.6600 1389.9800 1485.2600 1390.4600 ;
        RECT 1483.6600 1395.4200 1485.2600 1395.9000 ;
        RECT 1438.6600 1428.0600 1440.2600 1428.5400 ;
        RECT 1438.6600 1433.5000 1440.2600 1433.9800 ;
        RECT 1438.6600 1438.9400 1440.2600 1439.4200 ;
        RECT 1438.6600 1417.1800 1440.2600 1417.6600 ;
        RECT 1438.6600 1422.6200 1440.2600 1423.1000 ;
        RECT 1438.6600 1400.8600 1440.2600 1401.3400 ;
        RECT 1438.6600 1406.3000 1440.2600 1406.7800 ;
        RECT 1438.6600 1411.7400 1440.2600 1412.2200 ;
        RECT 1438.6600 1389.9800 1440.2600 1390.4600 ;
        RECT 1438.6600 1395.4200 1440.2600 1395.9000 ;
        RECT 1493.4000 1373.6600 1495.0000 1374.1400 ;
        RECT 1493.4000 1379.1000 1495.0000 1379.5800 ;
        RECT 1493.4000 1384.5400 1495.0000 1385.0200 ;
        RECT 1483.6600 1373.6600 1485.2600 1374.1400 ;
        RECT 1483.6600 1379.1000 1485.2600 1379.5800 ;
        RECT 1483.6600 1384.5400 1485.2600 1385.0200 ;
        RECT 1493.4000 1362.7800 1495.0000 1363.2600 ;
        RECT 1493.4000 1368.2200 1495.0000 1368.7000 ;
        RECT 1483.6600 1362.7800 1485.2600 1363.2600 ;
        RECT 1483.6600 1368.2200 1485.2600 1368.7000 ;
        RECT 1493.4000 1346.4600 1495.0000 1346.9400 ;
        RECT 1493.4000 1351.9000 1495.0000 1352.3800 ;
        RECT 1493.4000 1357.3400 1495.0000 1357.8200 ;
        RECT 1483.6600 1346.4600 1485.2600 1346.9400 ;
        RECT 1483.6600 1351.9000 1485.2600 1352.3800 ;
        RECT 1483.6600 1357.3400 1485.2600 1357.8200 ;
        RECT 1483.6600 1341.0200 1485.2600 1341.5000 ;
        RECT 1493.4000 1341.0200 1495.0000 1341.5000 ;
        RECT 1438.6600 1373.6600 1440.2600 1374.1400 ;
        RECT 1438.6600 1379.1000 1440.2600 1379.5800 ;
        RECT 1438.6600 1384.5400 1440.2600 1385.0200 ;
        RECT 1438.6600 1362.7800 1440.2600 1363.2600 ;
        RECT 1438.6600 1368.2200 1440.2600 1368.7000 ;
        RECT 1438.6600 1346.4600 1440.2600 1346.9400 ;
        RECT 1438.6600 1351.9000 1440.2600 1352.3800 ;
        RECT 1438.6600 1357.3400 1440.2600 1357.8200 ;
        RECT 1438.6600 1341.0200 1440.2600 1341.5000 ;
        RECT 1393.6600 1428.0600 1395.2600 1428.5400 ;
        RECT 1393.6600 1433.5000 1395.2600 1433.9800 ;
        RECT 1393.6600 1438.9400 1395.2600 1439.4200 ;
        RECT 1393.6600 1417.1800 1395.2600 1417.6600 ;
        RECT 1393.6600 1422.6200 1395.2600 1423.1000 ;
        RECT 1348.6600 1428.0600 1350.2600 1428.5400 ;
        RECT 1348.6600 1433.5000 1350.2600 1433.9800 ;
        RECT 1348.6600 1438.9400 1350.2600 1439.4200 ;
        RECT 1348.6600 1417.1800 1350.2600 1417.6600 ;
        RECT 1348.6600 1422.6200 1350.2600 1423.1000 ;
        RECT 1393.6600 1400.8600 1395.2600 1401.3400 ;
        RECT 1393.6600 1406.3000 1395.2600 1406.7800 ;
        RECT 1393.6600 1411.7400 1395.2600 1412.2200 ;
        RECT 1393.6600 1389.9800 1395.2600 1390.4600 ;
        RECT 1393.6600 1395.4200 1395.2600 1395.9000 ;
        RECT 1348.6600 1400.8600 1350.2600 1401.3400 ;
        RECT 1348.6600 1406.3000 1350.2600 1406.7800 ;
        RECT 1348.6600 1411.7400 1350.2600 1412.2200 ;
        RECT 1348.6600 1389.9800 1350.2600 1390.4600 ;
        RECT 1348.6600 1395.4200 1350.2600 1395.9000 ;
        RECT 1303.6600 1428.0600 1305.2600 1428.5400 ;
        RECT 1303.6600 1433.5000 1305.2600 1433.9800 ;
        RECT 1303.6600 1438.9400 1305.2600 1439.4200 ;
        RECT 1295.9000 1428.0600 1297.5000 1428.5400 ;
        RECT 1295.9000 1433.5000 1297.5000 1433.9800 ;
        RECT 1295.9000 1438.9400 1297.5000 1439.4200 ;
        RECT 1303.6600 1417.1800 1305.2600 1417.6600 ;
        RECT 1303.6600 1422.6200 1305.2600 1423.1000 ;
        RECT 1295.9000 1417.1800 1297.5000 1417.6600 ;
        RECT 1295.9000 1422.6200 1297.5000 1423.1000 ;
        RECT 1303.6600 1400.8600 1305.2600 1401.3400 ;
        RECT 1303.6600 1406.3000 1305.2600 1406.7800 ;
        RECT 1303.6600 1411.7400 1305.2600 1412.2200 ;
        RECT 1295.9000 1400.8600 1297.5000 1401.3400 ;
        RECT 1295.9000 1406.3000 1297.5000 1406.7800 ;
        RECT 1295.9000 1411.7400 1297.5000 1412.2200 ;
        RECT 1303.6600 1389.9800 1305.2600 1390.4600 ;
        RECT 1303.6600 1395.4200 1305.2600 1395.9000 ;
        RECT 1295.9000 1389.9800 1297.5000 1390.4600 ;
        RECT 1295.9000 1395.4200 1297.5000 1395.9000 ;
        RECT 1393.6600 1373.6600 1395.2600 1374.1400 ;
        RECT 1393.6600 1379.1000 1395.2600 1379.5800 ;
        RECT 1393.6600 1384.5400 1395.2600 1385.0200 ;
        RECT 1393.6600 1362.7800 1395.2600 1363.2600 ;
        RECT 1393.6600 1368.2200 1395.2600 1368.7000 ;
        RECT 1348.6600 1373.6600 1350.2600 1374.1400 ;
        RECT 1348.6600 1379.1000 1350.2600 1379.5800 ;
        RECT 1348.6600 1384.5400 1350.2600 1385.0200 ;
        RECT 1348.6600 1362.7800 1350.2600 1363.2600 ;
        RECT 1348.6600 1368.2200 1350.2600 1368.7000 ;
        RECT 1393.6600 1346.4600 1395.2600 1346.9400 ;
        RECT 1393.6600 1351.9000 1395.2600 1352.3800 ;
        RECT 1393.6600 1357.3400 1395.2600 1357.8200 ;
        RECT 1393.6600 1341.0200 1395.2600 1341.5000 ;
        RECT 1348.6600 1346.4600 1350.2600 1346.9400 ;
        RECT 1348.6600 1351.9000 1350.2600 1352.3800 ;
        RECT 1348.6600 1357.3400 1350.2600 1357.8200 ;
        RECT 1348.6600 1341.0200 1350.2600 1341.5000 ;
        RECT 1303.6600 1373.6600 1305.2600 1374.1400 ;
        RECT 1303.6600 1379.1000 1305.2600 1379.5800 ;
        RECT 1303.6600 1384.5400 1305.2600 1385.0200 ;
        RECT 1295.9000 1373.6600 1297.5000 1374.1400 ;
        RECT 1295.9000 1379.1000 1297.5000 1379.5800 ;
        RECT 1295.9000 1384.5400 1297.5000 1385.0200 ;
        RECT 1303.6600 1362.7800 1305.2600 1363.2600 ;
        RECT 1303.6600 1368.2200 1305.2600 1368.7000 ;
        RECT 1295.9000 1362.7800 1297.5000 1363.2600 ;
        RECT 1295.9000 1368.2200 1297.5000 1368.7000 ;
        RECT 1303.6600 1346.4600 1305.2600 1346.9400 ;
        RECT 1303.6600 1351.9000 1305.2600 1352.3800 ;
        RECT 1303.6600 1357.3400 1305.2600 1357.8200 ;
        RECT 1295.9000 1346.4600 1297.5000 1346.9400 ;
        RECT 1295.9000 1351.9000 1297.5000 1352.3800 ;
        RECT 1295.9000 1357.3400 1297.5000 1357.8200 ;
        RECT 1295.9000 1341.0200 1297.5000 1341.5000 ;
        RECT 1303.6600 1341.0200 1305.2600 1341.5000 ;
        RECT 1290.3400 1543.3300 1500.5600 1544.9300 ;
        RECT 1290.3400 1336.8300 1500.5600 1338.4300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1331.4000 1297.5000 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1549.4400 1297.5000 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1331.4000 1495.0000 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1549.4400 1495.0000 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1336.8300 1291.9400 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1336.8300 1500.5600 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1543.3300 1291.9400 1544.9300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1543.3300 1500.5600 1544.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 1107.1900 1485.2600 1315.2900 ;
        RECT 1438.6600 1107.1900 1440.2600 1315.2900 ;
        RECT 1393.6600 1107.1900 1395.2600 1315.2900 ;
        RECT 1348.6600 1107.1900 1350.2600 1315.2900 ;
        RECT 1303.6600 1107.1900 1305.2600 1315.2900 ;
        RECT 1493.4000 1101.7600 1495.0000 1321.4000 ;
        RECT 1295.9000 1101.7600 1297.5000 1321.4000 ;
      LAYER met3 ;
        RECT 1493.4000 1296.3400 1495.0000 1296.8200 ;
        RECT 1493.4000 1301.7800 1495.0000 1302.2600 ;
        RECT 1483.6600 1296.3400 1485.2600 1296.8200 ;
        RECT 1483.6600 1301.7800 1485.2600 1302.2600 ;
        RECT 1483.6600 1307.2200 1485.2600 1307.7000 ;
        RECT 1493.4000 1307.2200 1495.0000 1307.7000 ;
        RECT 1493.4000 1285.4600 1495.0000 1285.9400 ;
        RECT 1493.4000 1290.9000 1495.0000 1291.3800 ;
        RECT 1483.6600 1285.4600 1485.2600 1285.9400 ;
        RECT 1483.6600 1290.9000 1485.2600 1291.3800 ;
        RECT 1493.4000 1269.1400 1495.0000 1269.6200 ;
        RECT 1493.4000 1274.5800 1495.0000 1275.0600 ;
        RECT 1483.6600 1269.1400 1485.2600 1269.6200 ;
        RECT 1483.6600 1274.5800 1485.2600 1275.0600 ;
        RECT 1483.6600 1280.0200 1485.2600 1280.5000 ;
        RECT 1493.4000 1280.0200 1495.0000 1280.5000 ;
        RECT 1438.6600 1296.3400 1440.2600 1296.8200 ;
        RECT 1438.6600 1301.7800 1440.2600 1302.2600 ;
        RECT 1438.6600 1307.2200 1440.2600 1307.7000 ;
        RECT 1438.6600 1285.4600 1440.2600 1285.9400 ;
        RECT 1438.6600 1290.9000 1440.2600 1291.3800 ;
        RECT 1438.6600 1269.1400 1440.2600 1269.6200 ;
        RECT 1438.6600 1274.5800 1440.2600 1275.0600 ;
        RECT 1438.6600 1280.0200 1440.2600 1280.5000 ;
        RECT 1493.4000 1252.8200 1495.0000 1253.3000 ;
        RECT 1493.4000 1258.2600 1495.0000 1258.7400 ;
        RECT 1493.4000 1263.7000 1495.0000 1264.1800 ;
        RECT 1483.6600 1252.8200 1485.2600 1253.3000 ;
        RECT 1483.6600 1258.2600 1485.2600 1258.7400 ;
        RECT 1483.6600 1263.7000 1485.2600 1264.1800 ;
        RECT 1493.4000 1241.9400 1495.0000 1242.4200 ;
        RECT 1493.4000 1247.3800 1495.0000 1247.8600 ;
        RECT 1483.6600 1241.9400 1485.2600 1242.4200 ;
        RECT 1483.6600 1247.3800 1485.2600 1247.8600 ;
        RECT 1493.4000 1225.6200 1495.0000 1226.1000 ;
        RECT 1493.4000 1231.0600 1495.0000 1231.5400 ;
        RECT 1493.4000 1236.5000 1495.0000 1236.9800 ;
        RECT 1483.6600 1225.6200 1485.2600 1226.1000 ;
        RECT 1483.6600 1231.0600 1485.2600 1231.5400 ;
        RECT 1483.6600 1236.5000 1485.2600 1236.9800 ;
        RECT 1493.4000 1214.7400 1495.0000 1215.2200 ;
        RECT 1493.4000 1220.1800 1495.0000 1220.6600 ;
        RECT 1483.6600 1214.7400 1485.2600 1215.2200 ;
        RECT 1483.6600 1220.1800 1485.2600 1220.6600 ;
        RECT 1438.6600 1252.8200 1440.2600 1253.3000 ;
        RECT 1438.6600 1258.2600 1440.2600 1258.7400 ;
        RECT 1438.6600 1263.7000 1440.2600 1264.1800 ;
        RECT 1438.6600 1241.9400 1440.2600 1242.4200 ;
        RECT 1438.6600 1247.3800 1440.2600 1247.8600 ;
        RECT 1438.6600 1225.6200 1440.2600 1226.1000 ;
        RECT 1438.6600 1231.0600 1440.2600 1231.5400 ;
        RECT 1438.6600 1236.5000 1440.2600 1236.9800 ;
        RECT 1438.6600 1214.7400 1440.2600 1215.2200 ;
        RECT 1438.6600 1220.1800 1440.2600 1220.6600 ;
        RECT 1393.6600 1296.3400 1395.2600 1296.8200 ;
        RECT 1393.6600 1301.7800 1395.2600 1302.2600 ;
        RECT 1393.6600 1307.2200 1395.2600 1307.7000 ;
        RECT 1348.6600 1296.3400 1350.2600 1296.8200 ;
        RECT 1348.6600 1301.7800 1350.2600 1302.2600 ;
        RECT 1348.6600 1307.2200 1350.2600 1307.7000 ;
        RECT 1393.6600 1285.4600 1395.2600 1285.9400 ;
        RECT 1393.6600 1290.9000 1395.2600 1291.3800 ;
        RECT 1393.6600 1269.1400 1395.2600 1269.6200 ;
        RECT 1393.6600 1274.5800 1395.2600 1275.0600 ;
        RECT 1393.6600 1280.0200 1395.2600 1280.5000 ;
        RECT 1348.6600 1285.4600 1350.2600 1285.9400 ;
        RECT 1348.6600 1290.9000 1350.2600 1291.3800 ;
        RECT 1348.6600 1269.1400 1350.2600 1269.6200 ;
        RECT 1348.6600 1274.5800 1350.2600 1275.0600 ;
        RECT 1348.6600 1280.0200 1350.2600 1280.5000 ;
        RECT 1303.6600 1296.3400 1305.2600 1296.8200 ;
        RECT 1303.6600 1301.7800 1305.2600 1302.2600 ;
        RECT 1295.9000 1296.3400 1297.5000 1296.8200 ;
        RECT 1295.9000 1301.7800 1297.5000 1302.2600 ;
        RECT 1295.9000 1307.2200 1297.5000 1307.7000 ;
        RECT 1303.6600 1307.2200 1305.2600 1307.7000 ;
        RECT 1303.6600 1285.4600 1305.2600 1285.9400 ;
        RECT 1303.6600 1290.9000 1305.2600 1291.3800 ;
        RECT 1295.9000 1285.4600 1297.5000 1285.9400 ;
        RECT 1295.9000 1290.9000 1297.5000 1291.3800 ;
        RECT 1303.6600 1269.1400 1305.2600 1269.6200 ;
        RECT 1303.6600 1274.5800 1305.2600 1275.0600 ;
        RECT 1295.9000 1269.1400 1297.5000 1269.6200 ;
        RECT 1295.9000 1274.5800 1297.5000 1275.0600 ;
        RECT 1295.9000 1280.0200 1297.5000 1280.5000 ;
        RECT 1303.6600 1280.0200 1305.2600 1280.5000 ;
        RECT 1393.6600 1252.8200 1395.2600 1253.3000 ;
        RECT 1393.6600 1258.2600 1395.2600 1258.7400 ;
        RECT 1393.6600 1263.7000 1395.2600 1264.1800 ;
        RECT 1393.6600 1241.9400 1395.2600 1242.4200 ;
        RECT 1393.6600 1247.3800 1395.2600 1247.8600 ;
        RECT 1348.6600 1252.8200 1350.2600 1253.3000 ;
        RECT 1348.6600 1258.2600 1350.2600 1258.7400 ;
        RECT 1348.6600 1263.7000 1350.2600 1264.1800 ;
        RECT 1348.6600 1241.9400 1350.2600 1242.4200 ;
        RECT 1348.6600 1247.3800 1350.2600 1247.8600 ;
        RECT 1393.6600 1225.6200 1395.2600 1226.1000 ;
        RECT 1393.6600 1231.0600 1395.2600 1231.5400 ;
        RECT 1393.6600 1236.5000 1395.2600 1236.9800 ;
        RECT 1393.6600 1214.7400 1395.2600 1215.2200 ;
        RECT 1393.6600 1220.1800 1395.2600 1220.6600 ;
        RECT 1348.6600 1225.6200 1350.2600 1226.1000 ;
        RECT 1348.6600 1231.0600 1350.2600 1231.5400 ;
        RECT 1348.6600 1236.5000 1350.2600 1236.9800 ;
        RECT 1348.6600 1214.7400 1350.2600 1215.2200 ;
        RECT 1348.6600 1220.1800 1350.2600 1220.6600 ;
        RECT 1303.6600 1252.8200 1305.2600 1253.3000 ;
        RECT 1303.6600 1258.2600 1305.2600 1258.7400 ;
        RECT 1303.6600 1263.7000 1305.2600 1264.1800 ;
        RECT 1295.9000 1252.8200 1297.5000 1253.3000 ;
        RECT 1295.9000 1258.2600 1297.5000 1258.7400 ;
        RECT 1295.9000 1263.7000 1297.5000 1264.1800 ;
        RECT 1303.6600 1241.9400 1305.2600 1242.4200 ;
        RECT 1303.6600 1247.3800 1305.2600 1247.8600 ;
        RECT 1295.9000 1241.9400 1297.5000 1242.4200 ;
        RECT 1295.9000 1247.3800 1297.5000 1247.8600 ;
        RECT 1303.6600 1225.6200 1305.2600 1226.1000 ;
        RECT 1303.6600 1231.0600 1305.2600 1231.5400 ;
        RECT 1303.6600 1236.5000 1305.2600 1236.9800 ;
        RECT 1295.9000 1225.6200 1297.5000 1226.1000 ;
        RECT 1295.9000 1231.0600 1297.5000 1231.5400 ;
        RECT 1295.9000 1236.5000 1297.5000 1236.9800 ;
        RECT 1303.6600 1214.7400 1305.2600 1215.2200 ;
        RECT 1303.6600 1220.1800 1305.2600 1220.6600 ;
        RECT 1295.9000 1214.7400 1297.5000 1215.2200 ;
        RECT 1295.9000 1220.1800 1297.5000 1220.6600 ;
        RECT 1493.4000 1198.4200 1495.0000 1198.9000 ;
        RECT 1493.4000 1203.8600 1495.0000 1204.3400 ;
        RECT 1493.4000 1209.3000 1495.0000 1209.7800 ;
        RECT 1483.6600 1198.4200 1485.2600 1198.9000 ;
        RECT 1483.6600 1203.8600 1485.2600 1204.3400 ;
        RECT 1483.6600 1209.3000 1485.2600 1209.7800 ;
        RECT 1493.4000 1187.5400 1495.0000 1188.0200 ;
        RECT 1493.4000 1192.9800 1495.0000 1193.4600 ;
        RECT 1483.6600 1187.5400 1485.2600 1188.0200 ;
        RECT 1483.6600 1192.9800 1485.2600 1193.4600 ;
        RECT 1493.4000 1171.2200 1495.0000 1171.7000 ;
        RECT 1493.4000 1176.6600 1495.0000 1177.1400 ;
        RECT 1493.4000 1182.1000 1495.0000 1182.5800 ;
        RECT 1483.6600 1171.2200 1485.2600 1171.7000 ;
        RECT 1483.6600 1176.6600 1485.2600 1177.1400 ;
        RECT 1483.6600 1182.1000 1485.2600 1182.5800 ;
        RECT 1493.4000 1160.3400 1495.0000 1160.8200 ;
        RECT 1493.4000 1165.7800 1495.0000 1166.2600 ;
        RECT 1483.6600 1160.3400 1485.2600 1160.8200 ;
        RECT 1483.6600 1165.7800 1485.2600 1166.2600 ;
        RECT 1438.6600 1198.4200 1440.2600 1198.9000 ;
        RECT 1438.6600 1203.8600 1440.2600 1204.3400 ;
        RECT 1438.6600 1209.3000 1440.2600 1209.7800 ;
        RECT 1438.6600 1187.5400 1440.2600 1188.0200 ;
        RECT 1438.6600 1192.9800 1440.2600 1193.4600 ;
        RECT 1438.6600 1171.2200 1440.2600 1171.7000 ;
        RECT 1438.6600 1176.6600 1440.2600 1177.1400 ;
        RECT 1438.6600 1182.1000 1440.2600 1182.5800 ;
        RECT 1438.6600 1160.3400 1440.2600 1160.8200 ;
        RECT 1438.6600 1165.7800 1440.2600 1166.2600 ;
        RECT 1493.4000 1144.0200 1495.0000 1144.5000 ;
        RECT 1493.4000 1149.4600 1495.0000 1149.9400 ;
        RECT 1493.4000 1154.9000 1495.0000 1155.3800 ;
        RECT 1483.6600 1144.0200 1485.2600 1144.5000 ;
        RECT 1483.6600 1149.4600 1485.2600 1149.9400 ;
        RECT 1483.6600 1154.9000 1485.2600 1155.3800 ;
        RECT 1493.4000 1133.1400 1495.0000 1133.6200 ;
        RECT 1493.4000 1138.5800 1495.0000 1139.0600 ;
        RECT 1483.6600 1133.1400 1485.2600 1133.6200 ;
        RECT 1483.6600 1138.5800 1485.2600 1139.0600 ;
        RECT 1493.4000 1116.8200 1495.0000 1117.3000 ;
        RECT 1493.4000 1122.2600 1495.0000 1122.7400 ;
        RECT 1493.4000 1127.7000 1495.0000 1128.1800 ;
        RECT 1483.6600 1116.8200 1485.2600 1117.3000 ;
        RECT 1483.6600 1122.2600 1485.2600 1122.7400 ;
        RECT 1483.6600 1127.7000 1485.2600 1128.1800 ;
        RECT 1483.6600 1111.3800 1485.2600 1111.8600 ;
        RECT 1493.4000 1111.3800 1495.0000 1111.8600 ;
        RECT 1438.6600 1144.0200 1440.2600 1144.5000 ;
        RECT 1438.6600 1149.4600 1440.2600 1149.9400 ;
        RECT 1438.6600 1154.9000 1440.2600 1155.3800 ;
        RECT 1438.6600 1133.1400 1440.2600 1133.6200 ;
        RECT 1438.6600 1138.5800 1440.2600 1139.0600 ;
        RECT 1438.6600 1116.8200 1440.2600 1117.3000 ;
        RECT 1438.6600 1122.2600 1440.2600 1122.7400 ;
        RECT 1438.6600 1127.7000 1440.2600 1128.1800 ;
        RECT 1438.6600 1111.3800 1440.2600 1111.8600 ;
        RECT 1393.6600 1198.4200 1395.2600 1198.9000 ;
        RECT 1393.6600 1203.8600 1395.2600 1204.3400 ;
        RECT 1393.6600 1209.3000 1395.2600 1209.7800 ;
        RECT 1393.6600 1187.5400 1395.2600 1188.0200 ;
        RECT 1393.6600 1192.9800 1395.2600 1193.4600 ;
        RECT 1348.6600 1198.4200 1350.2600 1198.9000 ;
        RECT 1348.6600 1203.8600 1350.2600 1204.3400 ;
        RECT 1348.6600 1209.3000 1350.2600 1209.7800 ;
        RECT 1348.6600 1187.5400 1350.2600 1188.0200 ;
        RECT 1348.6600 1192.9800 1350.2600 1193.4600 ;
        RECT 1393.6600 1171.2200 1395.2600 1171.7000 ;
        RECT 1393.6600 1176.6600 1395.2600 1177.1400 ;
        RECT 1393.6600 1182.1000 1395.2600 1182.5800 ;
        RECT 1393.6600 1160.3400 1395.2600 1160.8200 ;
        RECT 1393.6600 1165.7800 1395.2600 1166.2600 ;
        RECT 1348.6600 1171.2200 1350.2600 1171.7000 ;
        RECT 1348.6600 1176.6600 1350.2600 1177.1400 ;
        RECT 1348.6600 1182.1000 1350.2600 1182.5800 ;
        RECT 1348.6600 1160.3400 1350.2600 1160.8200 ;
        RECT 1348.6600 1165.7800 1350.2600 1166.2600 ;
        RECT 1303.6600 1198.4200 1305.2600 1198.9000 ;
        RECT 1303.6600 1203.8600 1305.2600 1204.3400 ;
        RECT 1303.6600 1209.3000 1305.2600 1209.7800 ;
        RECT 1295.9000 1198.4200 1297.5000 1198.9000 ;
        RECT 1295.9000 1203.8600 1297.5000 1204.3400 ;
        RECT 1295.9000 1209.3000 1297.5000 1209.7800 ;
        RECT 1303.6600 1187.5400 1305.2600 1188.0200 ;
        RECT 1303.6600 1192.9800 1305.2600 1193.4600 ;
        RECT 1295.9000 1187.5400 1297.5000 1188.0200 ;
        RECT 1295.9000 1192.9800 1297.5000 1193.4600 ;
        RECT 1303.6600 1171.2200 1305.2600 1171.7000 ;
        RECT 1303.6600 1176.6600 1305.2600 1177.1400 ;
        RECT 1303.6600 1182.1000 1305.2600 1182.5800 ;
        RECT 1295.9000 1171.2200 1297.5000 1171.7000 ;
        RECT 1295.9000 1176.6600 1297.5000 1177.1400 ;
        RECT 1295.9000 1182.1000 1297.5000 1182.5800 ;
        RECT 1303.6600 1160.3400 1305.2600 1160.8200 ;
        RECT 1303.6600 1165.7800 1305.2600 1166.2600 ;
        RECT 1295.9000 1160.3400 1297.5000 1160.8200 ;
        RECT 1295.9000 1165.7800 1297.5000 1166.2600 ;
        RECT 1393.6600 1144.0200 1395.2600 1144.5000 ;
        RECT 1393.6600 1149.4600 1395.2600 1149.9400 ;
        RECT 1393.6600 1154.9000 1395.2600 1155.3800 ;
        RECT 1393.6600 1133.1400 1395.2600 1133.6200 ;
        RECT 1393.6600 1138.5800 1395.2600 1139.0600 ;
        RECT 1348.6600 1144.0200 1350.2600 1144.5000 ;
        RECT 1348.6600 1149.4600 1350.2600 1149.9400 ;
        RECT 1348.6600 1154.9000 1350.2600 1155.3800 ;
        RECT 1348.6600 1133.1400 1350.2600 1133.6200 ;
        RECT 1348.6600 1138.5800 1350.2600 1139.0600 ;
        RECT 1393.6600 1116.8200 1395.2600 1117.3000 ;
        RECT 1393.6600 1122.2600 1395.2600 1122.7400 ;
        RECT 1393.6600 1127.7000 1395.2600 1128.1800 ;
        RECT 1393.6600 1111.3800 1395.2600 1111.8600 ;
        RECT 1348.6600 1116.8200 1350.2600 1117.3000 ;
        RECT 1348.6600 1122.2600 1350.2600 1122.7400 ;
        RECT 1348.6600 1127.7000 1350.2600 1128.1800 ;
        RECT 1348.6600 1111.3800 1350.2600 1111.8600 ;
        RECT 1303.6600 1144.0200 1305.2600 1144.5000 ;
        RECT 1303.6600 1149.4600 1305.2600 1149.9400 ;
        RECT 1303.6600 1154.9000 1305.2600 1155.3800 ;
        RECT 1295.9000 1144.0200 1297.5000 1144.5000 ;
        RECT 1295.9000 1149.4600 1297.5000 1149.9400 ;
        RECT 1295.9000 1154.9000 1297.5000 1155.3800 ;
        RECT 1303.6600 1133.1400 1305.2600 1133.6200 ;
        RECT 1303.6600 1138.5800 1305.2600 1139.0600 ;
        RECT 1295.9000 1133.1400 1297.5000 1133.6200 ;
        RECT 1295.9000 1138.5800 1297.5000 1139.0600 ;
        RECT 1303.6600 1116.8200 1305.2600 1117.3000 ;
        RECT 1303.6600 1122.2600 1305.2600 1122.7400 ;
        RECT 1303.6600 1127.7000 1305.2600 1128.1800 ;
        RECT 1295.9000 1116.8200 1297.5000 1117.3000 ;
        RECT 1295.9000 1122.2600 1297.5000 1122.7400 ;
        RECT 1295.9000 1127.7000 1297.5000 1128.1800 ;
        RECT 1295.9000 1111.3800 1297.5000 1111.8600 ;
        RECT 1303.6600 1111.3800 1305.2600 1111.8600 ;
        RECT 1290.3400 1313.6900 1500.5600 1315.2900 ;
        RECT 1290.3400 1107.1900 1500.5600 1108.7900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1101.7600 1297.5000 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1319.8000 1297.5000 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1101.7600 1495.0000 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1319.8000 1495.0000 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1107.1900 1291.9400 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1107.1900 1500.5600 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1313.6900 1291.9400 1315.2900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1313.6900 1500.5600 1315.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 877.5500 1485.2600 1085.6500 ;
        RECT 1438.6600 877.5500 1440.2600 1085.6500 ;
        RECT 1393.6600 877.5500 1395.2600 1085.6500 ;
        RECT 1348.6600 877.5500 1350.2600 1085.6500 ;
        RECT 1303.6600 877.5500 1305.2600 1085.6500 ;
        RECT 1493.4000 872.1200 1495.0000 1091.7600 ;
        RECT 1295.9000 872.1200 1297.5000 1091.7600 ;
      LAYER met3 ;
        RECT 1493.4000 1066.7000 1495.0000 1067.1800 ;
        RECT 1493.4000 1072.1400 1495.0000 1072.6200 ;
        RECT 1483.6600 1066.7000 1485.2600 1067.1800 ;
        RECT 1483.6600 1072.1400 1485.2600 1072.6200 ;
        RECT 1483.6600 1077.5800 1485.2600 1078.0600 ;
        RECT 1493.4000 1077.5800 1495.0000 1078.0600 ;
        RECT 1493.4000 1055.8200 1495.0000 1056.3000 ;
        RECT 1493.4000 1061.2600 1495.0000 1061.7400 ;
        RECT 1483.6600 1055.8200 1485.2600 1056.3000 ;
        RECT 1483.6600 1061.2600 1485.2600 1061.7400 ;
        RECT 1493.4000 1039.5000 1495.0000 1039.9800 ;
        RECT 1493.4000 1044.9400 1495.0000 1045.4200 ;
        RECT 1483.6600 1039.5000 1485.2600 1039.9800 ;
        RECT 1483.6600 1044.9400 1485.2600 1045.4200 ;
        RECT 1483.6600 1050.3800 1485.2600 1050.8600 ;
        RECT 1493.4000 1050.3800 1495.0000 1050.8600 ;
        RECT 1438.6600 1066.7000 1440.2600 1067.1800 ;
        RECT 1438.6600 1072.1400 1440.2600 1072.6200 ;
        RECT 1438.6600 1077.5800 1440.2600 1078.0600 ;
        RECT 1438.6600 1055.8200 1440.2600 1056.3000 ;
        RECT 1438.6600 1061.2600 1440.2600 1061.7400 ;
        RECT 1438.6600 1039.5000 1440.2600 1039.9800 ;
        RECT 1438.6600 1044.9400 1440.2600 1045.4200 ;
        RECT 1438.6600 1050.3800 1440.2600 1050.8600 ;
        RECT 1493.4000 1023.1800 1495.0000 1023.6600 ;
        RECT 1493.4000 1028.6200 1495.0000 1029.1000 ;
        RECT 1493.4000 1034.0600 1495.0000 1034.5400 ;
        RECT 1483.6600 1023.1800 1485.2600 1023.6600 ;
        RECT 1483.6600 1028.6200 1485.2600 1029.1000 ;
        RECT 1483.6600 1034.0600 1485.2600 1034.5400 ;
        RECT 1493.4000 1012.3000 1495.0000 1012.7800 ;
        RECT 1493.4000 1017.7400 1495.0000 1018.2200 ;
        RECT 1483.6600 1012.3000 1485.2600 1012.7800 ;
        RECT 1483.6600 1017.7400 1485.2600 1018.2200 ;
        RECT 1493.4000 995.9800 1495.0000 996.4600 ;
        RECT 1493.4000 1001.4200 1495.0000 1001.9000 ;
        RECT 1493.4000 1006.8600 1495.0000 1007.3400 ;
        RECT 1483.6600 995.9800 1485.2600 996.4600 ;
        RECT 1483.6600 1001.4200 1485.2600 1001.9000 ;
        RECT 1483.6600 1006.8600 1485.2600 1007.3400 ;
        RECT 1493.4000 985.1000 1495.0000 985.5800 ;
        RECT 1493.4000 990.5400 1495.0000 991.0200 ;
        RECT 1483.6600 985.1000 1485.2600 985.5800 ;
        RECT 1483.6600 990.5400 1485.2600 991.0200 ;
        RECT 1438.6600 1023.1800 1440.2600 1023.6600 ;
        RECT 1438.6600 1028.6200 1440.2600 1029.1000 ;
        RECT 1438.6600 1034.0600 1440.2600 1034.5400 ;
        RECT 1438.6600 1012.3000 1440.2600 1012.7800 ;
        RECT 1438.6600 1017.7400 1440.2600 1018.2200 ;
        RECT 1438.6600 995.9800 1440.2600 996.4600 ;
        RECT 1438.6600 1001.4200 1440.2600 1001.9000 ;
        RECT 1438.6600 1006.8600 1440.2600 1007.3400 ;
        RECT 1438.6600 985.1000 1440.2600 985.5800 ;
        RECT 1438.6600 990.5400 1440.2600 991.0200 ;
        RECT 1393.6600 1066.7000 1395.2600 1067.1800 ;
        RECT 1393.6600 1072.1400 1395.2600 1072.6200 ;
        RECT 1393.6600 1077.5800 1395.2600 1078.0600 ;
        RECT 1348.6600 1066.7000 1350.2600 1067.1800 ;
        RECT 1348.6600 1072.1400 1350.2600 1072.6200 ;
        RECT 1348.6600 1077.5800 1350.2600 1078.0600 ;
        RECT 1393.6600 1055.8200 1395.2600 1056.3000 ;
        RECT 1393.6600 1061.2600 1395.2600 1061.7400 ;
        RECT 1393.6600 1039.5000 1395.2600 1039.9800 ;
        RECT 1393.6600 1044.9400 1395.2600 1045.4200 ;
        RECT 1393.6600 1050.3800 1395.2600 1050.8600 ;
        RECT 1348.6600 1055.8200 1350.2600 1056.3000 ;
        RECT 1348.6600 1061.2600 1350.2600 1061.7400 ;
        RECT 1348.6600 1039.5000 1350.2600 1039.9800 ;
        RECT 1348.6600 1044.9400 1350.2600 1045.4200 ;
        RECT 1348.6600 1050.3800 1350.2600 1050.8600 ;
        RECT 1303.6600 1066.7000 1305.2600 1067.1800 ;
        RECT 1303.6600 1072.1400 1305.2600 1072.6200 ;
        RECT 1295.9000 1066.7000 1297.5000 1067.1800 ;
        RECT 1295.9000 1072.1400 1297.5000 1072.6200 ;
        RECT 1295.9000 1077.5800 1297.5000 1078.0600 ;
        RECT 1303.6600 1077.5800 1305.2600 1078.0600 ;
        RECT 1303.6600 1055.8200 1305.2600 1056.3000 ;
        RECT 1303.6600 1061.2600 1305.2600 1061.7400 ;
        RECT 1295.9000 1055.8200 1297.5000 1056.3000 ;
        RECT 1295.9000 1061.2600 1297.5000 1061.7400 ;
        RECT 1303.6600 1039.5000 1305.2600 1039.9800 ;
        RECT 1303.6600 1044.9400 1305.2600 1045.4200 ;
        RECT 1295.9000 1039.5000 1297.5000 1039.9800 ;
        RECT 1295.9000 1044.9400 1297.5000 1045.4200 ;
        RECT 1295.9000 1050.3800 1297.5000 1050.8600 ;
        RECT 1303.6600 1050.3800 1305.2600 1050.8600 ;
        RECT 1393.6600 1023.1800 1395.2600 1023.6600 ;
        RECT 1393.6600 1028.6200 1395.2600 1029.1000 ;
        RECT 1393.6600 1034.0600 1395.2600 1034.5400 ;
        RECT 1393.6600 1012.3000 1395.2600 1012.7800 ;
        RECT 1393.6600 1017.7400 1395.2600 1018.2200 ;
        RECT 1348.6600 1023.1800 1350.2600 1023.6600 ;
        RECT 1348.6600 1028.6200 1350.2600 1029.1000 ;
        RECT 1348.6600 1034.0600 1350.2600 1034.5400 ;
        RECT 1348.6600 1012.3000 1350.2600 1012.7800 ;
        RECT 1348.6600 1017.7400 1350.2600 1018.2200 ;
        RECT 1393.6600 995.9800 1395.2600 996.4600 ;
        RECT 1393.6600 1001.4200 1395.2600 1001.9000 ;
        RECT 1393.6600 1006.8600 1395.2600 1007.3400 ;
        RECT 1393.6600 985.1000 1395.2600 985.5800 ;
        RECT 1393.6600 990.5400 1395.2600 991.0200 ;
        RECT 1348.6600 995.9800 1350.2600 996.4600 ;
        RECT 1348.6600 1001.4200 1350.2600 1001.9000 ;
        RECT 1348.6600 1006.8600 1350.2600 1007.3400 ;
        RECT 1348.6600 985.1000 1350.2600 985.5800 ;
        RECT 1348.6600 990.5400 1350.2600 991.0200 ;
        RECT 1303.6600 1023.1800 1305.2600 1023.6600 ;
        RECT 1303.6600 1028.6200 1305.2600 1029.1000 ;
        RECT 1303.6600 1034.0600 1305.2600 1034.5400 ;
        RECT 1295.9000 1023.1800 1297.5000 1023.6600 ;
        RECT 1295.9000 1028.6200 1297.5000 1029.1000 ;
        RECT 1295.9000 1034.0600 1297.5000 1034.5400 ;
        RECT 1303.6600 1012.3000 1305.2600 1012.7800 ;
        RECT 1303.6600 1017.7400 1305.2600 1018.2200 ;
        RECT 1295.9000 1012.3000 1297.5000 1012.7800 ;
        RECT 1295.9000 1017.7400 1297.5000 1018.2200 ;
        RECT 1303.6600 995.9800 1305.2600 996.4600 ;
        RECT 1303.6600 1001.4200 1305.2600 1001.9000 ;
        RECT 1303.6600 1006.8600 1305.2600 1007.3400 ;
        RECT 1295.9000 995.9800 1297.5000 996.4600 ;
        RECT 1295.9000 1001.4200 1297.5000 1001.9000 ;
        RECT 1295.9000 1006.8600 1297.5000 1007.3400 ;
        RECT 1303.6600 985.1000 1305.2600 985.5800 ;
        RECT 1303.6600 990.5400 1305.2600 991.0200 ;
        RECT 1295.9000 985.1000 1297.5000 985.5800 ;
        RECT 1295.9000 990.5400 1297.5000 991.0200 ;
        RECT 1493.4000 968.7800 1495.0000 969.2600 ;
        RECT 1493.4000 974.2200 1495.0000 974.7000 ;
        RECT 1493.4000 979.6600 1495.0000 980.1400 ;
        RECT 1483.6600 968.7800 1485.2600 969.2600 ;
        RECT 1483.6600 974.2200 1485.2600 974.7000 ;
        RECT 1483.6600 979.6600 1485.2600 980.1400 ;
        RECT 1493.4000 957.9000 1495.0000 958.3800 ;
        RECT 1493.4000 963.3400 1495.0000 963.8200 ;
        RECT 1483.6600 957.9000 1485.2600 958.3800 ;
        RECT 1483.6600 963.3400 1485.2600 963.8200 ;
        RECT 1493.4000 941.5800 1495.0000 942.0600 ;
        RECT 1493.4000 947.0200 1495.0000 947.5000 ;
        RECT 1493.4000 952.4600 1495.0000 952.9400 ;
        RECT 1483.6600 941.5800 1485.2600 942.0600 ;
        RECT 1483.6600 947.0200 1485.2600 947.5000 ;
        RECT 1483.6600 952.4600 1485.2600 952.9400 ;
        RECT 1493.4000 930.7000 1495.0000 931.1800 ;
        RECT 1493.4000 936.1400 1495.0000 936.6200 ;
        RECT 1483.6600 930.7000 1485.2600 931.1800 ;
        RECT 1483.6600 936.1400 1485.2600 936.6200 ;
        RECT 1438.6600 968.7800 1440.2600 969.2600 ;
        RECT 1438.6600 974.2200 1440.2600 974.7000 ;
        RECT 1438.6600 979.6600 1440.2600 980.1400 ;
        RECT 1438.6600 957.9000 1440.2600 958.3800 ;
        RECT 1438.6600 963.3400 1440.2600 963.8200 ;
        RECT 1438.6600 941.5800 1440.2600 942.0600 ;
        RECT 1438.6600 947.0200 1440.2600 947.5000 ;
        RECT 1438.6600 952.4600 1440.2600 952.9400 ;
        RECT 1438.6600 930.7000 1440.2600 931.1800 ;
        RECT 1438.6600 936.1400 1440.2600 936.6200 ;
        RECT 1493.4000 914.3800 1495.0000 914.8600 ;
        RECT 1493.4000 919.8200 1495.0000 920.3000 ;
        RECT 1493.4000 925.2600 1495.0000 925.7400 ;
        RECT 1483.6600 914.3800 1485.2600 914.8600 ;
        RECT 1483.6600 919.8200 1485.2600 920.3000 ;
        RECT 1483.6600 925.2600 1485.2600 925.7400 ;
        RECT 1493.4000 903.5000 1495.0000 903.9800 ;
        RECT 1493.4000 908.9400 1495.0000 909.4200 ;
        RECT 1483.6600 903.5000 1485.2600 903.9800 ;
        RECT 1483.6600 908.9400 1485.2600 909.4200 ;
        RECT 1493.4000 887.1800 1495.0000 887.6600 ;
        RECT 1493.4000 892.6200 1495.0000 893.1000 ;
        RECT 1493.4000 898.0600 1495.0000 898.5400 ;
        RECT 1483.6600 887.1800 1485.2600 887.6600 ;
        RECT 1483.6600 892.6200 1485.2600 893.1000 ;
        RECT 1483.6600 898.0600 1485.2600 898.5400 ;
        RECT 1483.6600 881.7400 1485.2600 882.2200 ;
        RECT 1493.4000 881.7400 1495.0000 882.2200 ;
        RECT 1438.6600 914.3800 1440.2600 914.8600 ;
        RECT 1438.6600 919.8200 1440.2600 920.3000 ;
        RECT 1438.6600 925.2600 1440.2600 925.7400 ;
        RECT 1438.6600 903.5000 1440.2600 903.9800 ;
        RECT 1438.6600 908.9400 1440.2600 909.4200 ;
        RECT 1438.6600 887.1800 1440.2600 887.6600 ;
        RECT 1438.6600 892.6200 1440.2600 893.1000 ;
        RECT 1438.6600 898.0600 1440.2600 898.5400 ;
        RECT 1438.6600 881.7400 1440.2600 882.2200 ;
        RECT 1393.6600 968.7800 1395.2600 969.2600 ;
        RECT 1393.6600 974.2200 1395.2600 974.7000 ;
        RECT 1393.6600 979.6600 1395.2600 980.1400 ;
        RECT 1393.6600 957.9000 1395.2600 958.3800 ;
        RECT 1393.6600 963.3400 1395.2600 963.8200 ;
        RECT 1348.6600 968.7800 1350.2600 969.2600 ;
        RECT 1348.6600 974.2200 1350.2600 974.7000 ;
        RECT 1348.6600 979.6600 1350.2600 980.1400 ;
        RECT 1348.6600 957.9000 1350.2600 958.3800 ;
        RECT 1348.6600 963.3400 1350.2600 963.8200 ;
        RECT 1393.6600 941.5800 1395.2600 942.0600 ;
        RECT 1393.6600 947.0200 1395.2600 947.5000 ;
        RECT 1393.6600 952.4600 1395.2600 952.9400 ;
        RECT 1393.6600 930.7000 1395.2600 931.1800 ;
        RECT 1393.6600 936.1400 1395.2600 936.6200 ;
        RECT 1348.6600 941.5800 1350.2600 942.0600 ;
        RECT 1348.6600 947.0200 1350.2600 947.5000 ;
        RECT 1348.6600 952.4600 1350.2600 952.9400 ;
        RECT 1348.6600 930.7000 1350.2600 931.1800 ;
        RECT 1348.6600 936.1400 1350.2600 936.6200 ;
        RECT 1303.6600 968.7800 1305.2600 969.2600 ;
        RECT 1303.6600 974.2200 1305.2600 974.7000 ;
        RECT 1303.6600 979.6600 1305.2600 980.1400 ;
        RECT 1295.9000 968.7800 1297.5000 969.2600 ;
        RECT 1295.9000 974.2200 1297.5000 974.7000 ;
        RECT 1295.9000 979.6600 1297.5000 980.1400 ;
        RECT 1303.6600 957.9000 1305.2600 958.3800 ;
        RECT 1303.6600 963.3400 1305.2600 963.8200 ;
        RECT 1295.9000 957.9000 1297.5000 958.3800 ;
        RECT 1295.9000 963.3400 1297.5000 963.8200 ;
        RECT 1303.6600 941.5800 1305.2600 942.0600 ;
        RECT 1303.6600 947.0200 1305.2600 947.5000 ;
        RECT 1303.6600 952.4600 1305.2600 952.9400 ;
        RECT 1295.9000 941.5800 1297.5000 942.0600 ;
        RECT 1295.9000 947.0200 1297.5000 947.5000 ;
        RECT 1295.9000 952.4600 1297.5000 952.9400 ;
        RECT 1303.6600 930.7000 1305.2600 931.1800 ;
        RECT 1303.6600 936.1400 1305.2600 936.6200 ;
        RECT 1295.9000 930.7000 1297.5000 931.1800 ;
        RECT 1295.9000 936.1400 1297.5000 936.6200 ;
        RECT 1393.6600 914.3800 1395.2600 914.8600 ;
        RECT 1393.6600 919.8200 1395.2600 920.3000 ;
        RECT 1393.6600 925.2600 1395.2600 925.7400 ;
        RECT 1393.6600 903.5000 1395.2600 903.9800 ;
        RECT 1393.6600 908.9400 1395.2600 909.4200 ;
        RECT 1348.6600 914.3800 1350.2600 914.8600 ;
        RECT 1348.6600 919.8200 1350.2600 920.3000 ;
        RECT 1348.6600 925.2600 1350.2600 925.7400 ;
        RECT 1348.6600 903.5000 1350.2600 903.9800 ;
        RECT 1348.6600 908.9400 1350.2600 909.4200 ;
        RECT 1393.6600 887.1800 1395.2600 887.6600 ;
        RECT 1393.6600 892.6200 1395.2600 893.1000 ;
        RECT 1393.6600 898.0600 1395.2600 898.5400 ;
        RECT 1393.6600 881.7400 1395.2600 882.2200 ;
        RECT 1348.6600 887.1800 1350.2600 887.6600 ;
        RECT 1348.6600 892.6200 1350.2600 893.1000 ;
        RECT 1348.6600 898.0600 1350.2600 898.5400 ;
        RECT 1348.6600 881.7400 1350.2600 882.2200 ;
        RECT 1303.6600 914.3800 1305.2600 914.8600 ;
        RECT 1303.6600 919.8200 1305.2600 920.3000 ;
        RECT 1303.6600 925.2600 1305.2600 925.7400 ;
        RECT 1295.9000 914.3800 1297.5000 914.8600 ;
        RECT 1295.9000 919.8200 1297.5000 920.3000 ;
        RECT 1295.9000 925.2600 1297.5000 925.7400 ;
        RECT 1303.6600 903.5000 1305.2600 903.9800 ;
        RECT 1303.6600 908.9400 1305.2600 909.4200 ;
        RECT 1295.9000 903.5000 1297.5000 903.9800 ;
        RECT 1295.9000 908.9400 1297.5000 909.4200 ;
        RECT 1303.6600 887.1800 1305.2600 887.6600 ;
        RECT 1303.6600 892.6200 1305.2600 893.1000 ;
        RECT 1303.6600 898.0600 1305.2600 898.5400 ;
        RECT 1295.9000 887.1800 1297.5000 887.6600 ;
        RECT 1295.9000 892.6200 1297.5000 893.1000 ;
        RECT 1295.9000 898.0600 1297.5000 898.5400 ;
        RECT 1295.9000 881.7400 1297.5000 882.2200 ;
        RECT 1303.6600 881.7400 1305.2600 882.2200 ;
        RECT 1290.3400 1084.0500 1500.5600 1085.6500 ;
        RECT 1290.3400 877.5500 1500.5600 879.1500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 872.1200 1297.5000 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 1090.1600 1297.5000 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 872.1200 1495.0000 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 1090.1600 1495.0000 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 877.5500 1291.9400 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 877.5500 1500.5600 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 1084.0500 1291.9400 1085.6500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 1084.0500 1500.5600 1085.6500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 647.9100 1485.2600 856.0100 ;
        RECT 1438.6600 647.9100 1440.2600 856.0100 ;
        RECT 1393.6600 647.9100 1395.2600 856.0100 ;
        RECT 1348.6600 647.9100 1350.2600 856.0100 ;
        RECT 1303.6600 647.9100 1305.2600 856.0100 ;
        RECT 1493.4000 642.4800 1495.0000 862.1200 ;
        RECT 1295.9000 642.4800 1297.5000 862.1200 ;
      LAYER met3 ;
        RECT 1493.4000 837.0600 1495.0000 837.5400 ;
        RECT 1493.4000 842.5000 1495.0000 842.9800 ;
        RECT 1483.6600 837.0600 1485.2600 837.5400 ;
        RECT 1483.6600 842.5000 1485.2600 842.9800 ;
        RECT 1483.6600 847.9400 1485.2600 848.4200 ;
        RECT 1493.4000 847.9400 1495.0000 848.4200 ;
        RECT 1493.4000 826.1800 1495.0000 826.6600 ;
        RECT 1493.4000 831.6200 1495.0000 832.1000 ;
        RECT 1483.6600 826.1800 1485.2600 826.6600 ;
        RECT 1483.6600 831.6200 1485.2600 832.1000 ;
        RECT 1493.4000 809.8600 1495.0000 810.3400 ;
        RECT 1493.4000 815.3000 1495.0000 815.7800 ;
        RECT 1483.6600 809.8600 1485.2600 810.3400 ;
        RECT 1483.6600 815.3000 1485.2600 815.7800 ;
        RECT 1483.6600 820.7400 1485.2600 821.2200 ;
        RECT 1493.4000 820.7400 1495.0000 821.2200 ;
        RECT 1438.6600 837.0600 1440.2600 837.5400 ;
        RECT 1438.6600 842.5000 1440.2600 842.9800 ;
        RECT 1438.6600 847.9400 1440.2600 848.4200 ;
        RECT 1438.6600 826.1800 1440.2600 826.6600 ;
        RECT 1438.6600 831.6200 1440.2600 832.1000 ;
        RECT 1438.6600 809.8600 1440.2600 810.3400 ;
        RECT 1438.6600 815.3000 1440.2600 815.7800 ;
        RECT 1438.6600 820.7400 1440.2600 821.2200 ;
        RECT 1493.4000 793.5400 1495.0000 794.0200 ;
        RECT 1493.4000 798.9800 1495.0000 799.4600 ;
        RECT 1493.4000 804.4200 1495.0000 804.9000 ;
        RECT 1483.6600 793.5400 1485.2600 794.0200 ;
        RECT 1483.6600 798.9800 1485.2600 799.4600 ;
        RECT 1483.6600 804.4200 1485.2600 804.9000 ;
        RECT 1493.4000 782.6600 1495.0000 783.1400 ;
        RECT 1493.4000 788.1000 1495.0000 788.5800 ;
        RECT 1483.6600 782.6600 1485.2600 783.1400 ;
        RECT 1483.6600 788.1000 1485.2600 788.5800 ;
        RECT 1493.4000 766.3400 1495.0000 766.8200 ;
        RECT 1493.4000 771.7800 1495.0000 772.2600 ;
        RECT 1493.4000 777.2200 1495.0000 777.7000 ;
        RECT 1483.6600 766.3400 1485.2600 766.8200 ;
        RECT 1483.6600 771.7800 1485.2600 772.2600 ;
        RECT 1483.6600 777.2200 1485.2600 777.7000 ;
        RECT 1493.4000 755.4600 1495.0000 755.9400 ;
        RECT 1493.4000 760.9000 1495.0000 761.3800 ;
        RECT 1483.6600 755.4600 1485.2600 755.9400 ;
        RECT 1483.6600 760.9000 1485.2600 761.3800 ;
        RECT 1438.6600 793.5400 1440.2600 794.0200 ;
        RECT 1438.6600 798.9800 1440.2600 799.4600 ;
        RECT 1438.6600 804.4200 1440.2600 804.9000 ;
        RECT 1438.6600 782.6600 1440.2600 783.1400 ;
        RECT 1438.6600 788.1000 1440.2600 788.5800 ;
        RECT 1438.6600 766.3400 1440.2600 766.8200 ;
        RECT 1438.6600 771.7800 1440.2600 772.2600 ;
        RECT 1438.6600 777.2200 1440.2600 777.7000 ;
        RECT 1438.6600 755.4600 1440.2600 755.9400 ;
        RECT 1438.6600 760.9000 1440.2600 761.3800 ;
        RECT 1393.6600 837.0600 1395.2600 837.5400 ;
        RECT 1393.6600 842.5000 1395.2600 842.9800 ;
        RECT 1393.6600 847.9400 1395.2600 848.4200 ;
        RECT 1348.6600 837.0600 1350.2600 837.5400 ;
        RECT 1348.6600 842.5000 1350.2600 842.9800 ;
        RECT 1348.6600 847.9400 1350.2600 848.4200 ;
        RECT 1393.6600 826.1800 1395.2600 826.6600 ;
        RECT 1393.6600 831.6200 1395.2600 832.1000 ;
        RECT 1393.6600 809.8600 1395.2600 810.3400 ;
        RECT 1393.6600 815.3000 1395.2600 815.7800 ;
        RECT 1393.6600 820.7400 1395.2600 821.2200 ;
        RECT 1348.6600 826.1800 1350.2600 826.6600 ;
        RECT 1348.6600 831.6200 1350.2600 832.1000 ;
        RECT 1348.6600 809.8600 1350.2600 810.3400 ;
        RECT 1348.6600 815.3000 1350.2600 815.7800 ;
        RECT 1348.6600 820.7400 1350.2600 821.2200 ;
        RECT 1303.6600 837.0600 1305.2600 837.5400 ;
        RECT 1303.6600 842.5000 1305.2600 842.9800 ;
        RECT 1295.9000 837.0600 1297.5000 837.5400 ;
        RECT 1295.9000 842.5000 1297.5000 842.9800 ;
        RECT 1295.9000 847.9400 1297.5000 848.4200 ;
        RECT 1303.6600 847.9400 1305.2600 848.4200 ;
        RECT 1303.6600 826.1800 1305.2600 826.6600 ;
        RECT 1303.6600 831.6200 1305.2600 832.1000 ;
        RECT 1295.9000 826.1800 1297.5000 826.6600 ;
        RECT 1295.9000 831.6200 1297.5000 832.1000 ;
        RECT 1303.6600 809.8600 1305.2600 810.3400 ;
        RECT 1303.6600 815.3000 1305.2600 815.7800 ;
        RECT 1295.9000 809.8600 1297.5000 810.3400 ;
        RECT 1295.9000 815.3000 1297.5000 815.7800 ;
        RECT 1295.9000 820.7400 1297.5000 821.2200 ;
        RECT 1303.6600 820.7400 1305.2600 821.2200 ;
        RECT 1393.6600 793.5400 1395.2600 794.0200 ;
        RECT 1393.6600 798.9800 1395.2600 799.4600 ;
        RECT 1393.6600 804.4200 1395.2600 804.9000 ;
        RECT 1393.6600 782.6600 1395.2600 783.1400 ;
        RECT 1393.6600 788.1000 1395.2600 788.5800 ;
        RECT 1348.6600 793.5400 1350.2600 794.0200 ;
        RECT 1348.6600 798.9800 1350.2600 799.4600 ;
        RECT 1348.6600 804.4200 1350.2600 804.9000 ;
        RECT 1348.6600 782.6600 1350.2600 783.1400 ;
        RECT 1348.6600 788.1000 1350.2600 788.5800 ;
        RECT 1393.6600 766.3400 1395.2600 766.8200 ;
        RECT 1393.6600 771.7800 1395.2600 772.2600 ;
        RECT 1393.6600 777.2200 1395.2600 777.7000 ;
        RECT 1393.6600 755.4600 1395.2600 755.9400 ;
        RECT 1393.6600 760.9000 1395.2600 761.3800 ;
        RECT 1348.6600 766.3400 1350.2600 766.8200 ;
        RECT 1348.6600 771.7800 1350.2600 772.2600 ;
        RECT 1348.6600 777.2200 1350.2600 777.7000 ;
        RECT 1348.6600 755.4600 1350.2600 755.9400 ;
        RECT 1348.6600 760.9000 1350.2600 761.3800 ;
        RECT 1303.6600 793.5400 1305.2600 794.0200 ;
        RECT 1303.6600 798.9800 1305.2600 799.4600 ;
        RECT 1303.6600 804.4200 1305.2600 804.9000 ;
        RECT 1295.9000 793.5400 1297.5000 794.0200 ;
        RECT 1295.9000 798.9800 1297.5000 799.4600 ;
        RECT 1295.9000 804.4200 1297.5000 804.9000 ;
        RECT 1303.6600 782.6600 1305.2600 783.1400 ;
        RECT 1303.6600 788.1000 1305.2600 788.5800 ;
        RECT 1295.9000 782.6600 1297.5000 783.1400 ;
        RECT 1295.9000 788.1000 1297.5000 788.5800 ;
        RECT 1303.6600 766.3400 1305.2600 766.8200 ;
        RECT 1303.6600 771.7800 1305.2600 772.2600 ;
        RECT 1303.6600 777.2200 1305.2600 777.7000 ;
        RECT 1295.9000 766.3400 1297.5000 766.8200 ;
        RECT 1295.9000 771.7800 1297.5000 772.2600 ;
        RECT 1295.9000 777.2200 1297.5000 777.7000 ;
        RECT 1303.6600 755.4600 1305.2600 755.9400 ;
        RECT 1303.6600 760.9000 1305.2600 761.3800 ;
        RECT 1295.9000 755.4600 1297.5000 755.9400 ;
        RECT 1295.9000 760.9000 1297.5000 761.3800 ;
        RECT 1493.4000 739.1400 1495.0000 739.6200 ;
        RECT 1493.4000 744.5800 1495.0000 745.0600 ;
        RECT 1493.4000 750.0200 1495.0000 750.5000 ;
        RECT 1483.6600 739.1400 1485.2600 739.6200 ;
        RECT 1483.6600 744.5800 1485.2600 745.0600 ;
        RECT 1483.6600 750.0200 1485.2600 750.5000 ;
        RECT 1493.4000 728.2600 1495.0000 728.7400 ;
        RECT 1493.4000 733.7000 1495.0000 734.1800 ;
        RECT 1483.6600 728.2600 1485.2600 728.7400 ;
        RECT 1483.6600 733.7000 1485.2600 734.1800 ;
        RECT 1493.4000 711.9400 1495.0000 712.4200 ;
        RECT 1493.4000 717.3800 1495.0000 717.8600 ;
        RECT 1493.4000 722.8200 1495.0000 723.3000 ;
        RECT 1483.6600 711.9400 1485.2600 712.4200 ;
        RECT 1483.6600 717.3800 1485.2600 717.8600 ;
        RECT 1483.6600 722.8200 1485.2600 723.3000 ;
        RECT 1493.4000 701.0600 1495.0000 701.5400 ;
        RECT 1493.4000 706.5000 1495.0000 706.9800 ;
        RECT 1483.6600 701.0600 1485.2600 701.5400 ;
        RECT 1483.6600 706.5000 1485.2600 706.9800 ;
        RECT 1438.6600 739.1400 1440.2600 739.6200 ;
        RECT 1438.6600 744.5800 1440.2600 745.0600 ;
        RECT 1438.6600 750.0200 1440.2600 750.5000 ;
        RECT 1438.6600 728.2600 1440.2600 728.7400 ;
        RECT 1438.6600 733.7000 1440.2600 734.1800 ;
        RECT 1438.6600 711.9400 1440.2600 712.4200 ;
        RECT 1438.6600 717.3800 1440.2600 717.8600 ;
        RECT 1438.6600 722.8200 1440.2600 723.3000 ;
        RECT 1438.6600 701.0600 1440.2600 701.5400 ;
        RECT 1438.6600 706.5000 1440.2600 706.9800 ;
        RECT 1493.4000 684.7400 1495.0000 685.2200 ;
        RECT 1493.4000 690.1800 1495.0000 690.6600 ;
        RECT 1493.4000 695.6200 1495.0000 696.1000 ;
        RECT 1483.6600 684.7400 1485.2600 685.2200 ;
        RECT 1483.6600 690.1800 1485.2600 690.6600 ;
        RECT 1483.6600 695.6200 1485.2600 696.1000 ;
        RECT 1493.4000 673.8600 1495.0000 674.3400 ;
        RECT 1493.4000 679.3000 1495.0000 679.7800 ;
        RECT 1483.6600 673.8600 1485.2600 674.3400 ;
        RECT 1483.6600 679.3000 1485.2600 679.7800 ;
        RECT 1493.4000 657.5400 1495.0000 658.0200 ;
        RECT 1493.4000 662.9800 1495.0000 663.4600 ;
        RECT 1493.4000 668.4200 1495.0000 668.9000 ;
        RECT 1483.6600 657.5400 1485.2600 658.0200 ;
        RECT 1483.6600 662.9800 1485.2600 663.4600 ;
        RECT 1483.6600 668.4200 1485.2600 668.9000 ;
        RECT 1483.6600 652.1000 1485.2600 652.5800 ;
        RECT 1493.4000 652.1000 1495.0000 652.5800 ;
        RECT 1438.6600 684.7400 1440.2600 685.2200 ;
        RECT 1438.6600 690.1800 1440.2600 690.6600 ;
        RECT 1438.6600 695.6200 1440.2600 696.1000 ;
        RECT 1438.6600 673.8600 1440.2600 674.3400 ;
        RECT 1438.6600 679.3000 1440.2600 679.7800 ;
        RECT 1438.6600 657.5400 1440.2600 658.0200 ;
        RECT 1438.6600 662.9800 1440.2600 663.4600 ;
        RECT 1438.6600 668.4200 1440.2600 668.9000 ;
        RECT 1438.6600 652.1000 1440.2600 652.5800 ;
        RECT 1393.6600 739.1400 1395.2600 739.6200 ;
        RECT 1393.6600 744.5800 1395.2600 745.0600 ;
        RECT 1393.6600 750.0200 1395.2600 750.5000 ;
        RECT 1393.6600 728.2600 1395.2600 728.7400 ;
        RECT 1393.6600 733.7000 1395.2600 734.1800 ;
        RECT 1348.6600 739.1400 1350.2600 739.6200 ;
        RECT 1348.6600 744.5800 1350.2600 745.0600 ;
        RECT 1348.6600 750.0200 1350.2600 750.5000 ;
        RECT 1348.6600 728.2600 1350.2600 728.7400 ;
        RECT 1348.6600 733.7000 1350.2600 734.1800 ;
        RECT 1393.6600 711.9400 1395.2600 712.4200 ;
        RECT 1393.6600 717.3800 1395.2600 717.8600 ;
        RECT 1393.6600 722.8200 1395.2600 723.3000 ;
        RECT 1393.6600 701.0600 1395.2600 701.5400 ;
        RECT 1393.6600 706.5000 1395.2600 706.9800 ;
        RECT 1348.6600 711.9400 1350.2600 712.4200 ;
        RECT 1348.6600 717.3800 1350.2600 717.8600 ;
        RECT 1348.6600 722.8200 1350.2600 723.3000 ;
        RECT 1348.6600 701.0600 1350.2600 701.5400 ;
        RECT 1348.6600 706.5000 1350.2600 706.9800 ;
        RECT 1303.6600 739.1400 1305.2600 739.6200 ;
        RECT 1303.6600 744.5800 1305.2600 745.0600 ;
        RECT 1303.6600 750.0200 1305.2600 750.5000 ;
        RECT 1295.9000 739.1400 1297.5000 739.6200 ;
        RECT 1295.9000 744.5800 1297.5000 745.0600 ;
        RECT 1295.9000 750.0200 1297.5000 750.5000 ;
        RECT 1303.6600 728.2600 1305.2600 728.7400 ;
        RECT 1303.6600 733.7000 1305.2600 734.1800 ;
        RECT 1295.9000 728.2600 1297.5000 728.7400 ;
        RECT 1295.9000 733.7000 1297.5000 734.1800 ;
        RECT 1303.6600 711.9400 1305.2600 712.4200 ;
        RECT 1303.6600 717.3800 1305.2600 717.8600 ;
        RECT 1303.6600 722.8200 1305.2600 723.3000 ;
        RECT 1295.9000 711.9400 1297.5000 712.4200 ;
        RECT 1295.9000 717.3800 1297.5000 717.8600 ;
        RECT 1295.9000 722.8200 1297.5000 723.3000 ;
        RECT 1303.6600 701.0600 1305.2600 701.5400 ;
        RECT 1303.6600 706.5000 1305.2600 706.9800 ;
        RECT 1295.9000 701.0600 1297.5000 701.5400 ;
        RECT 1295.9000 706.5000 1297.5000 706.9800 ;
        RECT 1393.6600 684.7400 1395.2600 685.2200 ;
        RECT 1393.6600 690.1800 1395.2600 690.6600 ;
        RECT 1393.6600 695.6200 1395.2600 696.1000 ;
        RECT 1393.6600 673.8600 1395.2600 674.3400 ;
        RECT 1393.6600 679.3000 1395.2600 679.7800 ;
        RECT 1348.6600 684.7400 1350.2600 685.2200 ;
        RECT 1348.6600 690.1800 1350.2600 690.6600 ;
        RECT 1348.6600 695.6200 1350.2600 696.1000 ;
        RECT 1348.6600 673.8600 1350.2600 674.3400 ;
        RECT 1348.6600 679.3000 1350.2600 679.7800 ;
        RECT 1393.6600 657.5400 1395.2600 658.0200 ;
        RECT 1393.6600 662.9800 1395.2600 663.4600 ;
        RECT 1393.6600 668.4200 1395.2600 668.9000 ;
        RECT 1393.6600 652.1000 1395.2600 652.5800 ;
        RECT 1348.6600 657.5400 1350.2600 658.0200 ;
        RECT 1348.6600 662.9800 1350.2600 663.4600 ;
        RECT 1348.6600 668.4200 1350.2600 668.9000 ;
        RECT 1348.6600 652.1000 1350.2600 652.5800 ;
        RECT 1303.6600 684.7400 1305.2600 685.2200 ;
        RECT 1303.6600 690.1800 1305.2600 690.6600 ;
        RECT 1303.6600 695.6200 1305.2600 696.1000 ;
        RECT 1295.9000 684.7400 1297.5000 685.2200 ;
        RECT 1295.9000 690.1800 1297.5000 690.6600 ;
        RECT 1295.9000 695.6200 1297.5000 696.1000 ;
        RECT 1303.6600 673.8600 1305.2600 674.3400 ;
        RECT 1303.6600 679.3000 1305.2600 679.7800 ;
        RECT 1295.9000 673.8600 1297.5000 674.3400 ;
        RECT 1295.9000 679.3000 1297.5000 679.7800 ;
        RECT 1303.6600 657.5400 1305.2600 658.0200 ;
        RECT 1303.6600 662.9800 1305.2600 663.4600 ;
        RECT 1303.6600 668.4200 1305.2600 668.9000 ;
        RECT 1295.9000 657.5400 1297.5000 658.0200 ;
        RECT 1295.9000 662.9800 1297.5000 663.4600 ;
        RECT 1295.9000 668.4200 1297.5000 668.9000 ;
        RECT 1295.9000 652.1000 1297.5000 652.5800 ;
        RECT 1303.6600 652.1000 1305.2600 652.5800 ;
        RECT 1290.3400 854.4100 1500.5600 856.0100 ;
        RECT 1290.3400 647.9100 1500.5600 649.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 642.4800 1297.5000 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 860.5200 1297.5000 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 642.4800 1495.0000 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 860.5200 1495.0000 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 647.9100 1291.9400 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 647.9100 1500.5600 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 854.4100 1291.9400 856.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 854.4100 1500.5600 856.0100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1483.6600 418.2700 1485.2600 626.3700 ;
        RECT 1438.6600 418.2700 1440.2600 626.3700 ;
        RECT 1393.6600 418.2700 1395.2600 626.3700 ;
        RECT 1348.6600 418.2700 1350.2600 626.3700 ;
        RECT 1303.6600 418.2700 1305.2600 626.3700 ;
        RECT 1493.4000 412.8400 1495.0000 632.4800 ;
        RECT 1295.9000 412.8400 1297.5000 632.4800 ;
      LAYER met3 ;
        RECT 1493.4000 607.4200 1495.0000 607.9000 ;
        RECT 1493.4000 612.8600 1495.0000 613.3400 ;
        RECT 1483.6600 607.4200 1485.2600 607.9000 ;
        RECT 1483.6600 612.8600 1485.2600 613.3400 ;
        RECT 1483.6600 618.3000 1485.2600 618.7800 ;
        RECT 1493.4000 618.3000 1495.0000 618.7800 ;
        RECT 1493.4000 596.5400 1495.0000 597.0200 ;
        RECT 1493.4000 601.9800 1495.0000 602.4600 ;
        RECT 1483.6600 596.5400 1485.2600 597.0200 ;
        RECT 1483.6600 601.9800 1485.2600 602.4600 ;
        RECT 1493.4000 580.2200 1495.0000 580.7000 ;
        RECT 1493.4000 585.6600 1495.0000 586.1400 ;
        RECT 1483.6600 580.2200 1485.2600 580.7000 ;
        RECT 1483.6600 585.6600 1485.2600 586.1400 ;
        RECT 1483.6600 591.1000 1485.2600 591.5800 ;
        RECT 1493.4000 591.1000 1495.0000 591.5800 ;
        RECT 1438.6600 607.4200 1440.2600 607.9000 ;
        RECT 1438.6600 612.8600 1440.2600 613.3400 ;
        RECT 1438.6600 618.3000 1440.2600 618.7800 ;
        RECT 1438.6600 596.5400 1440.2600 597.0200 ;
        RECT 1438.6600 601.9800 1440.2600 602.4600 ;
        RECT 1438.6600 580.2200 1440.2600 580.7000 ;
        RECT 1438.6600 585.6600 1440.2600 586.1400 ;
        RECT 1438.6600 591.1000 1440.2600 591.5800 ;
        RECT 1493.4000 563.9000 1495.0000 564.3800 ;
        RECT 1493.4000 569.3400 1495.0000 569.8200 ;
        RECT 1493.4000 574.7800 1495.0000 575.2600 ;
        RECT 1483.6600 563.9000 1485.2600 564.3800 ;
        RECT 1483.6600 569.3400 1485.2600 569.8200 ;
        RECT 1483.6600 574.7800 1485.2600 575.2600 ;
        RECT 1493.4000 553.0200 1495.0000 553.5000 ;
        RECT 1493.4000 558.4600 1495.0000 558.9400 ;
        RECT 1483.6600 553.0200 1485.2600 553.5000 ;
        RECT 1483.6600 558.4600 1485.2600 558.9400 ;
        RECT 1493.4000 536.7000 1495.0000 537.1800 ;
        RECT 1493.4000 542.1400 1495.0000 542.6200 ;
        RECT 1493.4000 547.5800 1495.0000 548.0600 ;
        RECT 1483.6600 536.7000 1485.2600 537.1800 ;
        RECT 1483.6600 542.1400 1485.2600 542.6200 ;
        RECT 1483.6600 547.5800 1485.2600 548.0600 ;
        RECT 1493.4000 525.8200 1495.0000 526.3000 ;
        RECT 1493.4000 531.2600 1495.0000 531.7400 ;
        RECT 1483.6600 525.8200 1485.2600 526.3000 ;
        RECT 1483.6600 531.2600 1485.2600 531.7400 ;
        RECT 1438.6600 563.9000 1440.2600 564.3800 ;
        RECT 1438.6600 569.3400 1440.2600 569.8200 ;
        RECT 1438.6600 574.7800 1440.2600 575.2600 ;
        RECT 1438.6600 553.0200 1440.2600 553.5000 ;
        RECT 1438.6600 558.4600 1440.2600 558.9400 ;
        RECT 1438.6600 536.7000 1440.2600 537.1800 ;
        RECT 1438.6600 542.1400 1440.2600 542.6200 ;
        RECT 1438.6600 547.5800 1440.2600 548.0600 ;
        RECT 1438.6600 525.8200 1440.2600 526.3000 ;
        RECT 1438.6600 531.2600 1440.2600 531.7400 ;
        RECT 1393.6600 607.4200 1395.2600 607.9000 ;
        RECT 1393.6600 612.8600 1395.2600 613.3400 ;
        RECT 1393.6600 618.3000 1395.2600 618.7800 ;
        RECT 1348.6600 607.4200 1350.2600 607.9000 ;
        RECT 1348.6600 612.8600 1350.2600 613.3400 ;
        RECT 1348.6600 618.3000 1350.2600 618.7800 ;
        RECT 1393.6600 596.5400 1395.2600 597.0200 ;
        RECT 1393.6600 601.9800 1395.2600 602.4600 ;
        RECT 1393.6600 580.2200 1395.2600 580.7000 ;
        RECT 1393.6600 585.6600 1395.2600 586.1400 ;
        RECT 1393.6600 591.1000 1395.2600 591.5800 ;
        RECT 1348.6600 596.5400 1350.2600 597.0200 ;
        RECT 1348.6600 601.9800 1350.2600 602.4600 ;
        RECT 1348.6600 580.2200 1350.2600 580.7000 ;
        RECT 1348.6600 585.6600 1350.2600 586.1400 ;
        RECT 1348.6600 591.1000 1350.2600 591.5800 ;
        RECT 1303.6600 607.4200 1305.2600 607.9000 ;
        RECT 1303.6600 612.8600 1305.2600 613.3400 ;
        RECT 1295.9000 607.4200 1297.5000 607.9000 ;
        RECT 1295.9000 612.8600 1297.5000 613.3400 ;
        RECT 1295.9000 618.3000 1297.5000 618.7800 ;
        RECT 1303.6600 618.3000 1305.2600 618.7800 ;
        RECT 1303.6600 596.5400 1305.2600 597.0200 ;
        RECT 1303.6600 601.9800 1305.2600 602.4600 ;
        RECT 1295.9000 596.5400 1297.5000 597.0200 ;
        RECT 1295.9000 601.9800 1297.5000 602.4600 ;
        RECT 1303.6600 580.2200 1305.2600 580.7000 ;
        RECT 1303.6600 585.6600 1305.2600 586.1400 ;
        RECT 1295.9000 580.2200 1297.5000 580.7000 ;
        RECT 1295.9000 585.6600 1297.5000 586.1400 ;
        RECT 1295.9000 591.1000 1297.5000 591.5800 ;
        RECT 1303.6600 591.1000 1305.2600 591.5800 ;
        RECT 1393.6600 563.9000 1395.2600 564.3800 ;
        RECT 1393.6600 569.3400 1395.2600 569.8200 ;
        RECT 1393.6600 574.7800 1395.2600 575.2600 ;
        RECT 1393.6600 553.0200 1395.2600 553.5000 ;
        RECT 1393.6600 558.4600 1395.2600 558.9400 ;
        RECT 1348.6600 563.9000 1350.2600 564.3800 ;
        RECT 1348.6600 569.3400 1350.2600 569.8200 ;
        RECT 1348.6600 574.7800 1350.2600 575.2600 ;
        RECT 1348.6600 553.0200 1350.2600 553.5000 ;
        RECT 1348.6600 558.4600 1350.2600 558.9400 ;
        RECT 1393.6600 536.7000 1395.2600 537.1800 ;
        RECT 1393.6600 542.1400 1395.2600 542.6200 ;
        RECT 1393.6600 547.5800 1395.2600 548.0600 ;
        RECT 1393.6600 525.8200 1395.2600 526.3000 ;
        RECT 1393.6600 531.2600 1395.2600 531.7400 ;
        RECT 1348.6600 536.7000 1350.2600 537.1800 ;
        RECT 1348.6600 542.1400 1350.2600 542.6200 ;
        RECT 1348.6600 547.5800 1350.2600 548.0600 ;
        RECT 1348.6600 525.8200 1350.2600 526.3000 ;
        RECT 1348.6600 531.2600 1350.2600 531.7400 ;
        RECT 1303.6600 563.9000 1305.2600 564.3800 ;
        RECT 1303.6600 569.3400 1305.2600 569.8200 ;
        RECT 1303.6600 574.7800 1305.2600 575.2600 ;
        RECT 1295.9000 563.9000 1297.5000 564.3800 ;
        RECT 1295.9000 569.3400 1297.5000 569.8200 ;
        RECT 1295.9000 574.7800 1297.5000 575.2600 ;
        RECT 1303.6600 553.0200 1305.2600 553.5000 ;
        RECT 1303.6600 558.4600 1305.2600 558.9400 ;
        RECT 1295.9000 553.0200 1297.5000 553.5000 ;
        RECT 1295.9000 558.4600 1297.5000 558.9400 ;
        RECT 1303.6600 536.7000 1305.2600 537.1800 ;
        RECT 1303.6600 542.1400 1305.2600 542.6200 ;
        RECT 1303.6600 547.5800 1305.2600 548.0600 ;
        RECT 1295.9000 536.7000 1297.5000 537.1800 ;
        RECT 1295.9000 542.1400 1297.5000 542.6200 ;
        RECT 1295.9000 547.5800 1297.5000 548.0600 ;
        RECT 1303.6600 525.8200 1305.2600 526.3000 ;
        RECT 1303.6600 531.2600 1305.2600 531.7400 ;
        RECT 1295.9000 525.8200 1297.5000 526.3000 ;
        RECT 1295.9000 531.2600 1297.5000 531.7400 ;
        RECT 1493.4000 509.5000 1495.0000 509.9800 ;
        RECT 1493.4000 514.9400 1495.0000 515.4200 ;
        RECT 1493.4000 520.3800 1495.0000 520.8600 ;
        RECT 1483.6600 509.5000 1485.2600 509.9800 ;
        RECT 1483.6600 514.9400 1485.2600 515.4200 ;
        RECT 1483.6600 520.3800 1485.2600 520.8600 ;
        RECT 1493.4000 498.6200 1495.0000 499.1000 ;
        RECT 1493.4000 504.0600 1495.0000 504.5400 ;
        RECT 1483.6600 498.6200 1485.2600 499.1000 ;
        RECT 1483.6600 504.0600 1485.2600 504.5400 ;
        RECT 1493.4000 482.3000 1495.0000 482.7800 ;
        RECT 1493.4000 487.7400 1495.0000 488.2200 ;
        RECT 1493.4000 493.1800 1495.0000 493.6600 ;
        RECT 1483.6600 482.3000 1485.2600 482.7800 ;
        RECT 1483.6600 487.7400 1485.2600 488.2200 ;
        RECT 1483.6600 493.1800 1485.2600 493.6600 ;
        RECT 1493.4000 471.4200 1495.0000 471.9000 ;
        RECT 1493.4000 476.8600 1495.0000 477.3400 ;
        RECT 1483.6600 471.4200 1485.2600 471.9000 ;
        RECT 1483.6600 476.8600 1485.2600 477.3400 ;
        RECT 1438.6600 509.5000 1440.2600 509.9800 ;
        RECT 1438.6600 514.9400 1440.2600 515.4200 ;
        RECT 1438.6600 520.3800 1440.2600 520.8600 ;
        RECT 1438.6600 498.6200 1440.2600 499.1000 ;
        RECT 1438.6600 504.0600 1440.2600 504.5400 ;
        RECT 1438.6600 482.3000 1440.2600 482.7800 ;
        RECT 1438.6600 487.7400 1440.2600 488.2200 ;
        RECT 1438.6600 493.1800 1440.2600 493.6600 ;
        RECT 1438.6600 471.4200 1440.2600 471.9000 ;
        RECT 1438.6600 476.8600 1440.2600 477.3400 ;
        RECT 1493.4000 455.1000 1495.0000 455.5800 ;
        RECT 1493.4000 460.5400 1495.0000 461.0200 ;
        RECT 1493.4000 465.9800 1495.0000 466.4600 ;
        RECT 1483.6600 455.1000 1485.2600 455.5800 ;
        RECT 1483.6600 460.5400 1485.2600 461.0200 ;
        RECT 1483.6600 465.9800 1485.2600 466.4600 ;
        RECT 1493.4000 444.2200 1495.0000 444.7000 ;
        RECT 1493.4000 449.6600 1495.0000 450.1400 ;
        RECT 1483.6600 444.2200 1485.2600 444.7000 ;
        RECT 1483.6600 449.6600 1485.2600 450.1400 ;
        RECT 1493.4000 427.9000 1495.0000 428.3800 ;
        RECT 1493.4000 433.3400 1495.0000 433.8200 ;
        RECT 1493.4000 438.7800 1495.0000 439.2600 ;
        RECT 1483.6600 427.9000 1485.2600 428.3800 ;
        RECT 1483.6600 433.3400 1485.2600 433.8200 ;
        RECT 1483.6600 438.7800 1485.2600 439.2600 ;
        RECT 1483.6600 422.4600 1485.2600 422.9400 ;
        RECT 1493.4000 422.4600 1495.0000 422.9400 ;
        RECT 1438.6600 455.1000 1440.2600 455.5800 ;
        RECT 1438.6600 460.5400 1440.2600 461.0200 ;
        RECT 1438.6600 465.9800 1440.2600 466.4600 ;
        RECT 1438.6600 444.2200 1440.2600 444.7000 ;
        RECT 1438.6600 449.6600 1440.2600 450.1400 ;
        RECT 1438.6600 427.9000 1440.2600 428.3800 ;
        RECT 1438.6600 433.3400 1440.2600 433.8200 ;
        RECT 1438.6600 438.7800 1440.2600 439.2600 ;
        RECT 1438.6600 422.4600 1440.2600 422.9400 ;
        RECT 1393.6600 509.5000 1395.2600 509.9800 ;
        RECT 1393.6600 514.9400 1395.2600 515.4200 ;
        RECT 1393.6600 520.3800 1395.2600 520.8600 ;
        RECT 1393.6600 498.6200 1395.2600 499.1000 ;
        RECT 1393.6600 504.0600 1395.2600 504.5400 ;
        RECT 1348.6600 509.5000 1350.2600 509.9800 ;
        RECT 1348.6600 514.9400 1350.2600 515.4200 ;
        RECT 1348.6600 520.3800 1350.2600 520.8600 ;
        RECT 1348.6600 498.6200 1350.2600 499.1000 ;
        RECT 1348.6600 504.0600 1350.2600 504.5400 ;
        RECT 1393.6600 482.3000 1395.2600 482.7800 ;
        RECT 1393.6600 487.7400 1395.2600 488.2200 ;
        RECT 1393.6600 493.1800 1395.2600 493.6600 ;
        RECT 1393.6600 471.4200 1395.2600 471.9000 ;
        RECT 1393.6600 476.8600 1395.2600 477.3400 ;
        RECT 1348.6600 482.3000 1350.2600 482.7800 ;
        RECT 1348.6600 487.7400 1350.2600 488.2200 ;
        RECT 1348.6600 493.1800 1350.2600 493.6600 ;
        RECT 1348.6600 471.4200 1350.2600 471.9000 ;
        RECT 1348.6600 476.8600 1350.2600 477.3400 ;
        RECT 1303.6600 509.5000 1305.2600 509.9800 ;
        RECT 1303.6600 514.9400 1305.2600 515.4200 ;
        RECT 1303.6600 520.3800 1305.2600 520.8600 ;
        RECT 1295.9000 509.5000 1297.5000 509.9800 ;
        RECT 1295.9000 514.9400 1297.5000 515.4200 ;
        RECT 1295.9000 520.3800 1297.5000 520.8600 ;
        RECT 1303.6600 498.6200 1305.2600 499.1000 ;
        RECT 1303.6600 504.0600 1305.2600 504.5400 ;
        RECT 1295.9000 498.6200 1297.5000 499.1000 ;
        RECT 1295.9000 504.0600 1297.5000 504.5400 ;
        RECT 1303.6600 482.3000 1305.2600 482.7800 ;
        RECT 1303.6600 487.7400 1305.2600 488.2200 ;
        RECT 1303.6600 493.1800 1305.2600 493.6600 ;
        RECT 1295.9000 482.3000 1297.5000 482.7800 ;
        RECT 1295.9000 487.7400 1297.5000 488.2200 ;
        RECT 1295.9000 493.1800 1297.5000 493.6600 ;
        RECT 1303.6600 471.4200 1305.2600 471.9000 ;
        RECT 1303.6600 476.8600 1305.2600 477.3400 ;
        RECT 1295.9000 471.4200 1297.5000 471.9000 ;
        RECT 1295.9000 476.8600 1297.5000 477.3400 ;
        RECT 1393.6600 455.1000 1395.2600 455.5800 ;
        RECT 1393.6600 460.5400 1395.2600 461.0200 ;
        RECT 1393.6600 465.9800 1395.2600 466.4600 ;
        RECT 1393.6600 444.2200 1395.2600 444.7000 ;
        RECT 1393.6600 449.6600 1395.2600 450.1400 ;
        RECT 1348.6600 455.1000 1350.2600 455.5800 ;
        RECT 1348.6600 460.5400 1350.2600 461.0200 ;
        RECT 1348.6600 465.9800 1350.2600 466.4600 ;
        RECT 1348.6600 444.2200 1350.2600 444.7000 ;
        RECT 1348.6600 449.6600 1350.2600 450.1400 ;
        RECT 1393.6600 427.9000 1395.2600 428.3800 ;
        RECT 1393.6600 433.3400 1395.2600 433.8200 ;
        RECT 1393.6600 438.7800 1395.2600 439.2600 ;
        RECT 1393.6600 422.4600 1395.2600 422.9400 ;
        RECT 1348.6600 427.9000 1350.2600 428.3800 ;
        RECT 1348.6600 433.3400 1350.2600 433.8200 ;
        RECT 1348.6600 438.7800 1350.2600 439.2600 ;
        RECT 1348.6600 422.4600 1350.2600 422.9400 ;
        RECT 1303.6600 455.1000 1305.2600 455.5800 ;
        RECT 1303.6600 460.5400 1305.2600 461.0200 ;
        RECT 1303.6600 465.9800 1305.2600 466.4600 ;
        RECT 1295.9000 455.1000 1297.5000 455.5800 ;
        RECT 1295.9000 460.5400 1297.5000 461.0200 ;
        RECT 1295.9000 465.9800 1297.5000 466.4600 ;
        RECT 1303.6600 444.2200 1305.2600 444.7000 ;
        RECT 1303.6600 449.6600 1305.2600 450.1400 ;
        RECT 1295.9000 444.2200 1297.5000 444.7000 ;
        RECT 1295.9000 449.6600 1297.5000 450.1400 ;
        RECT 1303.6600 427.9000 1305.2600 428.3800 ;
        RECT 1303.6600 433.3400 1305.2600 433.8200 ;
        RECT 1303.6600 438.7800 1305.2600 439.2600 ;
        RECT 1295.9000 427.9000 1297.5000 428.3800 ;
        RECT 1295.9000 433.3400 1297.5000 433.8200 ;
        RECT 1295.9000 438.7800 1297.5000 439.2600 ;
        RECT 1295.9000 422.4600 1297.5000 422.9400 ;
        RECT 1303.6600 422.4600 1305.2600 422.9400 ;
        RECT 1290.3400 624.7700 1500.5600 626.3700 ;
        RECT 1290.3400 418.2700 1500.5600 419.8700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 412.8400 1297.5000 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1295.9000 630.8800 1297.5000 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 412.8400 1495.0000 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.4000 630.8800 1495.0000 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 418.2700 1291.9400 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 418.2700 1500.5600 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1290.3400 624.7700 1291.9400 626.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1498.9600 624.7700 1500.5600 626.3700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1516.0200 2479.6000 1517.6200 2509.8600 ;
        RECT 1713.7200 2479.6000 1715.3200 2509.8600 ;
      LAYER met3 ;
        RECT 1713.7200 2497.3800 1715.3200 2497.8600 ;
        RECT 1516.0200 2497.3800 1517.6200 2497.8600 ;
        RECT 1713.7200 2491.9400 1715.3200 2492.4200 ;
        RECT 1713.7200 2486.5000 1715.3200 2486.9800 ;
        RECT 1516.0200 2491.9400 1517.6200 2492.4200 ;
        RECT 1516.0200 2486.5000 1517.6200 2486.9800 ;
        RECT 1510.5600 2503.1000 1720.7800 2504.7000 ;
        RECT 1510.5600 2483.5700 1720.7800 2485.1700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.0200 2479.6000 1517.6200 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.0200 2508.2600 1517.6200 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.7200 2479.6000 1715.3200 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.7200 2508.2600 1715.3200 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2483.5700 1512.1600 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2483.5700 1720.7800 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2503.1000 1512.1600 2504.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2503.1000 1720.7800 2504.7000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 188.6300 1705.4800 396.7300 ;
        RECT 1658.8800 188.6300 1660.4800 396.7300 ;
        RECT 1613.8800 188.6300 1615.4800 396.7300 ;
        RECT 1568.8800 188.6300 1570.4800 396.7300 ;
        RECT 1523.8800 188.6300 1525.4800 396.7300 ;
        RECT 1713.6200 183.2000 1715.2200 402.8400 ;
        RECT 1516.1200 183.2000 1517.7200 402.8400 ;
      LAYER met3 ;
        RECT 1713.6200 377.7800 1715.2200 378.2600 ;
        RECT 1713.6200 383.2200 1715.2200 383.7000 ;
        RECT 1703.8800 377.7800 1705.4800 378.2600 ;
        RECT 1703.8800 383.2200 1705.4800 383.7000 ;
        RECT 1703.8800 388.6600 1705.4800 389.1400 ;
        RECT 1713.6200 388.6600 1715.2200 389.1400 ;
        RECT 1713.6200 366.9000 1715.2200 367.3800 ;
        RECT 1713.6200 372.3400 1715.2200 372.8200 ;
        RECT 1703.8800 366.9000 1705.4800 367.3800 ;
        RECT 1703.8800 372.3400 1705.4800 372.8200 ;
        RECT 1713.6200 350.5800 1715.2200 351.0600 ;
        RECT 1713.6200 356.0200 1715.2200 356.5000 ;
        RECT 1703.8800 350.5800 1705.4800 351.0600 ;
        RECT 1703.8800 356.0200 1705.4800 356.5000 ;
        RECT 1703.8800 361.4600 1705.4800 361.9400 ;
        RECT 1713.6200 361.4600 1715.2200 361.9400 ;
        RECT 1658.8800 377.7800 1660.4800 378.2600 ;
        RECT 1658.8800 383.2200 1660.4800 383.7000 ;
        RECT 1658.8800 388.6600 1660.4800 389.1400 ;
        RECT 1658.8800 366.9000 1660.4800 367.3800 ;
        RECT 1658.8800 372.3400 1660.4800 372.8200 ;
        RECT 1658.8800 350.5800 1660.4800 351.0600 ;
        RECT 1658.8800 356.0200 1660.4800 356.5000 ;
        RECT 1658.8800 361.4600 1660.4800 361.9400 ;
        RECT 1713.6200 334.2600 1715.2200 334.7400 ;
        RECT 1713.6200 339.7000 1715.2200 340.1800 ;
        RECT 1713.6200 345.1400 1715.2200 345.6200 ;
        RECT 1703.8800 334.2600 1705.4800 334.7400 ;
        RECT 1703.8800 339.7000 1705.4800 340.1800 ;
        RECT 1703.8800 345.1400 1705.4800 345.6200 ;
        RECT 1713.6200 323.3800 1715.2200 323.8600 ;
        RECT 1713.6200 328.8200 1715.2200 329.3000 ;
        RECT 1703.8800 323.3800 1705.4800 323.8600 ;
        RECT 1703.8800 328.8200 1705.4800 329.3000 ;
        RECT 1713.6200 307.0600 1715.2200 307.5400 ;
        RECT 1713.6200 312.5000 1715.2200 312.9800 ;
        RECT 1713.6200 317.9400 1715.2200 318.4200 ;
        RECT 1703.8800 307.0600 1705.4800 307.5400 ;
        RECT 1703.8800 312.5000 1705.4800 312.9800 ;
        RECT 1703.8800 317.9400 1705.4800 318.4200 ;
        RECT 1713.6200 296.1800 1715.2200 296.6600 ;
        RECT 1713.6200 301.6200 1715.2200 302.1000 ;
        RECT 1703.8800 296.1800 1705.4800 296.6600 ;
        RECT 1703.8800 301.6200 1705.4800 302.1000 ;
        RECT 1658.8800 334.2600 1660.4800 334.7400 ;
        RECT 1658.8800 339.7000 1660.4800 340.1800 ;
        RECT 1658.8800 345.1400 1660.4800 345.6200 ;
        RECT 1658.8800 323.3800 1660.4800 323.8600 ;
        RECT 1658.8800 328.8200 1660.4800 329.3000 ;
        RECT 1658.8800 307.0600 1660.4800 307.5400 ;
        RECT 1658.8800 312.5000 1660.4800 312.9800 ;
        RECT 1658.8800 317.9400 1660.4800 318.4200 ;
        RECT 1658.8800 296.1800 1660.4800 296.6600 ;
        RECT 1658.8800 301.6200 1660.4800 302.1000 ;
        RECT 1613.8800 377.7800 1615.4800 378.2600 ;
        RECT 1613.8800 383.2200 1615.4800 383.7000 ;
        RECT 1613.8800 388.6600 1615.4800 389.1400 ;
        RECT 1568.8800 377.7800 1570.4800 378.2600 ;
        RECT 1568.8800 383.2200 1570.4800 383.7000 ;
        RECT 1568.8800 388.6600 1570.4800 389.1400 ;
        RECT 1613.8800 366.9000 1615.4800 367.3800 ;
        RECT 1613.8800 372.3400 1615.4800 372.8200 ;
        RECT 1613.8800 350.5800 1615.4800 351.0600 ;
        RECT 1613.8800 356.0200 1615.4800 356.5000 ;
        RECT 1613.8800 361.4600 1615.4800 361.9400 ;
        RECT 1568.8800 366.9000 1570.4800 367.3800 ;
        RECT 1568.8800 372.3400 1570.4800 372.8200 ;
        RECT 1568.8800 350.5800 1570.4800 351.0600 ;
        RECT 1568.8800 356.0200 1570.4800 356.5000 ;
        RECT 1568.8800 361.4600 1570.4800 361.9400 ;
        RECT 1523.8800 377.7800 1525.4800 378.2600 ;
        RECT 1523.8800 383.2200 1525.4800 383.7000 ;
        RECT 1516.1200 377.7800 1517.7200 378.2600 ;
        RECT 1516.1200 383.2200 1517.7200 383.7000 ;
        RECT 1516.1200 388.6600 1517.7200 389.1400 ;
        RECT 1523.8800 388.6600 1525.4800 389.1400 ;
        RECT 1523.8800 366.9000 1525.4800 367.3800 ;
        RECT 1523.8800 372.3400 1525.4800 372.8200 ;
        RECT 1516.1200 366.9000 1517.7200 367.3800 ;
        RECT 1516.1200 372.3400 1517.7200 372.8200 ;
        RECT 1523.8800 350.5800 1525.4800 351.0600 ;
        RECT 1523.8800 356.0200 1525.4800 356.5000 ;
        RECT 1516.1200 350.5800 1517.7200 351.0600 ;
        RECT 1516.1200 356.0200 1517.7200 356.5000 ;
        RECT 1516.1200 361.4600 1517.7200 361.9400 ;
        RECT 1523.8800 361.4600 1525.4800 361.9400 ;
        RECT 1613.8800 334.2600 1615.4800 334.7400 ;
        RECT 1613.8800 339.7000 1615.4800 340.1800 ;
        RECT 1613.8800 345.1400 1615.4800 345.6200 ;
        RECT 1613.8800 323.3800 1615.4800 323.8600 ;
        RECT 1613.8800 328.8200 1615.4800 329.3000 ;
        RECT 1568.8800 334.2600 1570.4800 334.7400 ;
        RECT 1568.8800 339.7000 1570.4800 340.1800 ;
        RECT 1568.8800 345.1400 1570.4800 345.6200 ;
        RECT 1568.8800 323.3800 1570.4800 323.8600 ;
        RECT 1568.8800 328.8200 1570.4800 329.3000 ;
        RECT 1613.8800 307.0600 1615.4800 307.5400 ;
        RECT 1613.8800 312.5000 1615.4800 312.9800 ;
        RECT 1613.8800 317.9400 1615.4800 318.4200 ;
        RECT 1613.8800 296.1800 1615.4800 296.6600 ;
        RECT 1613.8800 301.6200 1615.4800 302.1000 ;
        RECT 1568.8800 307.0600 1570.4800 307.5400 ;
        RECT 1568.8800 312.5000 1570.4800 312.9800 ;
        RECT 1568.8800 317.9400 1570.4800 318.4200 ;
        RECT 1568.8800 296.1800 1570.4800 296.6600 ;
        RECT 1568.8800 301.6200 1570.4800 302.1000 ;
        RECT 1523.8800 334.2600 1525.4800 334.7400 ;
        RECT 1523.8800 339.7000 1525.4800 340.1800 ;
        RECT 1523.8800 345.1400 1525.4800 345.6200 ;
        RECT 1516.1200 334.2600 1517.7200 334.7400 ;
        RECT 1516.1200 339.7000 1517.7200 340.1800 ;
        RECT 1516.1200 345.1400 1517.7200 345.6200 ;
        RECT 1523.8800 323.3800 1525.4800 323.8600 ;
        RECT 1523.8800 328.8200 1525.4800 329.3000 ;
        RECT 1516.1200 323.3800 1517.7200 323.8600 ;
        RECT 1516.1200 328.8200 1517.7200 329.3000 ;
        RECT 1523.8800 307.0600 1525.4800 307.5400 ;
        RECT 1523.8800 312.5000 1525.4800 312.9800 ;
        RECT 1523.8800 317.9400 1525.4800 318.4200 ;
        RECT 1516.1200 307.0600 1517.7200 307.5400 ;
        RECT 1516.1200 312.5000 1517.7200 312.9800 ;
        RECT 1516.1200 317.9400 1517.7200 318.4200 ;
        RECT 1523.8800 296.1800 1525.4800 296.6600 ;
        RECT 1523.8800 301.6200 1525.4800 302.1000 ;
        RECT 1516.1200 296.1800 1517.7200 296.6600 ;
        RECT 1516.1200 301.6200 1517.7200 302.1000 ;
        RECT 1713.6200 279.8600 1715.2200 280.3400 ;
        RECT 1713.6200 285.3000 1715.2200 285.7800 ;
        RECT 1713.6200 290.7400 1715.2200 291.2200 ;
        RECT 1703.8800 279.8600 1705.4800 280.3400 ;
        RECT 1703.8800 285.3000 1705.4800 285.7800 ;
        RECT 1703.8800 290.7400 1705.4800 291.2200 ;
        RECT 1713.6200 268.9800 1715.2200 269.4600 ;
        RECT 1713.6200 274.4200 1715.2200 274.9000 ;
        RECT 1703.8800 268.9800 1705.4800 269.4600 ;
        RECT 1703.8800 274.4200 1705.4800 274.9000 ;
        RECT 1713.6200 252.6600 1715.2200 253.1400 ;
        RECT 1713.6200 258.1000 1715.2200 258.5800 ;
        RECT 1713.6200 263.5400 1715.2200 264.0200 ;
        RECT 1703.8800 252.6600 1705.4800 253.1400 ;
        RECT 1703.8800 258.1000 1705.4800 258.5800 ;
        RECT 1703.8800 263.5400 1705.4800 264.0200 ;
        RECT 1713.6200 241.7800 1715.2200 242.2600 ;
        RECT 1713.6200 247.2200 1715.2200 247.7000 ;
        RECT 1703.8800 241.7800 1705.4800 242.2600 ;
        RECT 1703.8800 247.2200 1705.4800 247.7000 ;
        RECT 1658.8800 279.8600 1660.4800 280.3400 ;
        RECT 1658.8800 285.3000 1660.4800 285.7800 ;
        RECT 1658.8800 290.7400 1660.4800 291.2200 ;
        RECT 1658.8800 268.9800 1660.4800 269.4600 ;
        RECT 1658.8800 274.4200 1660.4800 274.9000 ;
        RECT 1658.8800 252.6600 1660.4800 253.1400 ;
        RECT 1658.8800 258.1000 1660.4800 258.5800 ;
        RECT 1658.8800 263.5400 1660.4800 264.0200 ;
        RECT 1658.8800 241.7800 1660.4800 242.2600 ;
        RECT 1658.8800 247.2200 1660.4800 247.7000 ;
        RECT 1713.6200 225.4600 1715.2200 225.9400 ;
        RECT 1713.6200 230.9000 1715.2200 231.3800 ;
        RECT 1713.6200 236.3400 1715.2200 236.8200 ;
        RECT 1703.8800 225.4600 1705.4800 225.9400 ;
        RECT 1703.8800 230.9000 1705.4800 231.3800 ;
        RECT 1703.8800 236.3400 1705.4800 236.8200 ;
        RECT 1713.6200 214.5800 1715.2200 215.0600 ;
        RECT 1713.6200 220.0200 1715.2200 220.5000 ;
        RECT 1703.8800 214.5800 1705.4800 215.0600 ;
        RECT 1703.8800 220.0200 1705.4800 220.5000 ;
        RECT 1713.6200 198.2600 1715.2200 198.7400 ;
        RECT 1713.6200 203.7000 1715.2200 204.1800 ;
        RECT 1713.6200 209.1400 1715.2200 209.6200 ;
        RECT 1703.8800 198.2600 1705.4800 198.7400 ;
        RECT 1703.8800 203.7000 1705.4800 204.1800 ;
        RECT 1703.8800 209.1400 1705.4800 209.6200 ;
        RECT 1703.8800 192.8200 1705.4800 193.3000 ;
        RECT 1713.6200 192.8200 1715.2200 193.3000 ;
        RECT 1658.8800 225.4600 1660.4800 225.9400 ;
        RECT 1658.8800 230.9000 1660.4800 231.3800 ;
        RECT 1658.8800 236.3400 1660.4800 236.8200 ;
        RECT 1658.8800 214.5800 1660.4800 215.0600 ;
        RECT 1658.8800 220.0200 1660.4800 220.5000 ;
        RECT 1658.8800 198.2600 1660.4800 198.7400 ;
        RECT 1658.8800 203.7000 1660.4800 204.1800 ;
        RECT 1658.8800 209.1400 1660.4800 209.6200 ;
        RECT 1658.8800 192.8200 1660.4800 193.3000 ;
        RECT 1613.8800 279.8600 1615.4800 280.3400 ;
        RECT 1613.8800 285.3000 1615.4800 285.7800 ;
        RECT 1613.8800 290.7400 1615.4800 291.2200 ;
        RECT 1613.8800 268.9800 1615.4800 269.4600 ;
        RECT 1613.8800 274.4200 1615.4800 274.9000 ;
        RECT 1568.8800 279.8600 1570.4800 280.3400 ;
        RECT 1568.8800 285.3000 1570.4800 285.7800 ;
        RECT 1568.8800 290.7400 1570.4800 291.2200 ;
        RECT 1568.8800 268.9800 1570.4800 269.4600 ;
        RECT 1568.8800 274.4200 1570.4800 274.9000 ;
        RECT 1613.8800 252.6600 1615.4800 253.1400 ;
        RECT 1613.8800 258.1000 1615.4800 258.5800 ;
        RECT 1613.8800 263.5400 1615.4800 264.0200 ;
        RECT 1613.8800 241.7800 1615.4800 242.2600 ;
        RECT 1613.8800 247.2200 1615.4800 247.7000 ;
        RECT 1568.8800 252.6600 1570.4800 253.1400 ;
        RECT 1568.8800 258.1000 1570.4800 258.5800 ;
        RECT 1568.8800 263.5400 1570.4800 264.0200 ;
        RECT 1568.8800 241.7800 1570.4800 242.2600 ;
        RECT 1568.8800 247.2200 1570.4800 247.7000 ;
        RECT 1523.8800 279.8600 1525.4800 280.3400 ;
        RECT 1523.8800 285.3000 1525.4800 285.7800 ;
        RECT 1523.8800 290.7400 1525.4800 291.2200 ;
        RECT 1516.1200 279.8600 1517.7200 280.3400 ;
        RECT 1516.1200 285.3000 1517.7200 285.7800 ;
        RECT 1516.1200 290.7400 1517.7200 291.2200 ;
        RECT 1523.8800 268.9800 1525.4800 269.4600 ;
        RECT 1523.8800 274.4200 1525.4800 274.9000 ;
        RECT 1516.1200 268.9800 1517.7200 269.4600 ;
        RECT 1516.1200 274.4200 1517.7200 274.9000 ;
        RECT 1523.8800 252.6600 1525.4800 253.1400 ;
        RECT 1523.8800 258.1000 1525.4800 258.5800 ;
        RECT 1523.8800 263.5400 1525.4800 264.0200 ;
        RECT 1516.1200 252.6600 1517.7200 253.1400 ;
        RECT 1516.1200 258.1000 1517.7200 258.5800 ;
        RECT 1516.1200 263.5400 1517.7200 264.0200 ;
        RECT 1523.8800 241.7800 1525.4800 242.2600 ;
        RECT 1523.8800 247.2200 1525.4800 247.7000 ;
        RECT 1516.1200 241.7800 1517.7200 242.2600 ;
        RECT 1516.1200 247.2200 1517.7200 247.7000 ;
        RECT 1613.8800 225.4600 1615.4800 225.9400 ;
        RECT 1613.8800 230.9000 1615.4800 231.3800 ;
        RECT 1613.8800 236.3400 1615.4800 236.8200 ;
        RECT 1613.8800 214.5800 1615.4800 215.0600 ;
        RECT 1613.8800 220.0200 1615.4800 220.5000 ;
        RECT 1568.8800 225.4600 1570.4800 225.9400 ;
        RECT 1568.8800 230.9000 1570.4800 231.3800 ;
        RECT 1568.8800 236.3400 1570.4800 236.8200 ;
        RECT 1568.8800 214.5800 1570.4800 215.0600 ;
        RECT 1568.8800 220.0200 1570.4800 220.5000 ;
        RECT 1613.8800 198.2600 1615.4800 198.7400 ;
        RECT 1613.8800 203.7000 1615.4800 204.1800 ;
        RECT 1613.8800 209.1400 1615.4800 209.6200 ;
        RECT 1613.8800 192.8200 1615.4800 193.3000 ;
        RECT 1568.8800 198.2600 1570.4800 198.7400 ;
        RECT 1568.8800 203.7000 1570.4800 204.1800 ;
        RECT 1568.8800 209.1400 1570.4800 209.6200 ;
        RECT 1568.8800 192.8200 1570.4800 193.3000 ;
        RECT 1523.8800 225.4600 1525.4800 225.9400 ;
        RECT 1523.8800 230.9000 1525.4800 231.3800 ;
        RECT 1523.8800 236.3400 1525.4800 236.8200 ;
        RECT 1516.1200 225.4600 1517.7200 225.9400 ;
        RECT 1516.1200 230.9000 1517.7200 231.3800 ;
        RECT 1516.1200 236.3400 1517.7200 236.8200 ;
        RECT 1523.8800 214.5800 1525.4800 215.0600 ;
        RECT 1523.8800 220.0200 1525.4800 220.5000 ;
        RECT 1516.1200 214.5800 1517.7200 215.0600 ;
        RECT 1516.1200 220.0200 1517.7200 220.5000 ;
        RECT 1523.8800 198.2600 1525.4800 198.7400 ;
        RECT 1523.8800 203.7000 1525.4800 204.1800 ;
        RECT 1523.8800 209.1400 1525.4800 209.6200 ;
        RECT 1516.1200 198.2600 1517.7200 198.7400 ;
        RECT 1516.1200 203.7000 1517.7200 204.1800 ;
        RECT 1516.1200 209.1400 1517.7200 209.6200 ;
        RECT 1516.1200 192.8200 1517.7200 193.3000 ;
        RECT 1523.8800 192.8200 1525.4800 193.3000 ;
        RECT 1510.5600 395.1300 1720.7800 396.7300 ;
        RECT 1510.5600 188.6300 1720.7800 190.2300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 183.2000 1517.7200 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 401.2400 1517.7200 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 183.2000 1715.2200 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 401.2400 1715.2200 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 188.6300 1512.1600 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 188.6300 1720.7800 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 395.1300 1512.1600 396.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 395.1300 1720.7800 396.7300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1516.0200 142.9400 1517.6200 173.2000 ;
        RECT 1713.7200 142.9400 1715.3200 173.2000 ;
      LAYER met3 ;
        RECT 1713.7200 160.7200 1715.3200 161.2000 ;
        RECT 1516.0200 160.7200 1517.6200 161.2000 ;
        RECT 1713.7200 155.2800 1715.3200 155.7600 ;
        RECT 1713.7200 149.8400 1715.3200 150.3200 ;
        RECT 1516.0200 155.2800 1517.6200 155.7600 ;
        RECT 1516.0200 149.8400 1517.6200 150.3200 ;
        RECT 1510.5600 166.4400 1720.7800 168.0400 ;
        RECT 1510.5600 146.9100 1720.7800 148.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.0200 142.9400 1517.6200 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.0200 171.6000 1517.6200 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.7200 142.9400 1715.3200 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.7200 171.6000 1715.3200 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 146.9100 1512.1600 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 146.9100 1720.7800 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 166.4400 1512.1600 168.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 166.4400 1720.7800 168.0400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 2255.3900 1705.4800 2463.4900 ;
        RECT 1658.8800 2255.3900 1660.4800 2463.4900 ;
        RECT 1613.8800 2255.3900 1615.4800 2463.4900 ;
        RECT 1568.8800 2255.3900 1570.4800 2463.4900 ;
        RECT 1523.8800 2255.3900 1525.4800 2463.4900 ;
        RECT 1713.6200 2249.9600 1715.2200 2469.6000 ;
        RECT 1516.1200 2249.9600 1517.7200 2469.6000 ;
      LAYER met3 ;
        RECT 1713.6200 2444.5400 1715.2200 2445.0200 ;
        RECT 1713.6200 2449.9800 1715.2200 2450.4600 ;
        RECT 1703.8800 2444.5400 1705.4800 2445.0200 ;
        RECT 1703.8800 2449.9800 1705.4800 2450.4600 ;
        RECT 1703.8800 2455.4200 1705.4800 2455.9000 ;
        RECT 1713.6200 2455.4200 1715.2200 2455.9000 ;
        RECT 1713.6200 2433.6600 1715.2200 2434.1400 ;
        RECT 1713.6200 2439.1000 1715.2200 2439.5800 ;
        RECT 1703.8800 2433.6600 1705.4800 2434.1400 ;
        RECT 1703.8800 2439.1000 1705.4800 2439.5800 ;
        RECT 1713.6200 2417.3400 1715.2200 2417.8200 ;
        RECT 1713.6200 2422.7800 1715.2200 2423.2600 ;
        RECT 1703.8800 2417.3400 1705.4800 2417.8200 ;
        RECT 1703.8800 2422.7800 1705.4800 2423.2600 ;
        RECT 1703.8800 2428.2200 1705.4800 2428.7000 ;
        RECT 1713.6200 2428.2200 1715.2200 2428.7000 ;
        RECT 1658.8800 2444.5400 1660.4800 2445.0200 ;
        RECT 1658.8800 2449.9800 1660.4800 2450.4600 ;
        RECT 1658.8800 2455.4200 1660.4800 2455.9000 ;
        RECT 1658.8800 2433.6600 1660.4800 2434.1400 ;
        RECT 1658.8800 2439.1000 1660.4800 2439.5800 ;
        RECT 1658.8800 2417.3400 1660.4800 2417.8200 ;
        RECT 1658.8800 2422.7800 1660.4800 2423.2600 ;
        RECT 1658.8800 2428.2200 1660.4800 2428.7000 ;
        RECT 1713.6200 2401.0200 1715.2200 2401.5000 ;
        RECT 1713.6200 2406.4600 1715.2200 2406.9400 ;
        RECT 1713.6200 2411.9000 1715.2200 2412.3800 ;
        RECT 1703.8800 2401.0200 1705.4800 2401.5000 ;
        RECT 1703.8800 2406.4600 1705.4800 2406.9400 ;
        RECT 1703.8800 2411.9000 1705.4800 2412.3800 ;
        RECT 1713.6200 2390.1400 1715.2200 2390.6200 ;
        RECT 1713.6200 2395.5800 1715.2200 2396.0600 ;
        RECT 1703.8800 2390.1400 1705.4800 2390.6200 ;
        RECT 1703.8800 2395.5800 1705.4800 2396.0600 ;
        RECT 1713.6200 2373.8200 1715.2200 2374.3000 ;
        RECT 1713.6200 2379.2600 1715.2200 2379.7400 ;
        RECT 1713.6200 2384.7000 1715.2200 2385.1800 ;
        RECT 1703.8800 2373.8200 1705.4800 2374.3000 ;
        RECT 1703.8800 2379.2600 1705.4800 2379.7400 ;
        RECT 1703.8800 2384.7000 1705.4800 2385.1800 ;
        RECT 1713.6200 2362.9400 1715.2200 2363.4200 ;
        RECT 1713.6200 2368.3800 1715.2200 2368.8600 ;
        RECT 1703.8800 2362.9400 1705.4800 2363.4200 ;
        RECT 1703.8800 2368.3800 1705.4800 2368.8600 ;
        RECT 1658.8800 2401.0200 1660.4800 2401.5000 ;
        RECT 1658.8800 2406.4600 1660.4800 2406.9400 ;
        RECT 1658.8800 2411.9000 1660.4800 2412.3800 ;
        RECT 1658.8800 2390.1400 1660.4800 2390.6200 ;
        RECT 1658.8800 2395.5800 1660.4800 2396.0600 ;
        RECT 1658.8800 2373.8200 1660.4800 2374.3000 ;
        RECT 1658.8800 2379.2600 1660.4800 2379.7400 ;
        RECT 1658.8800 2384.7000 1660.4800 2385.1800 ;
        RECT 1658.8800 2362.9400 1660.4800 2363.4200 ;
        RECT 1658.8800 2368.3800 1660.4800 2368.8600 ;
        RECT 1613.8800 2444.5400 1615.4800 2445.0200 ;
        RECT 1613.8800 2449.9800 1615.4800 2450.4600 ;
        RECT 1613.8800 2455.4200 1615.4800 2455.9000 ;
        RECT 1568.8800 2444.5400 1570.4800 2445.0200 ;
        RECT 1568.8800 2449.9800 1570.4800 2450.4600 ;
        RECT 1568.8800 2455.4200 1570.4800 2455.9000 ;
        RECT 1613.8800 2433.6600 1615.4800 2434.1400 ;
        RECT 1613.8800 2439.1000 1615.4800 2439.5800 ;
        RECT 1613.8800 2417.3400 1615.4800 2417.8200 ;
        RECT 1613.8800 2422.7800 1615.4800 2423.2600 ;
        RECT 1613.8800 2428.2200 1615.4800 2428.7000 ;
        RECT 1568.8800 2433.6600 1570.4800 2434.1400 ;
        RECT 1568.8800 2439.1000 1570.4800 2439.5800 ;
        RECT 1568.8800 2417.3400 1570.4800 2417.8200 ;
        RECT 1568.8800 2422.7800 1570.4800 2423.2600 ;
        RECT 1568.8800 2428.2200 1570.4800 2428.7000 ;
        RECT 1523.8800 2444.5400 1525.4800 2445.0200 ;
        RECT 1523.8800 2449.9800 1525.4800 2450.4600 ;
        RECT 1516.1200 2444.5400 1517.7200 2445.0200 ;
        RECT 1516.1200 2449.9800 1517.7200 2450.4600 ;
        RECT 1516.1200 2455.4200 1517.7200 2455.9000 ;
        RECT 1523.8800 2455.4200 1525.4800 2455.9000 ;
        RECT 1523.8800 2433.6600 1525.4800 2434.1400 ;
        RECT 1523.8800 2439.1000 1525.4800 2439.5800 ;
        RECT 1516.1200 2433.6600 1517.7200 2434.1400 ;
        RECT 1516.1200 2439.1000 1517.7200 2439.5800 ;
        RECT 1523.8800 2417.3400 1525.4800 2417.8200 ;
        RECT 1523.8800 2422.7800 1525.4800 2423.2600 ;
        RECT 1516.1200 2417.3400 1517.7200 2417.8200 ;
        RECT 1516.1200 2422.7800 1517.7200 2423.2600 ;
        RECT 1516.1200 2428.2200 1517.7200 2428.7000 ;
        RECT 1523.8800 2428.2200 1525.4800 2428.7000 ;
        RECT 1613.8800 2401.0200 1615.4800 2401.5000 ;
        RECT 1613.8800 2406.4600 1615.4800 2406.9400 ;
        RECT 1613.8800 2411.9000 1615.4800 2412.3800 ;
        RECT 1613.8800 2390.1400 1615.4800 2390.6200 ;
        RECT 1613.8800 2395.5800 1615.4800 2396.0600 ;
        RECT 1568.8800 2401.0200 1570.4800 2401.5000 ;
        RECT 1568.8800 2406.4600 1570.4800 2406.9400 ;
        RECT 1568.8800 2411.9000 1570.4800 2412.3800 ;
        RECT 1568.8800 2390.1400 1570.4800 2390.6200 ;
        RECT 1568.8800 2395.5800 1570.4800 2396.0600 ;
        RECT 1613.8800 2373.8200 1615.4800 2374.3000 ;
        RECT 1613.8800 2379.2600 1615.4800 2379.7400 ;
        RECT 1613.8800 2384.7000 1615.4800 2385.1800 ;
        RECT 1613.8800 2362.9400 1615.4800 2363.4200 ;
        RECT 1613.8800 2368.3800 1615.4800 2368.8600 ;
        RECT 1568.8800 2373.8200 1570.4800 2374.3000 ;
        RECT 1568.8800 2379.2600 1570.4800 2379.7400 ;
        RECT 1568.8800 2384.7000 1570.4800 2385.1800 ;
        RECT 1568.8800 2362.9400 1570.4800 2363.4200 ;
        RECT 1568.8800 2368.3800 1570.4800 2368.8600 ;
        RECT 1523.8800 2401.0200 1525.4800 2401.5000 ;
        RECT 1523.8800 2406.4600 1525.4800 2406.9400 ;
        RECT 1523.8800 2411.9000 1525.4800 2412.3800 ;
        RECT 1516.1200 2401.0200 1517.7200 2401.5000 ;
        RECT 1516.1200 2406.4600 1517.7200 2406.9400 ;
        RECT 1516.1200 2411.9000 1517.7200 2412.3800 ;
        RECT 1523.8800 2390.1400 1525.4800 2390.6200 ;
        RECT 1523.8800 2395.5800 1525.4800 2396.0600 ;
        RECT 1516.1200 2390.1400 1517.7200 2390.6200 ;
        RECT 1516.1200 2395.5800 1517.7200 2396.0600 ;
        RECT 1523.8800 2373.8200 1525.4800 2374.3000 ;
        RECT 1523.8800 2379.2600 1525.4800 2379.7400 ;
        RECT 1523.8800 2384.7000 1525.4800 2385.1800 ;
        RECT 1516.1200 2373.8200 1517.7200 2374.3000 ;
        RECT 1516.1200 2379.2600 1517.7200 2379.7400 ;
        RECT 1516.1200 2384.7000 1517.7200 2385.1800 ;
        RECT 1523.8800 2362.9400 1525.4800 2363.4200 ;
        RECT 1523.8800 2368.3800 1525.4800 2368.8600 ;
        RECT 1516.1200 2362.9400 1517.7200 2363.4200 ;
        RECT 1516.1200 2368.3800 1517.7200 2368.8600 ;
        RECT 1713.6200 2346.6200 1715.2200 2347.1000 ;
        RECT 1713.6200 2352.0600 1715.2200 2352.5400 ;
        RECT 1713.6200 2357.5000 1715.2200 2357.9800 ;
        RECT 1703.8800 2346.6200 1705.4800 2347.1000 ;
        RECT 1703.8800 2352.0600 1705.4800 2352.5400 ;
        RECT 1703.8800 2357.5000 1705.4800 2357.9800 ;
        RECT 1713.6200 2335.7400 1715.2200 2336.2200 ;
        RECT 1713.6200 2341.1800 1715.2200 2341.6600 ;
        RECT 1703.8800 2335.7400 1705.4800 2336.2200 ;
        RECT 1703.8800 2341.1800 1705.4800 2341.6600 ;
        RECT 1713.6200 2319.4200 1715.2200 2319.9000 ;
        RECT 1713.6200 2324.8600 1715.2200 2325.3400 ;
        RECT 1713.6200 2330.3000 1715.2200 2330.7800 ;
        RECT 1703.8800 2319.4200 1705.4800 2319.9000 ;
        RECT 1703.8800 2324.8600 1705.4800 2325.3400 ;
        RECT 1703.8800 2330.3000 1705.4800 2330.7800 ;
        RECT 1713.6200 2308.5400 1715.2200 2309.0200 ;
        RECT 1713.6200 2313.9800 1715.2200 2314.4600 ;
        RECT 1703.8800 2308.5400 1705.4800 2309.0200 ;
        RECT 1703.8800 2313.9800 1705.4800 2314.4600 ;
        RECT 1658.8800 2346.6200 1660.4800 2347.1000 ;
        RECT 1658.8800 2352.0600 1660.4800 2352.5400 ;
        RECT 1658.8800 2357.5000 1660.4800 2357.9800 ;
        RECT 1658.8800 2335.7400 1660.4800 2336.2200 ;
        RECT 1658.8800 2341.1800 1660.4800 2341.6600 ;
        RECT 1658.8800 2319.4200 1660.4800 2319.9000 ;
        RECT 1658.8800 2324.8600 1660.4800 2325.3400 ;
        RECT 1658.8800 2330.3000 1660.4800 2330.7800 ;
        RECT 1658.8800 2308.5400 1660.4800 2309.0200 ;
        RECT 1658.8800 2313.9800 1660.4800 2314.4600 ;
        RECT 1713.6200 2292.2200 1715.2200 2292.7000 ;
        RECT 1713.6200 2297.6600 1715.2200 2298.1400 ;
        RECT 1713.6200 2303.1000 1715.2200 2303.5800 ;
        RECT 1703.8800 2292.2200 1705.4800 2292.7000 ;
        RECT 1703.8800 2297.6600 1705.4800 2298.1400 ;
        RECT 1703.8800 2303.1000 1705.4800 2303.5800 ;
        RECT 1713.6200 2281.3400 1715.2200 2281.8200 ;
        RECT 1713.6200 2286.7800 1715.2200 2287.2600 ;
        RECT 1703.8800 2281.3400 1705.4800 2281.8200 ;
        RECT 1703.8800 2286.7800 1705.4800 2287.2600 ;
        RECT 1713.6200 2265.0200 1715.2200 2265.5000 ;
        RECT 1713.6200 2270.4600 1715.2200 2270.9400 ;
        RECT 1713.6200 2275.9000 1715.2200 2276.3800 ;
        RECT 1703.8800 2265.0200 1705.4800 2265.5000 ;
        RECT 1703.8800 2270.4600 1705.4800 2270.9400 ;
        RECT 1703.8800 2275.9000 1705.4800 2276.3800 ;
        RECT 1703.8800 2259.5800 1705.4800 2260.0600 ;
        RECT 1713.6200 2259.5800 1715.2200 2260.0600 ;
        RECT 1658.8800 2292.2200 1660.4800 2292.7000 ;
        RECT 1658.8800 2297.6600 1660.4800 2298.1400 ;
        RECT 1658.8800 2303.1000 1660.4800 2303.5800 ;
        RECT 1658.8800 2281.3400 1660.4800 2281.8200 ;
        RECT 1658.8800 2286.7800 1660.4800 2287.2600 ;
        RECT 1658.8800 2265.0200 1660.4800 2265.5000 ;
        RECT 1658.8800 2270.4600 1660.4800 2270.9400 ;
        RECT 1658.8800 2275.9000 1660.4800 2276.3800 ;
        RECT 1658.8800 2259.5800 1660.4800 2260.0600 ;
        RECT 1613.8800 2346.6200 1615.4800 2347.1000 ;
        RECT 1613.8800 2352.0600 1615.4800 2352.5400 ;
        RECT 1613.8800 2357.5000 1615.4800 2357.9800 ;
        RECT 1613.8800 2335.7400 1615.4800 2336.2200 ;
        RECT 1613.8800 2341.1800 1615.4800 2341.6600 ;
        RECT 1568.8800 2346.6200 1570.4800 2347.1000 ;
        RECT 1568.8800 2352.0600 1570.4800 2352.5400 ;
        RECT 1568.8800 2357.5000 1570.4800 2357.9800 ;
        RECT 1568.8800 2335.7400 1570.4800 2336.2200 ;
        RECT 1568.8800 2341.1800 1570.4800 2341.6600 ;
        RECT 1613.8800 2319.4200 1615.4800 2319.9000 ;
        RECT 1613.8800 2324.8600 1615.4800 2325.3400 ;
        RECT 1613.8800 2330.3000 1615.4800 2330.7800 ;
        RECT 1613.8800 2308.5400 1615.4800 2309.0200 ;
        RECT 1613.8800 2313.9800 1615.4800 2314.4600 ;
        RECT 1568.8800 2319.4200 1570.4800 2319.9000 ;
        RECT 1568.8800 2324.8600 1570.4800 2325.3400 ;
        RECT 1568.8800 2330.3000 1570.4800 2330.7800 ;
        RECT 1568.8800 2308.5400 1570.4800 2309.0200 ;
        RECT 1568.8800 2313.9800 1570.4800 2314.4600 ;
        RECT 1523.8800 2346.6200 1525.4800 2347.1000 ;
        RECT 1523.8800 2352.0600 1525.4800 2352.5400 ;
        RECT 1523.8800 2357.5000 1525.4800 2357.9800 ;
        RECT 1516.1200 2346.6200 1517.7200 2347.1000 ;
        RECT 1516.1200 2352.0600 1517.7200 2352.5400 ;
        RECT 1516.1200 2357.5000 1517.7200 2357.9800 ;
        RECT 1523.8800 2335.7400 1525.4800 2336.2200 ;
        RECT 1523.8800 2341.1800 1525.4800 2341.6600 ;
        RECT 1516.1200 2335.7400 1517.7200 2336.2200 ;
        RECT 1516.1200 2341.1800 1517.7200 2341.6600 ;
        RECT 1523.8800 2319.4200 1525.4800 2319.9000 ;
        RECT 1523.8800 2324.8600 1525.4800 2325.3400 ;
        RECT 1523.8800 2330.3000 1525.4800 2330.7800 ;
        RECT 1516.1200 2319.4200 1517.7200 2319.9000 ;
        RECT 1516.1200 2324.8600 1517.7200 2325.3400 ;
        RECT 1516.1200 2330.3000 1517.7200 2330.7800 ;
        RECT 1523.8800 2308.5400 1525.4800 2309.0200 ;
        RECT 1523.8800 2313.9800 1525.4800 2314.4600 ;
        RECT 1516.1200 2308.5400 1517.7200 2309.0200 ;
        RECT 1516.1200 2313.9800 1517.7200 2314.4600 ;
        RECT 1613.8800 2292.2200 1615.4800 2292.7000 ;
        RECT 1613.8800 2297.6600 1615.4800 2298.1400 ;
        RECT 1613.8800 2303.1000 1615.4800 2303.5800 ;
        RECT 1613.8800 2281.3400 1615.4800 2281.8200 ;
        RECT 1613.8800 2286.7800 1615.4800 2287.2600 ;
        RECT 1568.8800 2292.2200 1570.4800 2292.7000 ;
        RECT 1568.8800 2297.6600 1570.4800 2298.1400 ;
        RECT 1568.8800 2303.1000 1570.4800 2303.5800 ;
        RECT 1568.8800 2281.3400 1570.4800 2281.8200 ;
        RECT 1568.8800 2286.7800 1570.4800 2287.2600 ;
        RECT 1613.8800 2265.0200 1615.4800 2265.5000 ;
        RECT 1613.8800 2270.4600 1615.4800 2270.9400 ;
        RECT 1613.8800 2275.9000 1615.4800 2276.3800 ;
        RECT 1613.8800 2259.5800 1615.4800 2260.0600 ;
        RECT 1568.8800 2265.0200 1570.4800 2265.5000 ;
        RECT 1568.8800 2270.4600 1570.4800 2270.9400 ;
        RECT 1568.8800 2275.9000 1570.4800 2276.3800 ;
        RECT 1568.8800 2259.5800 1570.4800 2260.0600 ;
        RECT 1523.8800 2292.2200 1525.4800 2292.7000 ;
        RECT 1523.8800 2297.6600 1525.4800 2298.1400 ;
        RECT 1523.8800 2303.1000 1525.4800 2303.5800 ;
        RECT 1516.1200 2292.2200 1517.7200 2292.7000 ;
        RECT 1516.1200 2297.6600 1517.7200 2298.1400 ;
        RECT 1516.1200 2303.1000 1517.7200 2303.5800 ;
        RECT 1523.8800 2281.3400 1525.4800 2281.8200 ;
        RECT 1523.8800 2286.7800 1525.4800 2287.2600 ;
        RECT 1516.1200 2281.3400 1517.7200 2281.8200 ;
        RECT 1516.1200 2286.7800 1517.7200 2287.2600 ;
        RECT 1523.8800 2265.0200 1525.4800 2265.5000 ;
        RECT 1523.8800 2270.4600 1525.4800 2270.9400 ;
        RECT 1523.8800 2275.9000 1525.4800 2276.3800 ;
        RECT 1516.1200 2265.0200 1517.7200 2265.5000 ;
        RECT 1516.1200 2270.4600 1517.7200 2270.9400 ;
        RECT 1516.1200 2275.9000 1517.7200 2276.3800 ;
        RECT 1516.1200 2259.5800 1517.7200 2260.0600 ;
        RECT 1523.8800 2259.5800 1525.4800 2260.0600 ;
        RECT 1510.5600 2461.8900 1720.7800 2463.4900 ;
        RECT 1510.5600 2255.3900 1720.7800 2256.9900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 2249.9600 1517.7200 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 2468.0000 1517.7200 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 2249.9600 1715.2200 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 2468.0000 1715.2200 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2255.3900 1512.1600 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2255.3900 1720.7800 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2461.8900 1512.1600 2463.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2461.8900 1720.7800 2463.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 2025.7500 1705.4800 2233.8500 ;
        RECT 1658.8800 2025.7500 1660.4800 2233.8500 ;
        RECT 1613.8800 2025.7500 1615.4800 2233.8500 ;
        RECT 1568.8800 2025.7500 1570.4800 2233.8500 ;
        RECT 1523.8800 2025.7500 1525.4800 2233.8500 ;
        RECT 1713.6200 2020.3200 1715.2200 2239.9600 ;
        RECT 1516.1200 2020.3200 1517.7200 2239.9600 ;
      LAYER met3 ;
        RECT 1713.6200 2214.9000 1715.2200 2215.3800 ;
        RECT 1713.6200 2220.3400 1715.2200 2220.8200 ;
        RECT 1703.8800 2214.9000 1705.4800 2215.3800 ;
        RECT 1703.8800 2220.3400 1705.4800 2220.8200 ;
        RECT 1703.8800 2225.7800 1705.4800 2226.2600 ;
        RECT 1713.6200 2225.7800 1715.2200 2226.2600 ;
        RECT 1713.6200 2204.0200 1715.2200 2204.5000 ;
        RECT 1713.6200 2209.4600 1715.2200 2209.9400 ;
        RECT 1703.8800 2204.0200 1705.4800 2204.5000 ;
        RECT 1703.8800 2209.4600 1705.4800 2209.9400 ;
        RECT 1713.6200 2187.7000 1715.2200 2188.1800 ;
        RECT 1713.6200 2193.1400 1715.2200 2193.6200 ;
        RECT 1703.8800 2187.7000 1705.4800 2188.1800 ;
        RECT 1703.8800 2193.1400 1705.4800 2193.6200 ;
        RECT 1703.8800 2198.5800 1705.4800 2199.0600 ;
        RECT 1713.6200 2198.5800 1715.2200 2199.0600 ;
        RECT 1658.8800 2214.9000 1660.4800 2215.3800 ;
        RECT 1658.8800 2220.3400 1660.4800 2220.8200 ;
        RECT 1658.8800 2225.7800 1660.4800 2226.2600 ;
        RECT 1658.8800 2204.0200 1660.4800 2204.5000 ;
        RECT 1658.8800 2209.4600 1660.4800 2209.9400 ;
        RECT 1658.8800 2187.7000 1660.4800 2188.1800 ;
        RECT 1658.8800 2193.1400 1660.4800 2193.6200 ;
        RECT 1658.8800 2198.5800 1660.4800 2199.0600 ;
        RECT 1713.6200 2171.3800 1715.2200 2171.8600 ;
        RECT 1713.6200 2176.8200 1715.2200 2177.3000 ;
        RECT 1713.6200 2182.2600 1715.2200 2182.7400 ;
        RECT 1703.8800 2171.3800 1705.4800 2171.8600 ;
        RECT 1703.8800 2176.8200 1705.4800 2177.3000 ;
        RECT 1703.8800 2182.2600 1705.4800 2182.7400 ;
        RECT 1713.6200 2160.5000 1715.2200 2160.9800 ;
        RECT 1713.6200 2165.9400 1715.2200 2166.4200 ;
        RECT 1703.8800 2160.5000 1705.4800 2160.9800 ;
        RECT 1703.8800 2165.9400 1705.4800 2166.4200 ;
        RECT 1713.6200 2144.1800 1715.2200 2144.6600 ;
        RECT 1713.6200 2149.6200 1715.2200 2150.1000 ;
        RECT 1713.6200 2155.0600 1715.2200 2155.5400 ;
        RECT 1703.8800 2144.1800 1705.4800 2144.6600 ;
        RECT 1703.8800 2149.6200 1705.4800 2150.1000 ;
        RECT 1703.8800 2155.0600 1705.4800 2155.5400 ;
        RECT 1713.6200 2133.3000 1715.2200 2133.7800 ;
        RECT 1713.6200 2138.7400 1715.2200 2139.2200 ;
        RECT 1703.8800 2133.3000 1705.4800 2133.7800 ;
        RECT 1703.8800 2138.7400 1705.4800 2139.2200 ;
        RECT 1658.8800 2171.3800 1660.4800 2171.8600 ;
        RECT 1658.8800 2176.8200 1660.4800 2177.3000 ;
        RECT 1658.8800 2182.2600 1660.4800 2182.7400 ;
        RECT 1658.8800 2160.5000 1660.4800 2160.9800 ;
        RECT 1658.8800 2165.9400 1660.4800 2166.4200 ;
        RECT 1658.8800 2144.1800 1660.4800 2144.6600 ;
        RECT 1658.8800 2149.6200 1660.4800 2150.1000 ;
        RECT 1658.8800 2155.0600 1660.4800 2155.5400 ;
        RECT 1658.8800 2133.3000 1660.4800 2133.7800 ;
        RECT 1658.8800 2138.7400 1660.4800 2139.2200 ;
        RECT 1613.8800 2214.9000 1615.4800 2215.3800 ;
        RECT 1613.8800 2220.3400 1615.4800 2220.8200 ;
        RECT 1613.8800 2225.7800 1615.4800 2226.2600 ;
        RECT 1568.8800 2214.9000 1570.4800 2215.3800 ;
        RECT 1568.8800 2220.3400 1570.4800 2220.8200 ;
        RECT 1568.8800 2225.7800 1570.4800 2226.2600 ;
        RECT 1613.8800 2204.0200 1615.4800 2204.5000 ;
        RECT 1613.8800 2209.4600 1615.4800 2209.9400 ;
        RECT 1613.8800 2187.7000 1615.4800 2188.1800 ;
        RECT 1613.8800 2193.1400 1615.4800 2193.6200 ;
        RECT 1613.8800 2198.5800 1615.4800 2199.0600 ;
        RECT 1568.8800 2204.0200 1570.4800 2204.5000 ;
        RECT 1568.8800 2209.4600 1570.4800 2209.9400 ;
        RECT 1568.8800 2187.7000 1570.4800 2188.1800 ;
        RECT 1568.8800 2193.1400 1570.4800 2193.6200 ;
        RECT 1568.8800 2198.5800 1570.4800 2199.0600 ;
        RECT 1523.8800 2214.9000 1525.4800 2215.3800 ;
        RECT 1523.8800 2220.3400 1525.4800 2220.8200 ;
        RECT 1516.1200 2214.9000 1517.7200 2215.3800 ;
        RECT 1516.1200 2220.3400 1517.7200 2220.8200 ;
        RECT 1516.1200 2225.7800 1517.7200 2226.2600 ;
        RECT 1523.8800 2225.7800 1525.4800 2226.2600 ;
        RECT 1523.8800 2204.0200 1525.4800 2204.5000 ;
        RECT 1523.8800 2209.4600 1525.4800 2209.9400 ;
        RECT 1516.1200 2204.0200 1517.7200 2204.5000 ;
        RECT 1516.1200 2209.4600 1517.7200 2209.9400 ;
        RECT 1523.8800 2187.7000 1525.4800 2188.1800 ;
        RECT 1523.8800 2193.1400 1525.4800 2193.6200 ;
        RECT 1516.1200 2187.7000 1517.7200 2188.1800 ;
        RECT 1516.1200 2193.1400 1517.7200 2193.6200 ;
        RECT 1516.1200 2198.5800 1517.7200 2199.0600 ;
        RECT 1523.8800 2198.5800 1525.4800 2199.0600 ;
        RECT 1613.8800 2171.3800 1615.4800 2171.8600 ;
        RECT 1613.8800 2176.8200 1615.4800 2177.3000 ;
        RECT 1613.8800 2182.2600 1615.4800 2182.7400 ;
        RECT 1613.8800 2160.5000 1615.4800 2160.9800 ;
        RECT 1613.8800 2165.9400 1615.4800 2166.4200 ;
        RECT 1568.8800 2171.3800 1570.4800 2171.8600 ;
        RECT 1568.8800 2176.8200 1570.4800 2177.3000 ;
        RECT 1568.8800 2182.2600 1570.4800 2182.7400 ;
        RECT 1568.8800 2160.5000 1570.4800 2160.9800 ;
        RECT 1568.8800 2165.9400 1570.4800 2166.4200 ;
        RECT 1613.8800 2144.1800 1615.4800 2144.6600 ;
        RECT 1613.8800 2149.6200 1615.4800 2150.1000 ;
        RECT 1613.8800 2155.0600 1615.4800 2155.5400 ;
        RECT 1613.8800 2133.3000 1615.4800 2133.7800 ;
        RECT 1613.8800 2138.7400 1615.4800 2139.2200 ;
        RECT 1568.8800 2144.1800 1570.4800 2144.6600 ;
        RECT 1568.8800 2149.6200 1570.4800 2150.1000 ;
        RECT 1568.8800 2155.0600 1570.4800 2155.5400 ;
        RECT 1568.8800 2133.3000 1570.4800 2133.7800 ;
        RECT 1568.8800 2138.7400 1570.4800 2139.2200 ;
        RECT 1523.8800 2171.3800 1525.4800 2171.8600 ;
        RECT 1523.8800 2176.8200 1525.4800 2177.3000 ;
        RECT 1523.8800 2182.2600 1525.4800 2182.7400 ;
        RECT 1516.1200 2171.3800 1517.7200 2171.8600 ;
        RECT 1516.1200 2176.8200 1517.7200 2177.3000 ;
        RECT 1516.1200 2182.2600 1517.7200 2182.7400 ;
        RECT 1523.8800 2160.5000 1525.4800 2160.9800 ;
        RECT 1523.8800 2165.9400 1525.4800 2166.4200 ;
        RECT 1516.1200 2160.5000 1517.7200 2160.9800 ;
        RECT 1516.1200 2165.9400 1517.7200 2166.4200 ;
        RECT 1523.8800 2144.1800 1525.4800 2144.6600 ;
        RECT 1523.8800 2149.6200 1525.4800 2150.1000 ;
        RECT 1523.8800 2155.0600 1525.4800 2155.5400 ;
        RECT 1516.1200 2144.1800 1517.7200 2144.6600 ;
        RECT 1516.1200 2149.6200 1517.7200 2150.1000 ;
        RECT 1516.1200 2155.0600 1517.7200 2155.5400 ;
        RECT 1523.8800 2133.3000 1525.4800 2133.7800 ;
        RECT 1523.8800 2138.7400 1525.4800 2139.2200 ;
        RECT 1516.1200 2133.3000 1517.7200 2133.7800 ;
        RECT 1516.1200 2138.7400 1517.7200 2139.2200 ;
        RECT 1713.6200 2116.9800 1715.2200 2117.4600 ;
        RECT 1713.6200 2122.4200 1715.2200 2122.9000 ;
        RECT 1713.6200 2127.8600 1715.2200 2128.3400 ;
        RECT 1703.8800 2116.9800 1705.4800 2117.4600 ;
        RECT 1703.8800 2122.4200 1705.4800 2122.9000 ;
        RECT 1703.8800 2127.8600 1705.4800 2128.3400 ;
        RECT 1713.6200 2106.1000 1715.2200 2106.5800 ;
        RECT 1713.6200 2111.5400 1715.2200 2112.0200 ;
        RECT 1703.8800 2106.1000 1705.4800 2106.5800 ;
        RECT 1703.8800 2111.5400 1705.4800 2112.0200 ;
        RECT 1713.6200 2089.7800 1715.2200 2090.2600 ;
        RECT 1713.6200 2095.2200 1715.2200 2095.7000 ;
        RECT 1713.6200 2100.6600 1715.2200 2101.1400 ;
        RECT 1703.8800 2089.7800 1705.4800 2090.2600 ;
        RECT 1703.8800 2095.2200 1705.4800 2095.7000 ;
        RECT 1703.8800 2100.6600 1705.4800 2101.1400 ;
        RECT 1713.6200 2078.9000 1715.2200 2079.3800 ;
        RECT 1713.6200 2084.3400 1715.2200 2084.8200 ;
        RECT 1703.8800 2078.9000 1705.4800 2079.3800 ;
        RECT 1703.8800 2084.3400 1705.4800 2084.8200 ;
        RECT 1658.8800 2116.9800 1660.4800 2117.4600 ;
        RECT 1658.8800 2122.4200 1660.4800 2122.9000 ;
        RECT 1658.8800 2127.8600 1660.4800 2128.3400 ;
        RECT 1658.8800 2106.1000 1660.4800 2106.5800 ;
        RECT 1658.8800 2111.5400 1660.4800 2112.0200 ;
        RECT 1658.8800 2089.7800 1660.4800 2090.2600 ;
        RECT 1658.8800 2095.2200 1660.4800 2095.7000 ;
        RECT 1658.8800 2100.6600 1660.4800 2101.1400 ;
        RECT 1658.8800 2078.9000 1660.4800 2079.3800 ;
        RECT 1658.8800 2084.3400 1660.4800 2084.8200 ;
        RECT 1713.6200 2062.5800 1715.2200 2063.0600 ;
        RECT 1713.6200 2068.0200 1715.2200 2068.5000 ;
        RECT 1713.6200 2073.4600 1715.2200 2073.9400 ;
        RECT 1703.8800 2062.5800 1705.4800 2063.0600 ;
        RECT 1703.8800 2068.0200 1705.4800 2068.5000 ;
        RECT 1703.8800 2073.4600 1705.4800 2073.9400 ;
        RECT 1713.6200 2051.7000 1715.2200 2052.1800 ;
        RECT 1713.6200 2057.1400 1715.2200 2057.6200 ;
        RECT 1703.8800 2051.7000 1705.4800 2052.1800 ;
        RECT 1703.8800 2057.1400 1705.4800 2057.6200 ;
        RECT 1713.6200 2035.3800 1715.2200 2035.8600 ;
        RECT 1713.6200 2040.8200 1715.2200 2041.3000 ;
        RECT 1713.6200 2046.2600 1715.2200 2046.7400 ;
        RECT 1703.8800 2035.3800 1705.4800 2035.8600 ;
        RECT 1703.8800 2040.8200 1705.4800 2041.3000 ;
        RECT 1703.8800 2046.2600 1705.4800 2046.7400 ;
        RECT 1703.8800 2029.9400 1705.4800 2030.4200 ;
        RECT 1713.6200 2029.9400 1715.2200 2030.4200 ;
        RECT 1658.8800 2062.5800 1660.4800 2063.0600 ;
        RECT 1658.8800 2068.0200 1660.4800 2068.5000 ;
        RECT 1658.8800 2073.4600 1660.4800 2073.9400 ;
        RECT 1658.8800 2051.7000 1660.4800 2052.1800 ;
        RECT 1658.8800 2057.1400 1660.4800 2057.6200 ;
        RECT 1658.8800 2035.3800 1660.4800 2035.8600 ;
        RECT 1658.8800 2040.8200 1660.4800 2041.3000 ;
        RECT 1658.8800 2046.2600 1660.4800 2046.7400 ;
        RECT 1658.8800 2029.9400 1660.4800 2030.4200 ;
        RECT 1613.8800 2116.9800 1615.4800 2117.4600 ;
        RECT 1613.8800 2122.4200 1615.4800 2122.9000 ;
        RECT 1613.8800 2127.8600 1615.4800 2128.3400 ;
        RECT 1613.8800 2106.1000 1615.4800 2106.5800 ;
        RECT 1613.8800 2111.5400 1615.4800 2112.0200 ;
        RECT 1568.8800 2116.9800 1570.4800 2117.4600 ;
        RECT 1568.8800 2122.4200 1570.4800 2122.9000 ;
        RECT 1568.8800 2127.8600 1570.4800 2128.3400 ;
        RECT 1568.8800 2106.1000 1570.4800 2106.5800 ;
        RECT 1568.8800 2111.5400 1570.4800 2112.0200 ;
        RECT 1613.8800 2089.7800 1615.4800 2090.2600 ;
        RECT 1613.8800 2095.2200 1615.4800 2095.7000 ;
        RECT 1613.8800 2100.6600 1615.4800 2101.1400 ;
        RECT 1613.8800 2078.9000 1615.4800 2079.3800 ;
        RECT 1613.8800 2084.3400 1615.4800 2084.8200 ;
        RECT 1568.8800 2089.7800 1570.4800 2090.2600 ;
        RECT 1568.8800 2095.2200 1570.4800 2095.7000 ;
        RECT 1568.8800 2100.6600 1570.4800 2101.1400 ;
        RECT 1568.8800 2078.9000 1570.4800 2079.3800 ;
        RECT 1568.8800 2084.3400 1570.4800 2084.8200 ;
        RECT 1523.8800 2116.9800 1525.4800 2117.4600 ;
        RECT 1523.8800 2122.4200 1525.4800 2122.9000 ;
        RECT 1523.8800 2127.8600 1525.4800 2128.3400 ;
        RECT 1516.1200 2116.9800 1517.7200 2117.4600 ;
        RECT 1516.1200 2122.4200 1517.7200 2122.9000 ;
        RECT 1516.1200 2127.8600 1517.7200 2128.3400 ;
        RECT 1523.8800 2106.1000 1525.4800 2106.5800 ;
        RECT 1523.8800 2111.5400 1525.4800 2112.0200 ;
        RECT 1516.1200 2106.1000 1517.7200 2106.5800 ;
        RECT 1516.1200 2111.5400 1517.7200 2112.0200 ;
        RECT 1523.8800 2089.7800 1525.4800 2090.2600 ;
        RECT 1523.8800 2095.2200 1525.4800 2095.7000 ;
        RECT 1523.8800 2100.6600 1525.4800 2101.1400 ;
        RECT 1516.1200 2089.7800 1517.7200 2090.2600 ;
        RECT 1516.1200 2095.2200 1517.7200 2095.7000 ;
        RECT 1516.1200 2100.6600 1517.7200 2101.1400 ;
        RECT 1523.8800 2078.9000 1525.4800 2079.3800 ;
        RECT 1523.8800 2084.3400 1525.4800 2084.8200 ;
        RECT 1516.1200 2078.9000 1517.7200 2079.3800 ;
        RECT 1516.1200 2084.3400 1517.7200 2084.8200 ;
        RECT 1613.8800 2062.5800 1615.4800 2063.0600 ;
        RECT 1613.8800 2068.0200 1615.4800 2068.5000 ;
        RECT 1613.8800 2073.4600 1615.4800 2073.9400 ;
        RECT 1613.8800 2051.7000 1615.4800 2052.1800 ;
        RECT 1613.8800 2057.1400 1615.4800 2057.6200 ;
        RECT 1568.8800 2062.5800 1570.4800 2063.0600 ;
        RECT 1568.8800 2068.0200 1570.4800 2068.5000 ;
        RECT 1568.8800 2073.4600 1570.4800 2073.9400 ;
        RECT 1568.8800 2051.7000 1570.4800 2052.1800 ;
        RECT 1568.8800 2057.1400 1570.4800 2057.6200 ;
        RECT 1613.8800 2035.3800 1615.4800 2035.8600 ;
        RECT 1613.8800 2040.8200 1615.4800 2041.3000 ;
        RECT 1613.8800 2046.2600 1615.4800 2046.7400 ;
        RECT 1613.8800 2029.9400 1615.4800 2030.4200 ;
        RECT 1568.8800 2035.3800 1570.4800 2035.8600 ;
        RECT 1568.8800 2040.8200 1570.4800 2041.3000 ;
        RECT 1568.8800 2046.2600 1570.4800 2046.7400 ;
        RECT 1568.8800 2029.9400 1570.4800 2030.4200 ;
        RECT 1523.8800 2062.5800 1525.4800 2063.0600 ;
        RECT 1523.8800 2068.0200 1525.4800 2068.5000 ;
        RECT 1523.8800 2073.4600 1525.4800 2073.9400 ;
        RECT 1516.1200 2062.5800 1517.7200 2063.0600 ;
        RECT 1516.1200 2068.0200 1517.7200 2068.5000 ;
        RECT 1516.1200 2073.4600 1517.7200 2073.9400 ;
        RECT 1523.8800 2051.7000 1525.4800 2052.1800 ;
        RECT 1523.8800 2057.1400 1525.4800 2057.6200 ;
        RECT 1516.1200 2051.7000 1517.7200 2052.1800 ;
        RECT 1516.1200 2057.1400 1517.7200 2057.6200 ;
        RECT 1523.8800 2035.3800 1525.4800 2035.8600 ;
        RECT 1523.8800 2040.8200 1525.4800 2041.3000 ;
        RECT 1523.8800 2046.2600 1525.4800 2046.7400 ;
        RECT 1516.1200 2035.3800 1517.7200 2035.8600 ;
        RECT 1516.1200 2040.8200 1517.7200 2041.3000 ;
        RECT 1516.1200 2046.2600 1517.7200 2046.7400 ;
        RECT 1516.1200 2029.9400 1517.7200 2030.4200 ;
        RECT 1523.8800 2029.9400 1525.4800 2030.4200 ;
        RECT 1510.5600 2232.2500 1720.7800 2233.8500 ;
        RECT 1510.5600 2025.7500 1720.7800 2027.3500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 2020.3200 1517.7200 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 2238.3600 1517.7200 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 2020.3200 1715.2200 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 2238.3600 1715.2200 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2025.7500 1512.1600 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2025.7500 1720.7800 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2232.2500 1512.1600 2233.8500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2232.2500 1720.7800 2233.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 1796.1100 1705.4800 2004.2100 ;
        RECT 1658.8800 1796.1100 1660.4800 2004.2100 ;
        RECT 1613.8800 1796.1100 1615.4800 2004.2100 ;
        RECT 1568.8800 1796.1100 1570.4800 2004.2100 ;
        RECT 1523.8800 1796.1100 1525.4800 2004.2100 ;
        RECT 1713.6200 1790.6800 1715.2200 2010.3200 ;
        RECT 1516.1200 1790.6800 1517.7200 2010.3200 ;
      LAYER met3 ;
        RECT 1713.6200 1985.2600 1715.2200 1985.7400 ;
        RECT 1713.6200 1990.7000 1715.2200 1991.1800 ;
        RECT 1703.8800 1985.2600 1705.4800 1985.7400 ;
        RECT 1703.8800 1990.7000 1705.4800 1991.1800 ;
        RECT 1703.8800 1996.1400 1705.4800 1996.6200 ;
        RECT 1713.6200 1996.1400 1715.2200 1996.6200 ;
        RECT 1713.6200 1974.3800 1715.2200 1974.8600 ;
        RECT 1713.6200 1979.8200 1715.2200 1980.3000 ;
        RECT 1703.8800 1974.3800 1705.4800 1974.8600 ;
        RECT 1703.8800 1979.8200 1705.4800 1980.3000 ;
        RECT 1713.6200 1958.0600 1715.2200 1958.5400 ;
        RECT 1713.6200 1963.5000 1715.2200 1963.9800 ;
        RECT 1703.8800 1958.0600 1705.4800 1958.5400 ;
        RECT 1703.8800 1963.5000 1705.4800 1963.9800 ;
        RECT 1703.8800 1968.9400 1705.4800 1969.4200 ;
        RECT 1713.6200 1968.9400 1715.2200 1969.4200 ;
        RECT 1658.8800 1985.2600 1660.4800 1985.7400 ;
        RECT 1658.8800 1990.7000 1660.4800 1991.1800 ;
        RECT 1658.8800 1996.1400 1660.4800 1996.6200 ;
        RECT 1658.8800 1974.3800 1660.4800 1974.8600 ;
        RECT 1658.8800 1979.8200 1660.4800 1980.3000 ;
        RECT 1658.8800 1958.0600 1660.4800 1958.5400 ;
        RECT 1658.8800 1963.5000 1660.4800 1963.9800 ;
        RECT 1658.8800 1968.9400 1660.4800 1969.4200 ;
        RECT 1713.6200 1941.7400 1715.2200 1942.2200 ;
        RECT 1713.6200 1947.1800 1715.2200 1947.6600 ;
        RECT 1713.6200 1952.6200 1715.2200 1953.1000 ;
        RECT 1703.8800 1941.7400 1705.4800 1942.2200 ;
        RECT 1703.8800 1947.1800 1705.4800 1947.6600 ;
        RECT 1703.8800 1952.6200 1705.4800 1953.1000 ;
        RECT 1713.6200 1930.8600 1715.2200 1931.3400 ;
        RECT 1713.6200 1936.3000 1715.2200 1936.7800 ;
        RECT 1703.8800 1930.8600 1705.4800 1931.3400 ;
        RECT 1703.8800 1936.3000 1705.4800 1936.7800 ;
        RECT 1713.6200 1914.5400 1715.2200 1915.0200 ;
        RECT 1713.6200 1919.9800 1715.2200 1920.4600 ;
        RECT 1713.6200 1925.4200 1715.2200 1925.9000 ;
        RECT 1703.8800 1914.5400 1705.4800 1915.0200 ;
        RECT 1703.8800 1919.9800 1705.4800 1920.4600 ;
        RECT 1703.8800 1925.4200 1705.4800 1925.9000 ;
        RECT 1713.6200 1903.6600 1715.2200 1904.1400 ;
        RECT 1713.6200 1909.1000 1715.2200 1909.5800 ;
        RECT 1703.8800 1903.6600 1705.4800 1904.1400 ;
        RECT 1703.8800 1909.1000 1705.4800 1909.5800 ;
        RECT 1658.8800 1941.7400 1660.4800 1942.2200 ;
        RECT 1658.8800 1947.1800 1660.4800 1947.6600 ;
        RECT 1658.8800 1952.6200 1660.4800 1953.1000 ;
        RECT 1658.8800 1930.8600 1660.4800 1931.3400 ;
        RECT 1658.8800 1936.3000 1660.4800 1936.7800 ;
        RECT 1658.8800 1914.5400 1660.4800 1915.0200 ;
        RECT 1658.8800 1919.9800 1660.4800 1920.4600 ;
        RECT 1658.8800 1925.4200 1660.4800 1925.9000 ;
        RECT 1658.8800 1903.6600 1660.4800 1904.1400 ;
        RECT 1658.8800 1909.1000 1660.4800 1909.5800 ;
        RECT 1613.8800 1985.2600 1615.4800 1985.7400 ;
        RECT 1613.8800 1990.7000 1615.4800 1991.1800 ;
        RECT 1613.8800 1996.1400 1615.4800 1996.6200 ;
        RECT 1568.8800 1985.2600 1570.4800 1985.7400 ;
        RECT 1568.8800 1990.7000 1570.4800 1991.1800 ;
        RECT 1568.8800 1996.1400 1570.4800 1996.6200 ;
        RECT 1613.8800 1974.3800 1615.4800 1974.8600 ;
        RECT 1613.8800 1979.8200 1615.4800 1980.3000 ;
        RECT 1613.8800 1958.0600 1615.4800 1958.5400 ;
        RECT 1613.8800 1963.5000 1615.4800 1963.9800 ;
        RECT 1613.8800 1968.9400 1615.4800 1969.4200 ;
        RECT 1568.8800 1974.3800 1570.4800 1974.8600 ;
        RECT 1568.8800 1979.8200 1570.4800 1980.3000 ;
        RECT 1568.8800 1958.0600 1570.4800 1958.5400 ;
        RECT 1568.8800 1963.5000 1570.4800 1963.9800 ;
        RECT 1568.8800 1968.9400 1570.4800 1969.4200 ;
        RECT 1523.8800 1985.2600 1525.4800 1985.7400 ;
        RECT 1523.8800 1990.7000 1525.4800 1991.1800 ;
        RECT 1516.1200 1985.2600 1517.7200 1985.7400 ;
        RECT 1516.1200 1990.7000 1517.7200 1991.1800 ;
        RECT 1516.1200 1996.1400 1517.7200 1996.6200 ;
        RECT 1523.8800 1996.1400 1525.4800 1996.6200 ;
        RECT 1523.8800 1974.3800 1525.4800 1974.8600 ;
        RECT 1523.8800 1979.8200 1525.4800 1980.3000 ;
        RECT 1516.1200 1974.3800 1517.7200 1974.8600 ;
        RECT 1516.1200 1979.8200 1517.7200 1980.3000 ;
        RECT 1523.8800 1958.0600 1525.4800 1958.5400 ;
        RECT 1523.8800 1963.5000 1525.4800 1963.9800 ;
        RECT 1516.1200 1958.0600 1517.7200 1958.5400 ;
        RECT 1516.1200 1963.5000 1517.7200 1963.9800 ;
        RECT 1516.1200 1968.9400 1517.7200 1969.4200 ;
        RECT 1523.8800 1968.9400 1525.4800 1969.4200 ;
        RECT 1613.8800 1941.7400 1615.4800 1942.2200 ;
        RECT 1613.8800 1947.1800 1615.4800 1947.6600 ;
        RECT 1613.8800 1952.6200 1615.4800 1953.1000 ;
        RECT 1613.8800 1930.8600 1615.4800 1931.3400 ;
        RECT 1613.8800 1936.3000 1615.4800 1936.7800 ;
        RECT 1568.8800 1941.7400 1570.4800 1942.2200 ;
        RECT 1568.8800 1947.1800 1570.4800 1947.6600 ;
        RECT 1568.8800 1952.6200 1570.4800 1953.1000 ;
        RECT 1568.8800 1930.8600 1570.4800 1931.3400 ;
        RECT 1568.8800 1936.3000 1570.4800 1936.7800 ;
        RECT 1613.8800 1914.5400 1615.4800 1915.0200 ;
        RECT 1613.8800 1919.9800 1615.4800 1920.4600 ;
        RECT 1613.8800 1925.4200 1615.4800 1925.9000 ;
        RECT 1613.8800 1903.6600 1615.4800 1904.1400 ;
        RECT 1613.8800 1909.1000 1615.4800 1909.5800 ;
        RECT 1568.8800 1914.5400 1570.4800 1915.0200 ;
        RECT 1568.8800 1919.9800 1570.4800 1920.4600 ;
        RECT 1568.8800 1925.4200 1570.4800 1925.9000 ;
        RECT 1568.8800 1903.6600 1570.4800 1904.1400 ;
        RECT 1568.8800 1909.1000 1570.4800 1909.5800 ;
        RECT 1523.8800 1941.7400 1525.4800 1942.2200 ;
        RECT 1523.8800 1947.1800 1525.4800 1947.6600 ;
        RECT 1523.8800 1952.6200 1525.4800 1953.1000 ;
        RECT 1516.1200 1941.7400 1517.7200 1942.2200 ;
        RECT 1516.1200 1947.1800 1517.7200 1947.6600 ;
        RECT 1516.1200 1952.6200 1517.7200 1953.1000 ;
        RECT 1523.8800 1930.8600 1525.4800 1931.3400 ;
        RECT 1523.8800 1936.3000 1525.4800 1936.7800 ;
        RECT 1516.1200 1930.8600 1517.7200 1931.3400 ;
        RECT 1516.1200 1936.3000 1517.7200 1936.7800 ;
        RECT 1523.8800 1914.5400 1525.4800 1915.0200 ;
        RECT 1523.8800 1919.9800 1525.4800 1920.4600 ;
        RECT 1523.8800 1925.4200 1525.4800 1925.9000 ;
        RECT 1516.1200 1914.5400 1517.7200 1915.0200 ;
        RECT 1516.1200 1919.9800 1517.7200 1920.4600 ;
        RECT 1516.1200 1925.4200 1517.7200 1925.9000 ;
        RECT 1523.8800 1903.6600 1525.4800 1904.1400 ;
        RECT 1523.8800 1909.1000 1525.4800 1909.5800 ;
        RECT 1516.1200 1903.6600 1517.7200 1904.1400 ;
        RECT 1516.1200 1909.1000 1517.7200 1909.5800 ;
        RECT 1713.6200 1887.3400 1715.2200 1887.8200 ;
        RECT 1713.6200 1892.7800 1715.2200 1893.2600 ;
        RECT 1713.6200 1898.2200 1715.2200 1898.7000 ;
        RECT 1703.8800 1887.3400 1705.4800 1887.8200 ;
        RECT 1703.8800 1892.7800 1705.4800 1893.2600 ;
        RECT 1703.8800 1898.2200 1705.4800 1898.7000 ;
        RECT 1713.6200 1876.4600 1715.2200 1876.9400 ;
        RECT 1713.6200 1881.9000 1715.2200 1882.3800 ;
        RECT 1703.8800 1876.4600 1705.4800 1876.9400 ;
        RECT 1703.8800 1881.9000 1705.4800 1882.3800 ;
        RECT 1713.6200 1860.1400 1715.2200 1860.6200 ;
        RECT 1713.6200 1865.5800 1715.2200 1866.0600 ;
        RECT 1713.6200 1871.0200 1715.2200 1871.5000 ;
        RECT 1703.8800 1860.1400 1705.4800 1860.6200 ;
        RECT 1703.8800 1865.5800 1705.4800 1866.0600 ;
        RECT 1703.8800 1871.0200 1705.4800 1871.5000 ;
        RECT 1713.6200 1849.2600 1715.2200 1849.7400 ;
        RECT 1713.6200 1854.7000 1715.2200 1855.1800 ;
        RECT 1703.8800 1849.2600 1705.4800 1849.7400 ;
        RECT 1703.8800 1854.7000 1705.4800 1855.1800 ;
        RECT 1658.8800 1887.3400 1660.4800 1887.8200 ;
        RECT 1658.8800 1892.7800 1660.4800 1893.2600 ;
        RECT 1658.8800 1898.2200 1660.4800 1898.7000 ;
        RECT 1658.8800 1876.4600 1660.4800 1876.9400 ;
        RECT 1658.8800 1881.9000 1660.4800 1882.3800 ;
        RECT 1658.8800 1860.1400 1660.4800 1860.6200 ;
        RECT 1658.8800 1865.5800 1660.4800 1866.0600 ;
        RECT 1658.8800 1871.0200 1660.4800 1871.5000 ;
        RECT 1658.8800 1849.2600 1660.4800 1849.7400 ;
        RECT 1658.8800 1854.7000 1660.4800 1855.1800 ;
        RECT 1713.6200 1832.9400 1715.2200 1833.4200 ;
        RECT 1713.6200 1838.3800 1715.2200 1838.8600 ;
        RECT 1713.6200 1843.8200 1715.2200 1844.3000 ;
        RECT 1703.8800 1832.9400 1705.4800 1833.4200 ;
        RECT 1703.8800 1838.3800 1705.4800 1838.8600 ;
        RECT 1703.8800 1843.8200 1705.4800 1844.3000 ;
        RECT 1713.6200 1822.0600 1715.2200 1822.5400 ;
        RECT 1713.6200 1827.5000 1715.2200 1827.9800 ;
        RECT 1703.8800 1822.0600 1705.4800 1822.5400 ;
        RECT 1703.8800 1827.5000 1705.4800 1827.9800 ;
        RECT 1713.6200 1805.7400 1715.2200 1806.2200 ;
        RECT 1713.6200 1811.1800 1715.2200 1811.6600 ;
        RECT 1713.6200 1816.6200 1715.2200 1817.1000 ;
        RECT 1703.8800 1805.7400 1705.4800 1806.2200 ;
        RECT 1703.8800 1811.1800 1705.4800 1811.6600 ;
        RECT 1703.8800 1816.6200 1705.4800 1817.1000 ;
        RECT 1703.8800 1800.3000 1705.4800 1800.7800 ;
        RECT 1713.6200 1800.3000 1715.2200 1800.7800 ;
        RECT 1658.8800 1832.9400 1660.4800 1833.4200 ;
        RECT 1658.8800 1838.3800 1660.4800 1838.8600 ;
        RECT 1658.8800 1843.8200 1660.4800 1844.3000 ;
        RECT 1658.8800 1822.0600 1660.4800 1822.5400 ;
        RECT 1658.8800 1827.5000 1660.4800 1827.9800 ;
        RECT 1658.8800 1805.7400 1660.4800 1806.2200 ;
        RECT 1658.8800 1811.1800 1660.4800 1811.6600 ;
        RECT 1658.8800 1816.6200 1660.4800 1817.1000 ;
        RECT 1658.8800 1800.3000 1660.4800 1800.7800 ;
        RECT 1613.8800 1887.3400 1615.4800 1887.8200 ;
        RECT 1613.8800 1892.7800 1615.4800 1893.2600 ;
        RECT 1613.8800 1898.2200 1615.4800 1898.7000 ;
        RECT 1613.8800 1876.4600 1615.4800 1876.9400 ;
        RECT 1613.8800 1881.9000 1615.4800 1882.3800 ;
        RECT 1568.8800 1887.3400 1570.4800 1887.8200 ;
        RECT 1568.8800 1892.7800 1570.4800 1893.2600 ;
        RECT 1568.8800 1898.2200 1570.4800 1898.7000 ;
        RECT 1568.8800 1876.4600 1570.4800 1876.9400 ;
        RECT 1568.8800 1881.9000 1570.4800 1882.3800 ;
        RECT 1613.8800 1860.1400 1615.4800 1860.6200 ;
        RECT 1613.8800 1865.5800 1615.4800 1866.0600 ;
        RECT 1613.8800 1871.0200 1615.4800 1871.5000 ;
        RECT 1613.8800 1849.2600 1615.4800 1849.7400 ;
        RECT 1613.8800 1854.7000 1615.4800 1855.1800 ;
        RECT 1568.8800 1860.1400 1570.4800 1860.6200 ;
        RECT 1568.8800 1865.5800 1570.4800 1866.0600 ;
        RECT 1568.8800 1871.0200 1570.4800 1871.5000 ;
        RECT 1568.8800 1849.2600 1570.4800 1849.7400 ;
        RECT 1568.8800 1854.7000 1570.4800 1855.1800 ;
        RECT 1523.8800 1887.3400 1525.4800 1887.8200 ;
        RECT 1523.8800 1892.7800 1525.4800 1893.2600 ;
        RECT 1523.8800 1898.2200 1525.4800 1898.7000 ;
        RECT 1516.1200 1887.3400 1517.7200 1887.8200 ;
        RECT 1516.1200 1892.7800 1517.7200 1893.2600 ;
        RECT 1516.1200 1898.2200 1517.7200 1898.7000 ;
        RECT 1523.8800 1876.4600 1525.4800 1876.9400 ;
        RECT 1523.8800 1881.9000 1525.4800 1882.3800 ;
        RECT 1516.1200 1876.4600 1517.7200 1876.9400 ;
        RECT 1516.1200 1881.9000 1517.7200 1882.3800 ;
        RECT 1523.8800 1860.1400 1525.4800 1860.6200 ;
        RECT 1523.8800 1865.5800 1525.4800 1866.0600 ;
        RECT 1523.8800 1871.0200 1525.4800 1871.5000 ;
        RECT 1516.1200 1860.1400 1517.7200 1860.6200 ;
        RECT 1516.1200 1865.5800 1517.7200 1866.0600 ;
        RECT 1516.1200 1871.0200 1517.7200 1871.5000 ;
        RECT 1523.8800 1849.2600 1525.4800 1849.7400 ;
        RECT 1523.8800 1854.7000 1525.4800 1855.1800 ;
        RECT 1516.1200 1849.2600 1517.7200 1849.7400 ;
        RECT 1516.1200 1854.7000 1517.7200 1855.1800 ;
        RECT 1613.8800 1832.9400 1615.4800 1833.4200 ;
        RECT 1613.8800 1838.3800 1615.4800 1838.8600 ;
        RECT 1613.8800 1843.8200 1615.4800 1844.3000 ;
        RECT 1613.8800 1822.0600 1615.4800 1822.5400 ;
        RECT 1613.8800 1827.5000 1615.4800 1827.9800 ;
        RECT 1568.8800 1832.9400 1570.4800 1833.4200 ;
        RECT 1568.8800 1838.3800 1570.4800 1838.8600 ;
        RECT 1568.8800 1843.8200 1570.4800 1844.3000 ;
        RECT 1568.8800 1822.0600 1570.4800 1822.5400 ;
        RECT 1568.8800 1827.5000 1570.4800 1827.9800 ;
        RECT 1613.8800 1805.7400 1615.4800 1806.2200 ;
        RECT 1613.8800 1811.1800 1615.4800 1811.6600 ;
        RECT 1613.8800 1816.6200 1615.4800 1817.1000 ;
        RECT 1613.8800 1800.3000 1615.4800 1800.7800 ;
        RECT 1568.8800 1805.7400 1570.4800 1806.2200 ;
        RECT 1568.8800 1811.1800 1570.4800 1811.6600 ;
        RECT 1568.8800 1816.6200 1570.4800 1817.1000 ;
        RECT 1568.8800 1800.3000 1570.4800 1800.7800 ;
        RECT 1523.8800 1832.9400 1525.4800 1833.4200 ;
        RECT 1523.8800 1838.3800 1525.4800 1838.8600 ;
        RECT 1523.8800 1843.8200 1525.4800 1844.3000 ;
        RECT 1516.1200 1832.9400 1517.7200 1833.4200 ;
        RECT 1516.1200 1838.3800 1517.7200 1838.8600 ;
        RECT 1516.1200 1843.8200 1517.7200 1844.3000 ;
        RECT 1523.8800 1822.0600 1525.4800 1822.5400 ;
        RECT 1523.8800 1827.5000 1525.4800 1827.9800 ;
        RECT 1516.1200 1822.0600 1517.7200 1822.5400 ;
        RECT 1516.1200 1827.5000 1517.7200 1827.9800 ;
        RECT 1523.8800 1805.7400 1525.4800 1806.2200 ;
        RECT 1523.8800 1811.1800 1525.4800 1811.6600 ;
        RECT 1523.8800 1816.6200 1525.4800 1817.1000 ;
        RECT 1516.1200 1805.7400 1517.7200 1806.2200 ;
        RECT 1516.1200 1811.1800 1517.7200 1811.6600 ;
        RECT 1516.1200 1816.6200 1517.7200 1817.1000 ;
        RECT 1516.1200 1800.3000 1517.7200 1800.7800 ;
        RECT 1523.8800 1800.3000 1525.4800 1800.7800 ;
        RECT 1510.5600 2002.6100 1720.7800 2004.2100 ;
        RECT 1510.5600 1796.1100 1720.7800 1797.7100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1790.6800 1517.7200 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 2008.7200 1517.7200 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1790.6800 1715.2200 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 2008.7200 1715.2200 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1796.1100 1512.1600 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1796.1100 1720.7800 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 2002.6100 1512.1600 2004.2100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 2002.6100 1720.7800 2004.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 1566.4700 1705.4800 1774.5700 ;
        RECT 1658.8800 1566.4700 1660.4800 1774.5700 ;
        RECT 1613.8800 1566.4700 1615.4800 1774.5700 ;
        RECT 1568.8800 1566.4700 1570.4800 1774.5700 ;
        RECT 1523.8800 1566.4700 1525.4800 1774.5700 ;
        RECT 1713.6200 1561.0400 1715.2200 1780.6800 ;
        RECT 1516.1200 1561.0400 1517.7200 1780.6800 ;
      LAYER met3 ;
        RECT 1713.6200 1755.6200 1715.2200 1756.1000 ;
        RECT 1713.6200 1761.0600 1715.2200 1761.5400 ;
        RECT 1703.8800 1755.6200 1705.4800 1756.1000 ;
        RECT 1703.8800 1761.0600 1705.4800 1761.5400 ;
        RECT 1703.8800 1766.5000 1705.4800 1766.9800 ;
        RECT 1713.6200 1766.5000 1715.2200 1766.9800 ;
        RECT 1713.6200 1744.7400 1715.2200 1745.2200 ;
        RECT 1713.6200 1750.1800 1715.2200 1750.6600 ;
        RECT 1703.8800 1744.7400 1705.4800 1745.2200 ;
        RECT 1703.8800 1750.1800 1705.4800 1750.6600 ;
        RECT 1713.6200 1728.4200 1715.2200 1728.9000 ;
        RECT 1713.6200 1733.8600 1715.2200 1734.3400 ;
        RECT 1703.8800 1728.4200 1705.4800 1728.9000 ;
        RECT 1703.8800 1733.8600 1705.4800 1734.3400 ;
        RECT 1703.8800 1739.3000 1705.4800 1739.7800 ;
        RECT 1713.6200 1739.3000 1715.2200 1739.7800 ;
        RECT 1658.8800 1755.6200 1660.4800 1756.1000 ;
        RECT 1658.8800 1761.0600 1660.4800 1761.5400 ;
        RECT 1658.8800 1766.5000 1660.4800 1766.9800 ;
        RECT 1658.8800 1744.7400 1660.4800 1745.2200 ;
        RECT 1658.8800 1750.1800 1660.4800 1750.6600 ;
        RECT 1658.8800 1728.4200 1660.4800 1728.9000 ;
        RECT 1658.8800 1733.8600 1660.4800 1734.3400 ;
        RECT 1658.8800 1739.3000 1660.4800 1739.7800 ;
        RECT 1713.6200 1712.1000 1715.2200 1712.5800 ;
        RECT 1713.6200 1717.5400 1715.2200 1718.0200 ;
        RECT 1713.6200 1722.9800 1715.2200 1723.4600 ;
        RECT 1703.8800 1712.1000 1705.4800 1712.5800 ;
        RECT 1703.8800 1717.5400 1705.4800 1718.0200 ;
        RECT 1703.8800 1722.9800 1705.4800 1723.4600 ;
        RECT 1713.6200 1701.2200 1715.2200 1701.7000 ;
        RECT 1713.6200 1706.6600 1715.2200 1707.1400 ;
        RECT 1703.8800 1701.2200 1705.4800 1701.7000 ;
        RECT 1703.8800 1706.6600 1705.4800 1707.1400 ;
        RECT 1713.6200 1684.9000 1715.2200 1685.3800 ;
        RECT 1713.6200 1690.3400 1715.2200 1690.8200 ;
        RECT 1713.6200 1695.7800 1715.2200 1696.2600 ;
        RECT 1703.8800 1684.9000 1705.4800 1685.3800 ;
        RECT 1703.8800 1690.3400 1705.4800 1690.8200 ;
        RECT 1703.8800 1695.7800 1705.4800 1696.2600 ;
        RECT 1713.6200 1674.0200 1715.2200 1674.5000 ;
        RECT 1713.6200 1679.4600 1715.2200 1679.9400 ;
        RECT 1703.8800 1674.0200 1705.4800 1674.5000 ;
        RECT 1703.8800 1679.4600 1705.4800 1679.9400 ;
        RECT 1658.8800 1712.1000 1660.4800 1712.5800 ;
        RECT 1658.8800 1717.5400 1660.4800 1718.0200 ;
        RECT 1658.8800 1722.9800 1660.4800 1723.4600 ;
        RECT 1658.8800 1701.2200 1660.4800 1701.7000 ;
        RECT 1658.8800 1706.6600 1660.4800 1707.1400 ;
        RECT 1658.8800 1684.9000 1660.4800 1685.3800 ;
        RECT 1658.8800 1690.3400 1660.4800 1690.8200 ;
        RECT 1658.8800 1695.7800 1660.4800 1696.2600 ;
        RECT 1658.8800 1674.0200 1660.4800 1674.5000 ;
        RECT 1658.8800 1679.4600 1660.4800 1679.9400 ;
        RECT 1613.8800 1755.6200 1615.4800 1756.1000 ;
        RECT 1613.8800 1761.0600 1615.4800 1761.5400 ;
        RECT 1613.8800 1766.5000 1615.4800 1766.9800 ;
        RECT 1568.8800 1755.6200 1570.4800 1756.1000 ;
        RECT 1568.8800 1761.0600 1570.4800 1761.5400 ;
        RECT 1568.8800 1766.5000 1570.4800 1766.9800 ;
        RECT 1613.8800 1744.7400 1615.4800 1745.2200 ;
        RECT 1613.8800 1750.1800 1615.4800 1750.6600 ;
        RECT 1613.8800 1728.4200 1615.4800 1728.9000 ;
        RECT 1613.8800 1733.8600 1615.4800 1734.3400 ;
        RECT 1613.8800 1739.3000 1615.4800 1739.7800 ;
        RECT 1568.8800 1744.7400 1570.4800 1745.2200 ;
        RECT 1568.8800 1750.1800 1570.4800 1750.6600 ;
        RECT 1568.8800 1728.4200 1570.4800 1728.9000 ;
        RECT 1568.8800 1733.8600 1570.4800 1734.3400 ;
        RECT 1568.8800 1739.3000 1570.4800 1739.7800 ;
        RECT 1523.8800 1755.6200 1525.4800 1756.1000 ;
        RECT 1523.8800 1761.0600 1525.4800 1761.5400 ;
        RECT 1516.1200 1755.6200 1517.7200 1756.1000 ;
        RECT 1516.1200 1761.0600 1517.7200 1761.5400 ;
        RECT 1516.1200 1766.5000 1517.7200 1766.9800 ;
        RECT 1523.8800 1766.5000 1525.4800 1766.9800 ;
        RECT 1523.8800 1744.7400 1525.4800 1745.2200 ;
        RECT 1523.8800 1750.1800 1525.4800 1750.6600 ;
        RECT 1516.1200 1744.7400 1517.7200 1745.2200 ;
        RECT 1516.1200 1750.1800 1517.7200 1750.6600 ;
        RECT 1523.8800 1728.4200 1525.4800 1728.9000 ;
        RECT 1523.8800 1733.8600 1525.4800 1734.3400 ;
        RECT 1516.1200 1728.4200 1517.7200 1728.9000 ;
        RECT 1516.1200 1733.8600 1517.7200 1734.3400 ;
        RECT 1516.1200 1739.3000 1517.7200 1739.7800 ;
        RECT 1523.8800 1739.3000 1525.4800 1739.7800 ;
        RECT 1613.8800 1712.1000 1615.4800 1712.5800 ;
        RECT 1613.8800 1717.5400 1615.4800 1718.0200 ;
        RECT 1613.8800 1722.9800 1615.4800 1723.4600 ;
        RECT 1613.8800 1701.2200 1615.4800 1701.7000 ;
        RECT 1613.8800 1706.6600 1615.4800 1707.1400 ;
        RECT 1568.8800 1712.1000 1570.4800 1712.5800 ;
        RECT 1568.8800 1717.5400 1570.4800 1718.0200 ;
        RECT 1568.8800 1722.9800 1570.4800 1723.4600 ;
        RECT 1568.8800 1701.2200 1570.4800 1701.7000 ;
        RECT 1568.8800 1706.6600 1570.4800 1707.1400 ;
        RECT 1613.8800 1684.9000 1615.4800 1685.3800 ;
        RECT 1613.8800 1690.3400 1615.4800 1690.8200 ;
        RECT 1613.8800 1695.7800 1615.4800 1696.2600 ;
        RECT 1613.8800 1674.0200 1615.4800 1674.5000 ;
        RECT 1613.8800 1679.4600 1615.4800 1679.9400 ;
        RECT 1568.8800 1684.9000 1570.4800 1685.3800 ;
        RECT 1568.8800 1690.3400 1570.4800 1690.8200 ;
        RECT 1568.8800 1695.7800 1570.4800 1696.2600 ;
        RECT 1568.8800 1674.0200 1570.4800 1674.5000 ;
        RECT 1568.8800 1679.4600 1570.4800 1679.9400 ;
        RECT 1523.8800 1712.1000 1525.4800 1712.5800 ;
        RECT 1523.8800 1717.5400 1525.4800 1718.0200 ;
        RECT 1523.8800 1722.9800 1525.4800 1723.4600 ;
        RECT 1516.1200 1712.1000 1517.7200 1712.5800 ;
        RECT 1516.1200 1717.5400 1517.7200 1718.0200 ;
        RECT 1516.1200 1722.9800 1517.7200 1723.4600 ;
        RECT 1523.8800 1701.2200 1525.4800 1701.7000 ;
        RECT 1523.8800 1706.6600 1525.4800 1707.1400 ;
        RECT 1516.1200 1701.2200 1517.7200 1701.7000 ;
        RECT 1516.1200 1706.6600 1517.7200 1707.1400 ;
        RECT 1523.8800 1684.9000 1525.4800 1685.3800 ;
        RECT 1523.8800 1690.3400 1525.4800 1690.8200 ;
        RECT 1523.8800 1695.7800 1525.4800 1696.2600 ;
        RECT 1516.1200 1684.9000 1517.7200 1685.3800 ;
        RECT 1516.1200 1690.3400 1517.7200 1690.8200 ;
        RECT 1516.1200 1695.7800 1517.7200 1696.2600 ;
        RECT 1523.8800 1674.0200 1525.4800 1674.5000 ;
        RECT 1523.8800 1679.4600 1525.4800 1679.9400 ;
        RECT 1516.1200 1674.0200 1517.7200 1674.5000 ;
        RECT 1516.1200 1679.4600 1517.7200 1679.9400 ;
        RECT 1713.6200 1657.7000 1715.2200 1658.1800 ;
        RECT 1713.6200 1663.1400 1715.2200 1663.6200 ;
        RECT 1713.6200 1668.5800 1715.2200 1669.0600 ;
        RECT 1703.8800 1657.7000 1705.4800 1658.1800 ;
        RECT 1703.8800 1663.1400 1705.4800 1663.6200 ;
        RECT 1703.8800 1668.5800 1705.4800 1669.0600 ;
        RECT 1713.6200 1646.8200 1715.2200 1647.3000 ;
        RECT 1713.6200 1652.2600 1715.2200 1652.7400 ;
        RECT 1703.8800 1646.8200 1705.4800 1647.3000 ;
        RECT 1703.8800 1652.2600 1705.4800 1652.7400 ;
        RECT 1713.6200 1630.5000 1715.2200 1630.9800 ;
        RECT 1713.6200 1635.9400 1715.2200 1636.4200 ;
        RECT 1713.6200 1641.3800 1715.2200 1641.8600 ;
        RECT 1703.8800 1630.5000 1705.4800 1630.9800 ;
        RECT 1703.8800 1635.9400 1705.4800 1636.4200 ;
        RECT 1703.8800 1641.3800 1705.4800 1641.8600 ;
        RECT 1713.6200 1619.6200 1715.2200 1620.1000 ;
        RECT 1713.6200 1625.0600 1715.2200 1625.5400 ;
        RECT 1703.8800 1619.6200 1705.4800 1620.1000 ;
        RECT 1703.8800 1625.0600 1705.4800 1625.5400 ;
        RECT 1658.8800 1657.7000 1660.4800 1658.1800 ;
        RECT 1658.8800 1663.1400 1660.4800 1663.6200 ;
        RECT 1658.8800 1668.5800 1660.4800 1669.0600 ;
        RECT 1658.8800 1646.8200 1660.4800 1647.3000 ;
        RECT 1658.8800 1652.2600 1660.4800 1652.7400 ;
        RECT 1658.8800 1630.5000 1660.4800 1630.9800 ;
        RECT 1658.8800 1635.9400 1660.4800 1636.4200 ;
        RECT 1658.8800 1641.3800 1660.4800 1641.8600 ;
        RECT 1658.8800 1619.6200 1660.4800 1620.1000 ;
        RECT 1658.8800 1625.0600 1660.4800 1625.5400 ;
        RECT 1713.6200 1603.3000 1715.2200 1603.7800 ;
        RECT 1713.6200 1608.7400 1715.2200 1609.2200 ;
        RECT 1713.6200 1614.1800 1715.2200 1614.6600 ;
        RECT 1703.8800 1603.3000 1705.4800 1603.7800 ;
        RECT 1703.8800 1608.7400 1705.4800 1609.2200 ;
        RECT 1703.8800 1614.1800 1705.4800 1614.6600 ;
        RECT 1713.6200 1592.4200 1715.2200 1592.9000 ;
        RECT 1713.6200 1597.8600 1715.2200 1598.3400 ;
        RECT 1703.8800 1592.4200 1705.4800 1592.9000 ;
        RECT 1703.8800 1597.8600 1705.4800 1598.3400 ;
        RECT 1713.6200 1576.1000 1715.2200 1576.5800 ;
        RECT 1713.6200 1581.5400 1715.2200 1582.0200 ;
        RECT 1713.6200 1586.9800 1715.2200 1587.4600 ;
        RECT 1703.8800 1576.1000 1705.4800 1576.5800 ;
        RECT 1703.8800 1581.5400 1705.4800 1582.0200 ;
        RECT 1703.8800 1586.9800 1705.4800 1587.4600 ;
        RECT 1703.8800 1570.6600 1705.4800 1571.1400 ;
        RECT 1713.6200 1570.6600 1715.2200 1571.1400 ;
        RECT 1658.8800 1603.3000 1660.4800 1603.7800 ;
        RECT 1658.8800 1608.7400 1660.4800 1609.2200 ;
        RECT 1658.8800 1614.1800 1660.4800 1614.6600 ;
        RECT 1658.8800 1592.4200 1660.4800 1592.9000 ;
        RECT 1658.8800 1597.8600 1660.4800 1598.3400 ;
        RECT 1658.8800 1576.1000 1660.4800 1576.5800 ;
        RECT 1658.8800 1581.5400 1660.4800 1582.0200 ;
        RECT 1658.8800 1586.9800 1660.4800 1587.4600 ;
        RECT 1658.8800 1570.6600 1660.4800 1571.1400 ;
        RECT 1613.8800 1657.7000 1615.4800 1658.1800 ;
        RECT 1613.8800 1663.1400 1615.4800 1663.6200 ;
        RECT 1613.8800 1668.5800 1615.4800 1669.0600 ;
        RECT 1613.8800 1646.8200 1615.4800 1647.3000 ;
        RECT 1613.8800 1652.2600 1615.4800 1652.7400 ;
        RECT 1568.8800 1657.7000 1570.4800 1658.1800 ;
        RECT 1568.8800 1663.1400 1570.4800 1663.6200 ;
        RECT 1568.8800 1668.5800 1570.4800 1669.0600 ;
        RECT 1568.8800 1646.8200 1570.4800 1647.3000 ;
        RECT 1568.8800 1652.2600 1570.4800 1652.7400 ;
        RECT 1613.8800 1630.5000 1615.4800 1630.9800 ;
        RECT 1613.8800 1635.9400 1615.4800 1636.4200 ;
        RECT 1613.8800 1641.3800 1615.4800 1641.8600 ;
        RECT 1613.8800 1619.6200 1615.4800 1620.1000 ;
        RECT 1613.8800 1625.0600 1615.4800 1625.5400 ;
        RECT 1568.8800 1630.5000 1570.4800 1630.9800 ;
        RECT 1568.8800 1635.9400 1570.4800 1636.4200 ;
        RECT 1568.8800 1641.3800 1570.4800 1641.8600 ;
        RECT 1568.8800 1619.6200 1570.4800 1620.1000 ;
        RECT 1568.8800 1625.0600 1570.4800 1625.5400 ;
        RECT 1523.8800 1657.7000 1525.4800 1658.1800 ;
        RECT 1523.8800 1663.1400 1525.4800 1663.6200 ;
        RECT 1523.8800 1668.5800 1525.4800 1669.0600 ;
        RECT 1516.1200 1657.7000 1517.7200 1658.1800 ;
        RECT 1516.1200 1663.1400 1517.7200 1663.6200 ;
        RECT 1516.1200 1668.5800 1517.7200 1669.0600 ;
        RECT 1523.8800 1646.8200 1525.4800 1647.3000 ;
        RECT 1523.8800 1652.2600 1525.4800 1652.7400 ;
        RECT 1516.1200 1646.8200 1517.7200 1647.3000 ;
        RECT 1516.1200 1652.2600 1517.7200 1652.7400 ;
        RECT 1523.8800 1630.5000 1525.4800 1630.9800 ;
        RECT 1523.8800 1635.9400 1525.4800 1636.4200 ;
        RECT 1523.8800 1641.3800 1525.4800 1641.8600 ;
        RECT 1516.1200 1630.5000 1517.7200 1630.9800 ;
        RECT 1516.1200 1635.9400 1517.7200 1636.4200 ;
        RECT 1516.1200 1641.3800 1517.7200 1641.8600 ;
        RECT 1523.8800 1619.6200 1525.4800 1620.1000 ;
        RECT 1523.8800 1625.0600 1525.4800 1625.5400 ;
        RECT 1516.1200 1619.6200 1517.7200 1620.1000 ;
        RECT 1516.1200 1625.0600 1517.7200 1625.5400 ;
        RECT 1613.8800 1603.3000 1615.4800 1603.7800 ;
        RECT 1613.8800 1608.7400 1615.4800 1609.2200 ;
        RECT 1613.8800 1614.1800 1615.4800 1614.6600 ;
        RECT 1613.8800 1592.4200 1615.4800 1592.9000 ;
        RECT 1613.8800 1597.8600 1615.4800 1598.3400 ;
        RECT 1568.8800 1603.3000 1570.4800 1603.7800 ;
        RECT 1568.8800 1608.7400 1570.4800 1609.2200 ;
        RECT 1568.8800 1614.1800 1570.4800 1614.6600 ;
        RECT 1568.8800 1592.4200 1570.4800 1592.9000 ;
        RECT 1568.8800 1597.8600 1570.4800 1598.3400 ;
        RECT 1613.8800 1576.1000 1615.4800 1576.5800 ;
        RECT 1613.8800 1581.5400 1615.4800 1582.0200 ;
        RECT 1613.8800 1586.9800 1615.4800 1587.4600 ;
        RECT 1613.8800 1570.6600 1615.4800 1571.1400 ;
        RECT 1568.8800 1576.1000 1570.4800 1576.5800 ;
        RECT 1568.8800 1581.5400 1570.4800 1582.0200 ;
        RECT 1568.8800 1586.9800 1570.4800 1587.4600 ;
        RECT 1568.8800 1570.6600 1570.4800 1571.1400 ;
        RECT 1523.8800 1603.3000 1525.4800 1603.7800 ;
        RECT 1523.8800 1608.7400 1525.4800 1609.2200 ;
        RECT 1523.8800 1614.1800 1525.4800 1614.6600 ;
        RECT 1516.1200 1603.3000 1517.7200 1603.7800 ;
        RECT 1516.1200 1608.7400 1517.7200 1609.2200 ;
        RECT 1516.1200 1614.1800 1517.7200 1614.6600 ;
        RECT 1523.8800 1592.4200 1525.4800 1592.9000 ;
        RECT 1523.8800 1597.8600 1525.4800 1598.3400 ;
        RECT 1516.1200 1592.4200 1517.7200 1592.9000 ;
        RECT 1516.1200 1597.8600 1517.7200 1598.3400 ;
        RECT 1523.8800 1576.1000 1525.4800 1576.5800 ;
        RECT 1523.8800 1581.5400 1525.4800 1582.0200 ;
        RECT 1523.8800 1586.9800 1525.4800 1587.4600 ;
        RECT 1516.1200 1576.1000 1517.7200 1576.5800 ;
        RECT 1516.1200 1581.5400 1517.7200 1582.0200 ;
        RECT 1516.1200 1586.9800 1517.7200 1587.4600 ;
        RECT 1516.1200 1570.6600 1517.7200 1571.1400 ;
        RECT 1523.8800 1570.6600 1525.4800 1571.1400 ;
        RECT 1510.5600 1772.9700 1720.7800 1774.5700 ;
        RECT 1510.5600 1566.4700 1720.7800 1568.0700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1561.0400 1517.7200 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1779.0800 1517.7200 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1561.0400 1715.2200 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1779.0800 1715.2200 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1566.4700 1512.1600 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1566.4700 1720.7800 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1772.9700 1512.1600 1774.5700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1772.9700 1720.7800 1774.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 1336.8300 1705.4800 1544.9300 ;
        RECT 1658.8800 1336.8300 1660.4800 1544.9300 ;
        RECT 1613.8800 1336.8300 1615.4800 1544.9300 ;
        RECT 1568.8800 1336.8300 1570.4800 1544.9300 ;
        RECT 1523.8800 1336.8300 1525.4800 1544.9300 ;
        RECT 1713.6200 1331.4000 1715.2200 1551.0400 ;
        RECT 1516.1200 1331.4000 1517.7200 1551.0400 ;
      LAYER met3 ;
        RECT 1713.6200 1525.9800 1715.2200 1526.4600 ;
        RECT 1713.6200 1531.4200 1715.2200 1531.9000 ;
        RECT 1703.8800 1525.9800 1705.4800 1526.4600 ;
        RECT 1703.8800 1531.4200 1705.4800 1531.9000 ;
        RECT 1703.8800 1536.8600 1705.4800 1537.3400 ;
        RECT 1713.6200 1536.8600 1715.2200 1537.3400 ;
        RECT 1713.6200 1515.1000 1715.2200 1515.5800 ;
        RECT 1713.6200 1520.5400 1715.2200 1521.0200 ;
        RECT 1703.8800 1515.1000 1705.4800 1515.5800 ;
        RECT 1703.8800 1520.5400 1705.4800 1521.0200 ;
        RECT 1713.6200 1498.7800 1715.2200 1499.2600 ;
        RECT 1713.6200 1504.2200 1715.2200 1504.7000 ;
        RECT 1703.8800 1498.7800 1705.4800 1499.2600 ;
        RECT 1703.8800 1504.2200 1705.4800 1504.7000 ;
        RECT 1703.8800 1509.6600 1705.4800 1510.1400 ;
        RECT 1713.6200 1509.6600 1715.2200 1510.1400 ;
        RECT 1658.8800 1525.9800 1660.4800 1526.4600 ;
        RECT 1658.8800 1531.4200 1660.4800 1531.9000 ;
        RECT 1658.8800 1536.8600 1660.4800 1537.3400 ;
        RECT 1658.8800 1515.1000 1660.4800 1515.5800 ;
        RECT 1658.8800 1520.5400 1660.4800 1521.0200 ;
        RECT 1658.8800 1498.7800 1660.4800 1499.2600 ;
        RECT 1658.8800 1504.2200 1660.4800 1504.7000 ;
        RECT 1658.8800 1509.6600 1660.4800 1510.1400 ;
        RECT 1713.6200 1482.4600 1715.2200 1482.9400 ;
        RECT 1713.6200 1487.9000 1715.2200 1488.3800 ;
        RECT 1713.6200 1493.3400 1715.2200 1493.8200 ;
        RECT 1703.8800 1482.4600 1705.4800 1482.9400 ;
        RECT 1703.8800 1487.9000 1705.4800 1488.3800 ;
        RECT 1703.8800 1493.3400 1705.4800 1493.8200 ;
        RECT 1713.6200 1471.5800 1715.2200 1472.0600 ;
        RECT 1713.6200 1477.0200 1715.2200 1477.5000 ;
        RECT 1703.8800 1471.5800 1705.4800 1472.0600 ;
        RECT 1703.8800 1477.0200 1705.4800 1477.5000 ;
        RECT 1713.6200 1455.2600 1715.2200 1455.7400 ;
        RECT 1713.6200 1460.7000 1715.2200 1461.1800 ;
        RECT 1713.6200 1466.1400 1715.2200 1466.6200 ;
        RECT 1703.8800 1455.2600 1705.4800 1455.7400 ;
        RECT 1703.8800 1460.7000 1705.4800 1461.1800 ;
        RECT 1703.8800 1466.1400 1705.4800 1466.6200 ;
        RECT 1713.6200 1444.3800 1715.2200 1444.8600 ;
        RECT 1713.6200 1449.8200 1715.2200 1450.3000 ;
        RECT 1703.8800 1444.3800 1705.4800 1444.8600 ;
        RECT 1703.8800 1449.8200 1705.4800 1450.3000 ;
        RECT 1658.8800 1482.4600 1660.4800 1482.9400 ;
        RECT 1658.8800 1487.9000 1660.4800 1488.3800 ;
        RECT 1658.8800 1493.3400 1660.4800 1493.8200 ;
        RECT 1658.8800 1471.5800 1660.4800 1472.0600 ;
        RECT 1658.8800 1477.0200 1660.4800 1477.5000 ;
        RECT 1658.8800 1455.2600 1660.4800 1455.7400 ;
        RECT 1658.8800 1460.7000 1660.4800 1461.1800 ;
        RECT 1658.8800 1466.1400 1660.4800 1466.6200 ;
        RECT 1658.8800 1444.3800 1660.4800 1444.8600 ;
        RECT 1658.8800 1449.8200 1660.4800 1450.3000 ;
        RECT 1613.8800 1525.9800 1615.4800 1526.4600 ;
        RECT 1613.8800 1531.4200 1615.4800 1531.9000 ;
        RECT 1613.8800 1536.8600 1615.4800 1537.3400 ;
        RECT 1568.8800 1525.9800 1570.4800 1526.4600 ;
        RECT 1568.8800 1531.4200 1570.4800 1531.9000 ;
        RECT 1568.8800 1536.8600 1570.4800 1537.3400 ;
        RECT 1613.8800 1515.1000 1615.4800 1515.5800 ;
        RECT 1613.8800 1520.5400 1615.4800 1521.0200 ;
        RECT 1613.8800 1498.7800 1615.4800 1499.2600 ;
        RECT 1613.8800 1504.2200 1615.4800 1504.7000 ;
        RECT 1613.8800 1509.6600 1615.4800 1510.1400 ;
        RECT 1568.8800 1515.1000 1570.4800 1515.5800 ;
        RECT 1568.8800 1520.5400 1570.4800 1521.0200 ;
        RECT 1568.8800 1498.7800 1570.4800 1499.2600 ;
        RECT 1568.8800 1504.2200 1570.4800 1504.7000 ;
        RECT 1568.8800 1509.6600 1570.4800 1510.1400 ;
        RECT 1523.8800 1525.9800 1525.4800 1526.4600 ;
        RECT 1523.8800 1531.4200 1525.4800 1531.9000 ;
        RECT 1516.1200 1525.9800 1517.7200 1526.4600 ;
        RECT 1516.1200 1531.4200 1517.7200 1531.9000 ;
        RECT 1516.1200 1536.8600 1517.7200 1537.3400 ;
        RECT 1523.8800 1536.8600 1525.4800 1537.3400 ;
        RECT 1523.8800 1515.1000 1525.4800 1515.5800 ;
        RECT 1523.8800 1520.5400 1525.4800 1521.0200 ;
        RECT 1516.1200 1515.1000 1517.7200 1515.5800 ;
        RECT 1516.1200 1520.5400 1517.7200 1521.0200 ;
        RECT 1523.8800 1498.7800 1525.4800 1499.2600 ;
        RECT 1523.8800 1504.2200 1525.4800 1504.7000 ;
        RECT 1516.1200 1498.7800 1517.7200 1499.2600 ;
        RECT 1516.1200 1504.2200 1517.7200 1504.7000 ;
        RECT 1516.1200 1509.6600 1517.7200 1510.1400 ;
        RECT 1523.8800 1509.6600 1525.4800 1510.1400 ;
        RECT 1613.8800 1482.4600 1615.4800 1482.9400 ;
        RECT 1613.8800 1487.9000 1615.4800 1488.3800 ;
        RECT 1613.8800 1493.3400 1615.4800 1493.8200 ;
        RECT 1613.8800 1471.5800 1615.4800 1472.0600 ;
        RECT 1613.8800 1477.0200 1615.4800 1477.5000 ;
        RECT 1568.8800 1482.4600 1570.4800 1482.9400 ;
        RECT 1568.8800 1487.9000 1570.4800 1488.3800 ;
        RECT 1568.8800 1493.3400 1570.4800 1493.8200 ;
        RECT 1568.8800 1471.5800 1570.4800 1472.0600 ;
        RECT 1568.8800 1477.0200 1570.4800 1477.5000 ;
        RECT 1613.8800 1455.2600 1615.4800 1455.7400 ;
        RECT 1613.8800 1460.7000 1615.4800 1461.1800 ;
        RECT 1613.8800 1466.1400 1615.4800 1466.6200 ;
        RECT 1613.8800 1444.3800 1615.4800 1444.8600 ;
        RECT 1613.8800 1449.8200 1615.4800 1450.3000 ;
        RECT 1568.8800 1455.2600 1570.4800 1455.7400 ;
        RECT 1568.8800 1460.7000 1570.4800 1461.1800 ;
        RECT 1568.8800 1466.1400 1570.4800 1466.6200 ;
        RECT 1568.8800 1444.3800 1570.4800 1444.8600 ;
        RECT 1568.8800 1449.8200 1570.4800 1450.3000 ;
        RECT 1523.8800 1482.4600 1525.4800 1482.9400 ;
        RECT 1523.8800 1487.9000 1525.4800 1488.3800 ;
        RECT 1523.8800 1493.3400 1525.4800 1493.8200 ;
        RECT 1516.1200 1482.4600 1517.7200 1482.9400 ;
        RECT 1516.1200 1487.9000 1517.7200 1488.3800 ;
        RECT 1516.1200 1493.3400 1517.7200 1493.8200 ;
        RECT 1523.8800 1471.5800 1525.4800 1472.0600 ;
        RECT 1523.8800 1477.0200 1525.4800 1477.5000 ;
        RECT 1516.1200 1471.5800 1517.7200 1472.0600 ;
        RECT 1516.1200 1477.0200 1517.7200 1477.5000 ;
        RECT 1523.8800 1455.2600 1525.4800 1455.7400 ;
        RECT 1523.8800 1460.7000 1525.4800 1461.1800 ;
        RECT 1523.8800 1466.1400 1525.4800 1466.6200 ;
        RECT 1516.1200 1455.2600 1517.7200 1455.7400 ;
        RECT 1516.1200 1460.7000 1517.7200 1461.1800 ;
        RECT 1516.1200 1466.1400 1517.7200 1466.6200 ;
        RECT 1523.8800 1444.3800 1525.4800 1444.8600 ;
        RECT 1523.8800 1449.8200 1525.4800 1450.3000 ;
        RECT 1516.1200 1444.3800 1517.7200 1444.8600 ;
        RECT 1516.1200 1449.8200 1517.7200 1450.3000 ;
        RECT 1713.6200 1428.0600 1715.2200 1428.5400 ;
        RECT 1713.6200 1433.5000 1715.2200 1433.9800 ;
        RECT 1713.6200 1438.9400 1715.2200 1439.4200 ;
        RECT 1703.8800 1428.0600 1705.4800 1428.5400 ;
        RECT 1703.8800 1433.5000 1705.4800 1433.9800 ;
        RECT 1703.8800 1438.9400 1705.4800 1439.4200 ;
        RECT 1713.6200 1417.1800 1715.2200 1417.6600 ;
        RECT 1713.6200 1422.6200 1715.2200 1423.1000 ;
        RECT 1703.8800 1417.1800 1705.4800 1417.6600 ;
        RECT 1703.8800 1422.6200 1705.4800 1423.1000 ;
        RECT 1713.6200 1400.8600 1715.2200 1401.3400 ;
        RECT 1713.6200 1406.3000 1715.2200 1406.7800 ;
        RECT 1713.6200 1411.7400 1715.2200 1412.2200 ;
        RECT 1703.8800 1400.8600 1705.4800 1401.3400 ;
        RECT 1703.8800 1406.3000 1705.4800 1406.7800 ;
        RECT 1703.8800 1411.7400 1705.4800 1412.2200 ;
        RECT 1713.6200 1389.9800 1715.2200 1390.4600 ;
        RECT 1713.6200 1395.4200 1715.2200 1395.9000 ;
        RECT 1703.8800 1389.9800 1705.4800 1390.4600 ;
        RECT 1703.8800 1395.4200 1705.4800 1395.9000 ;
        RECT 1658.8800 1428.0600 1660.4800 1428.5400 ;
        RECT 1658.8800 1433.5000 1660.4800 1433.9800 ;
        RECT 1658.8800 1438.9400 1660.4800 1439.4200 ;
        RECT 1658.8800 1417.1800 1660.4800 1417.6600 ;
        RECT 1658.8800 1422.6200 1660.4800 1423.1000 ;
        RECT 1658.8800 1400.8600 1660.4800 1401.3400 ;
        RECT 1658.8800 1406.3000 1660.4800 1406.7800 ;
        RECT 1658.8800 1411.7400 1660.4800 1412.2200 ;
        RECT 1658.8800 1389.9800 1660.4800 1390.4600 ;
        RECT 1658.8800 1395.4200 1660.4800 1395.9000 ;
        RECT 1713.6200 1373.6600 1715.2200 1374.1400 ;
        RECT 1713.6200 1379.1000 1715.2200 1379.5800 ;
        RECT 1713.6200 1384.5400 1715.2200 1385.0200 ;
        RECT 1703.8800 1373.6600 1705.4800 1374.1400 ;
        RECT 1703.8800 1379.1000 1705.4800 1379.5800 ;
        RECT 1703.8800 1384.5400 1705.4800 1385.0200 ;
        RECT 1713.6200 1362.7800 1715.2200 1363.2600 ;
        RECT 1713.6200 1368.2200 1715.2200 1368.7000 ;
        RECT 1703.8800 1362.7800 1705.4800 1363.2600 ;
        RECT 1703.8800 1368.2200 1705.4800 1368.7000 ;
        RECT 1713.6200 1346.4600 1715.2200 1346.9400 ;
        RECT 1713.6200 1351.9000 1715.2200 1352.3800 ;
        RECT 1713.6200 1357.3400 1715.2200 1357.8200 ;
        RECT 1703.8800 1346.4600 1705.4800 1346.9400 ;
        RECT 1703.8800 1351.9000 1705.4800 1352.3800 ;
        RECT 1703.8800 1357.3400 1705.4800 1357.8200 ;
        RECT 1703.8800 1341.0200 1705.4800 1341.5000 ;
        RECT 1713.6200 1341.0200 1715.2200 1341.5000 ;
        RECT 1658.8800 1373.6600 1660.4800 1374.1400 ;
        RECT 1658.8800 1379.1000 1660.4800 1379.5800 ;
        RECT 1658.8800 1384.5400 1660.4800 1385.0200 ;
        RECT 1658.8800 1362.7800 1660.4800 1363.2600 ;
        RECT 1658.8800 1368.2200 1660.4800 1368.7000 ;
        RECT 1658.8800 1346.4600 1660.4800 1346.9400 ;
        RECT 1658.8800 1351.9000 1660.4800 1352.3800 ;
        RECT 1658.8800 1357.3400 1660.4800 1357.8200 ;
        RECT 1658.8800 1341.0200 1660.4800 1341.5000 ;
        RECT 1613.8800 1428.0600 1615.4800 1428.5400 ;
        RECT 1613.8800 1433.5000 1615.4800 1433.9800 ;
        RECT 1613.8800 1438.9400 1615.4800 1439.4200 ;
        RECT 1613.8800 1417.1800 1615.4800 1417.6600 ;
        RECT 1613.8800 1422.6200 1615.4800 1423.1000 ;
        RECT 1568.8800 1428.0600 1570.4800 1428.5400 ;
        RECT 1568.8800 1433.5000 1570.4800 1433.9800 ;
        RECT 1568.8800 1438.9400 1570.4800 1439.4200 ;
        RECT 1568.8800 1417.1800 1570.4800 1417.6600 ;
        RECT 1568.8800 1422.6200 1570.4800 1423.1000 ;
        RECT 1613.8800 1400.8600 1615.4800 1401.3400 ;
        RECT 1613.8800 1406.3000 1615.4800 1406.7800 ;
        RECT 1613.8800 1411.7400 1615.4800 1412.2200 ;
        RECT 1613.8800 1389.9800 1615.4800 1390.4600 ;
        RECT 1613.8800 1395.4200 1615.4800 1395.9000 ;
        RECT 1568.8800 1400.8600 1570.4800 1401.3400 ;
        RECT 1568.8800 1406.3000 1570.4800 1406.7800 ;
        RECT 1568.8800 1411.7400 1570.4800 1412.2200 ;
        RECT 1568.8800 1389.9800 1570.4800 1390.4600 ;
        RECT 1568.8800 1395.4200 1570.4800 1395.9000 ;
        RECT 1523.8800 1428.0600 1525.4800 1428.5400 ;
        RECT 1523.8800 1433.5000 1525.4800 1433.9800 ;
        RECT 1523.8800 1438.9400 1525.4800 1439.4200 ;
        RECT 1516.1200 1428.0600 1517.7200 1428.5400 ;
        RECT 1516.1200 1433.5000 1517.7200 1433.9800 ;
        RECT 1516.1200 1438.9400 1517.7200 1439.4200 ;
        RECT 1523.8800 1417.1800 1525.4800 1417.6600 ;
        RECT 1523.8800 1422.6200 1525.4800 1423.1000 ;
        RECT 1516.1200 1417.1800 1517.7200 1417.6600 ;
        RECT 1516.1200 1422.6200 1517.7200 1423.1000 ;
        RECT 1523.8800 1400.8600 1525.4800 1401.3400 ;
        RECT 1523.8800 1406.3000 1525.4800 1406.7800 ;
        RECT 1523.8800 1411.7400 1525.4800 1412.2200 ;
        RECT 1516.1200 1400.8600 1517.7200 1401.3400 ;
        RECT 1516.1200 1406.3000 1517.7200 1406.7800 ;
        RECT 1516.1200 1411.7400 1517.7200 1412.2200 ;
        RECT 1523.8800 1389.9800 1525.4800 1390.4600 ;
        RECT 1523.8800 1395.4200 1525.4800 1395.9000 ;
        RECT 1516.1200 1389.9800 1517.7200 1390.4600 ;
        RECT 1516.1200 1395.4200 1517.7200 1395.9000 ;
        RECT 1613.8800 1373.6600 1615.4800 1374.1400 ;
        RECT 1613.8800 1379.1000 1615.4800 1379.5800 ;
        RECT 1613.8800 1384.5400 1615.4800 1385.0200 ;
        RECT 1613.8800 1362.7800 1615.4800 1363.2600 ;
        RECT 1613.8800 1368.2200 1615.4800 1368.7000 ;
        RECT 1568.8800 1373.6600 1570.4800 1374.1400 ;
        RECT 1568.8800 1379.1000 1570.4800 1379.5800 ;
        RECT 1568.8800 1384.5400 1570.4800 1385.0200 ;
        RECT 1568.8800 1362.7800 1570.4800 1363.2600 ;
        RECT 1568.8800 1368.2200 1570.4800 1368.7000 ;
        RECT 1613.8800 1346.4600 1615.4800 1346.9400 ;
        RECT 1613.8800 1351.9000 1615.4800 1352.3800 ;
        RECT 1613.8800 1357.3400 1615.4800 1357.8200 ;
        RECT 1613.8800 1341.0200 1615.4800 1341.5000 ;
        RECT 1568.8800 1346.4600 1570.4800 1346.9400 ;
        RECT 1568.8800 1351.9000 1570.4800 1352.3800 ;
        RECT 1568.8800 1357.3400 1570.4800 1357.8200 ;
        RECT 1568.8800 1341.0200 1570.4800 1341.5000 ;
        RECT 1523.8800 1373.6600 1525.4800 1374.1400 ;
        RECT 1523.8800 1379.1000 1525.4800 1379.5800 ;
        RECT 1523.8800 1384.5400 1525.4800 1385.0200 ;
        RECT 1516.1200 1373.6600 1517.7200 1374.1400 ;
        RECT 1516.1200 1379.1000 1517.7200 1379.5800 ;
        RECT 1516.1200 1384.5400 1517.7200 1385.0200 ;
        RECT 1523.8800 1362.7800 1525.4800 1363.2600 ;
        RECT 1523.8800 1368.2200 1525.4800 1368.7000 ;
        RECT 1516.1200 1362.7800 1517.7200 1363.2600 ;
        RECT 1516.1200 1368.2200 1517.7200 1368.7000 ;
        RECT 1523.8800 1346.4600 1525.4800 1346.9400 ;
        RECT 1523.8800 1351.9000 1525.4800 1352.3800 ;
        RECT 1523.8800 1357.3400 1525.4800 1357.8200 ;
        RECT 1516.1200 1346.4600 1517.7200 1346.9400 ;
        RECT 1516.1200 1351.9000 1517.7200 1352.3800 ;
        RECT 1516.1200 1357.3400 1517.7200 1357.8200 ;
        RECT 1516.1200 1341.0200 1517.7200 1341.5000 ;
        RECT 1523.8800 1341.0200 1525.4800 1341.5000 ;
        RECT 1510.5600 1543.3300 1720.7800 1544.9300 ;
        RECT 1510.5600 1336.8300 1720.7800 1338.4300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1331.4000 1517.7200 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1549.4400 1517.7200 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1331.4000 1715.2200 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1549.4400 1715.2200 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1336.8300 1512.1600 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1336.8300 1720.7800 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1543.3300 1512.1600 1544.9300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1543.3300 1720.7800 1544.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 1107.1900 1705.4800 1315.2900 ;
        RECT 1658.8800 1107.1900 1660.4800 1315.2900 ;
        RECT 1613.8800 1107.1900 1615.4800 1315.2900 ;
        RECT 1568.8800 1107.1900 1570.4800 1315.2900 ;
        RECT 1523.8800 1107.1900 1525.4800 1315.2900 ;
        RECT 1713.6200 1101.7600 1715.2200 1321.4000 ;
        RECT 1516.1200 1101.7600 1517.7200 1321.4000 ;
      LAYER met3 ;
        RECT 1713.6200 1296.3400 1715.2200 1296.8200 ;
        RECT 1713.6200 1301.7800 1715.2200 1302.2600 ;
        RECT 1703.8800 1296.3400 1705.4800 1296.8200 ;
        RECT 1703.8800 1301.7800 1705.4800 1302.2600 ;
        RECT 1703.8800 1307.2200 1705.4800 1307.7000 ;
        RECT 1713.6200 1307.2200 1715.2200 1307.7000 ;
        RECT 1713.6200 1285.4600 1715.2200 1285.9400 ;
        RECT 1713.6200 1290.9000 1715.2200 1291.3800 ;
        RECT 1703.8800 1285.4600 1705.4800 1285.9400 ;
        RECT 1703.8800 1290.9000 1705.4800 1291.3800 ;
        RECT 1713.6200 1269.1400 1715.2200 1269.6200 ;
        RECT 1713.6200 1274.5800 1715.2200 1275.0600 ;
        RECT 1703.8800 1269.1400 1705.4800 1269.6200 ;
        RECT 1703.8800 1274.5800 1705.4800 1275.0600 ;
        RECT 1703.8800 1280.0200 1705.4800 1280.5000 ;
        RECT 1713.6200 1280.0200 1715.2200 1280.5000 ;
        RECT 1658.8800 1296.3400 1660.4800 1296.8200 ;
        RECT 1658.8800 1301.7800 1660.4800 1302.2600 ;
        RECT 1658.8800 1307.2200 1660.4800 1307.7000 ;
        RECT 1658.8800 1285.4600 1660.4800 1285.9400 ;
        RECT 1658.8800 1290.9000 1660.4800 1291.3800 ;
        RECT 1658.8800 1269.1400 1660.4800 1269.6200 ;
        RECT 1658.8800 1274.5800 1660.4800 1275.0600 ;
        RECT 1658.8800 1280.0200 1660.4800 1280.5000 ;
        RECT 1713.6200 1252.8200 1715.2200 1253.3000 ;
        RECT 1713.6200 1258.2600 1715.2200 1258.7400 ;
        RECT 1713.6200 1263.7000 1715.2200 1264.1800 ;
        RECT 1703.8800 1252.8200 1705.4800 1253.3000 ;
        RECT 1703.8800 1258.2600 1705.4800 1258.7400 ;
        RECT 1703.8800 1263.7000 1705.4800 1264.1800 ;
        RECT 1713.6200 1241.9400 1715.2200 1242.4200 ;
        RECT 1713.6200 1247.3800 1715.2200 1247.8600 ;
        RECT 1703.8800 1241.9400 1705.4800 1242.4200 ;
        RECT 1703.8800 1247.3800 1705.4800 1247.8600 ;
        RECT 1713.6200 1225.6200 1715.2200 1226.1000 ;
        RECT 1713.6200 1231.0600 1715.2200 1231.5400 ;
        RECT 1713.6200 1236.5000 1715.2200 1236.9800 ;
        RECT 1703.8800 1225.6200 1705.4800 1226.1000 ;
        RECT 1703.8800 1231.0600 1705.4800 1231.5400 ;
        RECT 1703.8800 1236.5000 1705.4800 1236.9800 ;
        RECT 1713.6200 1214.7400 1715.2200 1215.2200 ;
        RECT 1713.6200 1220.1800 1715.2200 1220.6600 ;
        RECT 1703.8800 1214.7400 1705.4800 1215.2200 ;
        RECT 1703.8800 1220.1800 1705.4800 1220.6600 ;
        RECT 1658.8800 1252.8200 1660.4800 1253.3000 ;
        RECT 1658.8800 1258.2600 1660.4800 1258.7400 ;
        RECT 1658.8800 1263.7000 1660.4800 1264.1800 ;
        RECT 1658.8800 1241.9400 1660.4800 1242.4200 ;
        RECT 1658.8800 1247.3800 1660.4800 1247.8600 ;
        RECT 1658.8800 1225.6200 1660.4800 1226.1000 ;
        RECT 1658.8800 1231.0600 1660.4800 1231.5400 ;
        RECT 1658.8800 1236.5000 1660.4800 1236.9800 ;
        RECT 1658.8800 1214.7400 1660.4800 1215.2200 ;
        RECT 1658.8800 1220.1800 1660.4800 1220.6600 ;
        RECT 1613.8800 1296.3400 1615.4800 1296.8200 ;
        RECT 1613.8800 1301.7800 1615.4800 1302.2600 ;
        RECT 1613.8800 1307.2200 1615.4800 1307.7000 ;
        RECT 1568.8800 1296.3400 1570.4800 1296.8200 ;
        RECT 1568.8800 1301.7800 1570.4800 1302.2600 ;
        RECT 1568.8800 1307.2200 1570.4800 1307.7000 ;
        RECT 1613.8800 1285.4600 1615.4800 1285.9400 ;
        RECT 1613.8800 1290.9000 1615.4800 1291.3800 ;
        RECT 1613.8800 1269.1400 1615.4800 1269.6200 ;
        RECT 1613.8800 1274.5800 1615.4800 1275.0600 ;
        RECT 1613.8800 1280.0200 1615.4800 1280.5000 ;
        RECT 1568.8800 1285.4600 1570.4800 1285.9400 ;
        RECT 1568.8800 1290.9000 1570.4800 1291.3800 ;
        RECT 1568.8800 1269.1400 1570.4800 1269.6200 ;
        RECT 1568.8800 1274.5800 1570.4800 1275.0600 ;
        RECT 1568.8800 1280.0200 1570.4800 1280.5000 ;
        RECT 1523.8800 1296.3400 1525.4800 1296.8200 ;
        RECT 1523.8800 1301.7800 1525.4800 1302.2600 ;
        RECT 1516.1200 1296.3400 1517.7200 1296.8200 ;
        RECT 1516.1200 1301.7800 1517.7200 1302.2600 ;
        RECT 1516.1200 1307.2200 1517.7200 1307.7000 ;
        RECT 1523.8800 1307.2200 1525.4800 1307.7000 ;
        RECT 1523.8800 1285.4600 1525.4800 1285.9400 ;
        RECT 1523.8800 1290.9000 1525.4800 1291.3800 ;
        RECT 1516.1200 1285.4600 1517.7200 1285.9400 ;
        RECT 1516.1200 1290.9000 1517.7200 1291.3800 ;
        RECT 1523.8800 1269.1400 1525.4800 1269.6200 ;
        RECT 1523.8800 1274.5800 1525.4800 1275.0600 ;
        RECT 1516.1200 1269.1400 1517.7200 1269.6200 ;
        RECT 1516.1200 1274.5800 1517.7200 1275.0600 ;
        RECT 1516.1200 1280.0200 1517.7200 1280.5000 ;
        RECT 1523.8800 1280.0200 1525.4800 1280.5000 ;
        RECT 1613.8800 1252.8200 1615.4800 1253.3000 ;
        RECT 1613.8800 1258.2600 1615.4800 1258.7400 ;
        RECT 1613.8800 1263.7000 1615.4800 1264.1800 ;
        RECT 1613.8800 1241.9400 1615.4800 1242.4200 ;
        RECT 1613.8800 1247.3800 1615.4800 1247.8600 ;
        RECT 1568.8800 1252.8200 1570.4800 1253.3000 ;
        RECT 1568.8800 1258.2600 1570.4800 1258.7400 ;
        RECT 1568.8800 1263.7000 1570.4800 1264.1800 ;
        RECT 1568.8800 1241.9400 1570.4800 1242.4200 ;
        RECT 1568.8800 1247.3800 1570.4800 1247.8600 ;
        RECT 1613.8800 1225.6200 1615.4800 1226.1000 ;
        RECT 1613.8800 1231.0600 1615.4800 1231.5400 ;
        RECT 1613.8800 1236.5000 1615.4800 1236.9800 ;
        RECT 1613.8800 1214.7400 1615.4800 1215.2200 ;
        RECT 1613.8800 1220.1800 1615.4800 1220.6600 ;
        RECT 1568.8800 1225.6200 1570.4800 1226.1000 ;
        RECT 1568.8800 1231.0600 1570.4800 1231.5400 ;
        RECT 1568.8800 1236.5000 1570.4800 1236.9800 ;
        RECT 1568.8800 1214.7400 1570.4800 1215.2200 ;
        RECT 1568.8800 1220.1800 1570.4800 1220.6600 ;
        RECT 1523.8800 1252.8200 1525.4800 1253.3000 ;
        RECT 1523.8800 1258.2600 1525.4800 1258.7400 ;
        RECT 1523.8800 1263.7000 1525.4800 1264.1800 ;
        RECT 1516.1200 1252.8200 1517.7200 1253.3000 ;
        RECT 1516.1200 1258.2600 1517.7200 1258.7400 ;
        RECT 1516.1200 1263.7000 1517.7200 1264.1800 ;
        RECT 1523.8800 1241.9400 1525.4800 1242.4200 ;
        RECT 1523.8800 1247.3800 1525.4800 1247.8600 ;
        RECT 1516.1200 1241.9400 1517.7200 1242.4200 ;
        RECT 1516.1200 1247.3800 1517.7200 1247.8600 ;
        RECT 1523.8800 1225.6200 1525.4800 1226.1000 ;
        RECT 1523.8800 1231.0600 1525.4800 1231.5400 ;
        RECT 1523.8800 1236.5000 1525.4800 1236.9800 ;
        RECT 1516.1200 1225.6200 1517.7200 1226.1000 ;
        RECT 1516.1200 1231.0600 1517.7200 1231.5400 ;
        RECT 1516.1200 1236.5000 1517.7200 1236.9800 ;
        RECT 1523.8800 1214.7400 1525.4800 1215.2200 ;
        RECT 1523.8800 1220.1800 1525.4800 1220.6600 ;
        RECT 1516.1200 1214.7400 1517.7200 1215.2200 ;
        RECT 1516.1200 1220.1800 1517.7200 1220.6600 ;
        RECT 1713.6200 1198.4200 1715.2200 1198.9000 ;
        RECT 1713.6200 1203.8600 1715.2200 1204.3400 ;
        RECT 1713.6200 1209.3000 1715.2200 1209.7800 ;
        RECT 1703.8800 1198.4200 1705.4800 1198.9000 ;
        RECT 1703.8800 1203.8600 1705.4800 1204.3400 ;
        RECT 1703.8800 1209.3000 1705.4800 1209.7800 ;
        RECT 1713.6200 1187.5400 1715.2200 1188.0200 ;
        RECT 1713.6200 1192.9800 1715.2200 1193.4600 ;
        RECT 1703.8800 1187.5400 1705.4800 1188.0200 ;
        RECT 1703.8800 1192.9800 1705.4800 1193.4600 ;
        RECT 1713.6200 1171.2200 1715.2200 1171.7000 ;
        RECT 1713.6200 1176.6600 1715.2200 1177.1400 ;
        RECT 1713.6200 1182.1000 1715.2200 1182.5800 ;
        RECT 1703.8800 1171.2200 1705.4800 1171.7000 ;
        RECT 1703.8800 1176.6600 1705.4800 1177.1400 ;
        RECT 1703.8800 1182.1000 1705.4800 1182.5800 ;
        RECT 1713.6200 1160.3400 1715.2200 1160.8200 ;
        RECT 1713.6200 1165.7800 1715.2200 1166.2600 ;
        RECT 1703.8800 1160.3400 1705.4800 1160.8200 ;
        RECT 1703.8800 1165.7800 1705.4800 1166.2600 ;
        RECT 1658.8800 1198.4200 1660.4800 1198.9000 ;
        RECT 1658.8800 1203.8600 1660.4800 1204.3400 ;
        RECT 1658.8800 1209.3000 1660.4800 1209.7800 ;
        RECT 1658.8800 1187.5400 1660.4800 1188.0200 ;
        RECT 1658.8800 1192.9800 1660.4800 1193.4600 ;
        RECT 1658.8800 1171.2200 1660.4800 1171.7000 ;
        RECT 1658.8800 1176.6600 1660.4800 1177.1400 ;
        RECT 1658.8800 1182.1000 1660.4800 1182.5800 ;
        RECT 1658.8800 1160.3400 1660.4800 1160.8200 ;
        RECT 1658.8800 1165.7800 1660.4800 1166.2600 ;
        RECT 1713.6200 1144.0200 1715.2200 1144.5000 ;
        RECT 1713.6200 1149.4600 1715.2200 1149.9400 ;
        RECT 1713.6200 1154.9000 1715.2200 1155.3800 ;
        RECT 1703.8800 1144.0200 1705.4800 1144.5000 ;
        RECT 1703.8800 1149.4600 1705.4800 1149.9400 ;
        RECT 1703.8800 1154.9000 1705.4800 1155.3800 ;
        RECT 1713.6200 1133.1400 1715.2200 1133.6200 ;
        RECT 1713.6200 1138.5800 1715.2200 1139.0600 ;
        RECT 1703.8800 1133.1400 1705.4800 1133.6200 ;
        RECT 1703.8800 1138.5800 1705.4800 1139.0600 ;
        RECT 1713.6200 1116.8200 1715.2200 1117.3000 ;
        RECT 1713.6200 1122.2600 1715.2200 1122.7400 ;
        RECT 1713.6200 1127.7000 1715.2200 1128.1800 ;
        RECT 1703.8800 1116.8200 1705.4800 1117.3000 ;
        RECT 1703.8800 1122.2600 1705.4800 1122.7400 ;
        RECT 1703.8800 1127.7000 1705.4800 1128.1800 ;
        RECT 1703.8800 1111.3800 1705.4800 1111.8600 ;
        RECT 1713.6200 1111.3800 1715.2200 1111.8600 ;
        RECT 1658.8800 1144.0200 1660.4800 1144.5000 ;
        RECT 1658.8800 1149.4600 1660.4800 1149.9400 ;
        RECT 1658.8800 1154.9000 1660.4800 1155.3800 ;
        RECT 1658.8800 1133.1400 1660.4800 1133.6200 ;
        RECT 1658.8800 1138.5800 1660.4800 1139.0600 ;
        RECT 1658.8800 1116.8200 1660.4800 1117.3000 ;
        RECT 1658.8800 1122.2600 1660.4800 1122.7400 ;
        RECT 1658.8800 1127.7000 1660.4800 1128.1800 ;
        RECT 1658.8800 1111.3800 1660.4800 1111.8600 ;
        RECT 1613.8800 1198.4200 1615.4800 1198.9000 ;
        RECT 1613.8800 1203.8600 1615.4800 1204.3400 ;
        RECT 1613.8800 1209.3000 1615.4800 1209.7800 ;
        RECT 1613.8800 1187.5400 1615.4800 1188.0200 ;
        RECT 1613.8800 1192.9800 1615.4800 1193.4600 ;
        RECT 1568.8800 1198.4200 1570.4800 1198.9000 ;
        RECT 1568.8800 1203.8600 1570.4800 1204.3400 ;
        RECT 1568.8800 1209.3000 1570.4800 1209.7800 ;
        RECT 1568.8800 1187.5400 1570.4800 1188.0200 ;
        RECT 1568.8800 1192.9800 1570.4800 1193.4600 ;
        RECT 1613.8800 1171.2200 1615.4800 1171.7000 ;
        RECT 1613.8800 1176.6600 1615.4800 1177.1400 ;
        RECT 1613.8800 1182.1000 1615.4800 1182.5800 ;
        RECT 1613.8800 1160.3400 1615.4800 1160.8200 ;
        RECT 1613.8800 1165.7800 1615.4800 1166.2600 ;
        RECT 1568.8800 1171.2200 1570.4800 1171.7000 ;
        RECT 1568.8800 1176.6600 1570.4800 1177.1400 ;
        RECT 1568.8800 1182.1000 1570.4800 1182.5800 ;
        RECT 1568.8800 1160.3400 1570.4800 1160.8200 ;
        RECT 1568.8800 1165.7800 1570.4800 1166.2600 ;
        RECT 1523.8800 1198.4200 1525.4800 1198.9000 ;
        RECT 1523.8800 1203.8600 1525.4800 1204.3400 ;
        RECT 1523.8800 1209.3000 1525.4800 1209.7800 ;
        RECT 1516.1200 1198.4200 1517.7200 1198.9000 ;
        RECT 1516.1200 1203.8600 1517.7200 1204.3400 ;
        RECT 1516.1200 1209.3000 1517.7200 1209.7800 ;
        RECT 1523.8800 1187.5400 1525.4800 1188.0200 ;
        RECT 1523.8800 1192.9800 1525.4800 1193.4600 ;
        RECT 1516.1200 1187.5400 1517.7200 1188.0200 ;
        RECT 1516.1200 1192.9800 1517.7200 1193.4600 ;
        RECT 1523.8800 1171.2200 1525.4800 1171.7000 ;
        RECT 1523.8800 1176.6600 1525.4800 1177.1400 ;
        RECT 1523.8800 1182.1000 1525.4800 1182.5800 ;
        RECT 1516.1200 1171.2200 1517.7200 1171.7000 ;
        RECT 1516.1200 1176.6600 1517.7200 1177.1400 ;
        RECT 1516.1200 1182.1000 1517.7200 1182.5800 ;
        RECT 1523.8800 1160.3400 1525.4800 1160.8200 ;
        RECT 1523.8800 1165.7800 1525.4800 1166.2600 ;
        RECT 1516.1200 1160.3400 1517.7200 1160.8200 ;
        RECT 1516.1200 1165.7800 1517.7200 1166.2600 ;
        RECT 1613.8800 1144.0200 1615.4800 1144.5000 ;
        RECT 1613.8800 1149.4600 1615.4800 1149.9400 ;
        RECT 1613.8800 1154.9000 1615.4800 1155.3800 ;
        RECT 1613.8800 1133.1400 1615.4800 1133.6200 ;
        RECT 1613.8800 1138.5800 1615.4800 1139.0600 ;
        RECT 1568.8800 1144.0200 1570.4800 1144.5000 ;
        RECT 1568.8800 1149.4600 1570.4800 1149.9400 ;
        RECT 1568.8800 1154.9000 1570.4800 1155.3800 ;
        RECT 1568.8800 1133.1400 1570.4800 1133.6200 ;
        RECT 1568.8800 1138.5800 1570.4800 1139.0600 ;
        RECT 1613.8800 1116.8200 1615.4800 1117.3000 ;
        RECT 1613.8800 1122.2600 1615.4800 1122.7400 ;
        RECT 1613.8800 1127.7000 1615.4800 1128.1800 ;
        RECT 1613.8800 1111.3800 1615.4800 1111.8600 ;
        RECT 1568.8800 1116.8200 1570.4800 1117.3000 ;
        RECT 1568.8800 1122.2600 1570.4800 1122.7400 ;
        RECT 1568.8800 1127.7000 1570.4800 1128.1800 ;
        RECT 1568.8800 1111.3800 1570.4800 1111.8600 ;
        RECT 1523.8800 1144.0200 1525.4800 1144.5000 ;
        RECT 1523.8800 1149.4600 1525.4800 1149.9400 ;
        RECT 1523.8800 1154.9000 1525.4800 1155.3800 ;
        RECT 1516.1200 1144.0200 1517.7200 1144.5000 ;
        RECT 1516.1200 1149.4600 1517.7200 1149.9400 ;
        RECT 1516.1200 1154.9000 1517.7200 1155.3800 ;
        RECT 1523.8800 1133.1400 1525.4800 1133.6200 ;
        RECT 1523.8800 1138.5800 1525.4800 1139.0600 ;
        RECT 1516.1200 1133.1400 1517.7200 1133.6200 ;
        RECT 1516.1200 1138.5800 1517.7200 1139.0600 ;
        RECT 1523.8800 1116.8200 1525.4800 1117.3000 ;
        RECT 1523.8800 1122.2600 1525.4800 1122.7400 ;
        RECT 1523.8800 1127.7000 1525.4800 1128.1800 ;
        RECT 1516.1200 1116.8200 1517.7200 1117.3000 ;
        RECT 1516.1200 1122.2600 1517.7200 1122.7400 ;
        RECT 1516.1200 1127.7000 1517.7200 1128.1800 ;
        RECT 1516.1200 1111.3800 1517.7200 1111.8600 ;
        RECT 1523.8800 1111.3800 1525.4800 1111.8600 ;
        RECT 1510.5600 1313.6900 1720.7800 1315.2900 ;
        RECT 1510.5600 1107.1900 1720.7800 1108.7900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1101.7600 1517.7200 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1319.8000 1517.7200 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1101.7600 1715.2200 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1319.8000 1715.2200 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1107.1900 1512.1600 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1107.1900 1720.7800 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1313.6900 1512.1600 1315.2900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1313.6900 1720.7800 1315.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 877.5500 1705.4800 1085.6500 ;
        RECT 1658.8800 877.5500 1660.4800 1085.6500 ;
        RECT 1613.8800 877.5500 1615.4800 1085.6500 ;
        RECT 1568.8800 877.5500 1570.4800 1085.6500 ;
        RECT 1523.8800 877.5500 1525.4800 1085.6500 ;
        RECT 1713.6200 872.1200 1715.2200 1091.7600 ;
        RECT 1516.1200 872.1200 1517.7200 1091.7600 ;
      LAYER met3 ;
        RECT 1713.6200 1066.7000 1715.2200 1067.1800 ;
        RECT 1713.6200 1072.1400 1715.2200 1072.6200 ;
        RECT 1703.8800 1066.7000 1705.4800 1067.1800 ;
        RECT 1703.8800 1072.1400 1705.4800 1072.6200 ;
        RECT 1703.8800 1077.5800 1705.4800 1078.0600 ;
        RECT 1713.6200 1077.5800 1715.2200 1078.0600 ;
        RECT 1713.6200 1055.8200 1715.2200 1056.3000 ;
        RECT 1713.6200 1061.2600 1715.2200 1061.7400 ;
        RECT 1703.8800 1055.8200 1705.4800 1056.3000 ;
        RECT 1703.8800 1061.2600 1705.4800 1061.7400 ;
        RECT 1713.6200 1039.5000 1715.2200 1039.9800 ;
        RECT 1713.6200 1044.9400 1715.2200 1045.4200 ;
        RECT 1703.8800 1039.5000 1705.4800 1039.9800 ;
        RECT 1703.8800 1044.9400 1705.4800 1045.4200 ;
        RECT 1703.8800 1050.3800 1705.4800 1050.8600 ;
        RECT 1713.6200 1050.3800 1715.2200 1050.8600 ;
        RECT 1658.8800 1066.7000 1660.4800 1067.1800 ;
        RECT 1658.8800 1072.1400 1660.4800 1072.6200 ;
        RECT 1658.8800 1077.5800 1660.4800 1078.0600 ;
        RECT 1658.8800 1055.8200 1660.4800 1056.3000 ;
        RECT 1658.8800 1061.2600 1660.4800 1061.7400 ;
        RECT 1658.8800 1039.5000 1660.4800 1039.9800 ;
        RECT 1658.8800 1044.9400 1660.4800 1045.4200 ;
        RECT 1658.8800 1050.3800 1660.4800 1050.8600 ;
        RECT 1713.6200 1023.1800 1715.2200 1023.6600 ;
        RECT 1713.6200 1028.6200 1715.2200 1029.1000 ;
        RECT 1713.6200 1034.0600 1715.2200 1034.5400 ;
        RECT 1703.8800 1023.1800 1705.4800 1023.6600 ;
        RECT 1703.8800 1028.6200 1705.4800 1029.1000 ;
        RECT 1703.8800 1034.0600 1705.4800 1034.5400 ;
        RECT 1713.6200 1012.3000 1715.2200 1012.7800 ;
        RECT 1713.6200 1017.7400 1715.2200 1018.2200 ;
        RECT 1703.8800 1012.3000 1705.4800 1012.7800 ;
        RECT 1703.8800 1017.7400 1705.4800 1018.2200 ;
        RECT 1713.6200 995.9800 1715.2200 996.4600 ;
        RECT 1713.6200 1001.4200 1715.2200 1001.9000 ;
        RECT 1713.6200 1006.8600 1715.2200 1007.3400 ;
        RECT 1703.8800 995.9800 1705.4800 996.4600 ;
        RECT 1703.8800 1001.4200 1705.4800 1001.9000 ;
        RECT 1703.8800 1006.8600 1705.4800 1007.3400 ;
        RECT 1713.6200 985.1000 1715.2200 985.5800 ;
        RECT 1713.6200 990.5400 1715.2200 991.0200 ;
        RECT 1703.8800 985.1000 1705.4800 985.5800 ;
        RECT 1703.8800 990.5400 1705.4800 991.0200 ;
        RECT 1658.8800 1023.1800 1660.4800 1023.6600 ;
        RECT 1658.8800 1028.6200 1660.4800 1029.1000 ;
        RECT 1658.8800 1034.0600 1660.4800 1034.5400 ;
        RECT 1658.8800 1012.3000 1660.4800 1012.7800 ;
        RECT 1658.8800 1017.7400 1660.4800 1018.2200 ;
        RECT 1658.8800 995.9800 1660.4800 996.4600 ;
        RECT 1658.8800 1001.4200 1660.4800 1001.9000 ;
        RECT 1658.8800 1006.8600 1660.4800 1007.3400 ;
        RECT 1658.8800 985.1000 1660.4800 985.5800 ;
        RECT 1658.8800 990.5400 1660.4800 991.0200 ;
        RECT 1613.8800 1066.7000 1615.4800 1067.1800 ;
        RECT 1613.8800 1072.1400 1615.4800 1072.6200 ;
        RECT 1613.8800 1077.5800 1615.4800 1078.0600 ;
        RECT 1568.8800 1066.7000 1570.4800 1067.1800 ;
        RECT 1568.8800 1072.1400 1570.4800 1072.6200 ;
        RECT 1568.8800 1077.5800 1570.4800 1078.0600 ;
        RECT 1613.8800 1055.8200 1615.4800 1056.3000 ;
        RECT 1613.8800 1061.2600 1615.4800 1061.7400 ;
        RECT 1613.8800 1039.5000 1615.4800 1039.9800 ;
        RECT 1613.8800 1044.9400 1615.4800 1045.4200 ;
        RECT 1613.8800 1050.3800 1615.4800 1050.8600 ;
        RECT 1568.8800 1055.8200 1570.4800 1056.3000 ;
        RECT 1568.8800 1061.2600 1570.4800 1061.7400 ;
        RECT 1568.8800 1039.5000 1570.4800 1039.9800 ;
        RECT 1568.8800 1044.9400 1570.4800 1045.4200 ;
        RECT 1568.8800 1050.3800 1570.4800 1050.8600 ;
        RECT 1523.8800 1066.7000 1525.4800 1067.1800 ;
        RECT 1523.8800 1072.1400 1525.4800 1072.6200 ;
        RECT 1516.1200 1066.7000 1517.7200 1067.1800 ;
        RECT 1516.1200 1072.1400 1517.7200 1072.6200 ;
        RECT 1516.1200 1077.5800 1517.7200 1078.0600 ;
        RECT 1523.8800 1077.5800 1525.4800 1078.0600 ;
        RECT 1523.8800 1055.8200 1525.4800 1056.3000 ;
        RECT 1523.8800 1061.2600 1525.4800 1061.7400 ;
        RECT 1516.1200 1055.8200 1517.7200 1056.3000 ;
        RECT 1516.1200 1061.2600 1517.7200 1061.7400 ;
        RECT 1523.8800 1039.5000 1525.4800 1039.9800 ;
        RECT 1523.8800 1044.9400 1525.4800 1045.4200 ;
        RECT 1516.1200 1039.5000 1517.7200 1039.9800 ;
        RECT 1516.1200 1044.9400 1517.7200 1045.4200 ;
        RECT 1516.1200 1050.3800 1517.7200 1050.8600 ;
        RECT 1523.8800 1050.3800 1525.4800 1050.8600 ;
        RECT 1613.8800 1023.1800 1615.4800 1023.6600 ;
        RECT 1613.8800 1028.6200 1615.4800 1029.1000 ;
        RECT 1613.8800 1034.0600 1615.4800 1034.5400 ;
        RECT 1613.8800 1012.3000 1615.4800 1012.7800 ;
        RECT 1613.8800 1017.7400 1615.4800 1018.2200 ;
        RECT 1568.8800 1023.1800 1570.4800 1023.6600 ;
        RECT 1568.8800 1028.6200 1570.4800 1029.1000 ;
        RECT 1568.8800 1034.0600 1570.4800 1034.5400 ;
        RECT 1568.8800 1012.3000 1570.4800 1012.7800 ;
        RECT 1568.8800 1017.7400 1570.4800 1018.2200 ;
        RECT 1613.8800 995.9800 1615.4800 996.4600 ;
        RECT 1613.8800 1001.4200 1615.4800 1001.9000 ;
        RECT 1613.8800 1006.8600 1615.4800 1007.3400 ;
        RECT 1613.8800 985.1000 1615.4800 985.5800 ;
        RECT 1613.8800 990.5400 1615.4800 991.0200 ;
        RECT 1568.8800 995.9800 1570.4800 996.4600 ;
        RECT 1568.8800 1001.4200 1570.4800 1001.9000 ;
        RECT 1568.8800 1006.8600 1570.4800 1007.3400 ;
        RECT 1568.8800 985.1000 1570.4800 985.5800 ;
        RECT 1568.8800 990.5400 1570.4800 991.0200 ;
        RECT 1523.8800 1023.1800 1525.4800 1023.6600 ;
        RECT 1523.8800 1028.6200 1525.4800 1029.1000 ;
        RECT 1523.8800 1034.0600 1525.4800 1034.5400 ;
        RECT 1516.1200 1023.1800 1517.7200 1023.6600 ;
        RECT 1516.1200 1028.6200 1517.7200 1029.1000 ;
        RECT 1516.1200 1034.0600 1517.7200 1034.5400 ;
        RECT 1523.8800 1012.3000 1525.4800 1012.7800 ;
        RECT 1523.8800 1017.7400 1525.4800 1018.2200 ;
        RECT 1516.1200 1012.3000 1517.7200 1012.7800 ;
        RECT 1516.1200 1017.7400 1517.7200 1018.2200 ;
        RECT 1523.8800 995.9800 1525.4800 996.4600 ;
        RECT 1523.8800 1001.4200 1525.4800 1001.9000 ;
        RECT 1523.8800 1006.8600 1525.4800 1007.3400 ;
        RECT 1516.1200 995.9800 1517.7200 996.4600 ;
        RECT 1516.1200 1001.4200 1517.7200 1001.9000 ;
        RECT 1516.1200 1006.8600 1517.7200 1007.3400 ;
        RECT 1523.8800 985.1000 1525.4800 985.5800 ;
        RECT 1523.8800 990.5400 1525.4800 991.0200 ;
        RECT 1516.1200 985.1000 1517.7200 985.5800 ;
        RECT 1516.1200 990.5400 1517.7200 991.0200 ;
        RECT 1713.6200 968.7800 1715.2200 969.2600 ;
        RECT 1713.6200 974.2200 1715.2200 974.7000 ;
        RECT 1713.6200 979.6600 1715.2200 980.1400 ;
        RECT 1703.8800 968.7800 1705.4800 969.2600 ;
        RECT 1703.8800 974.2200 1705.4800 974.7000 ;
        RECT 1703.8800 979.6600 1705.4800 980.1400 ;
        RECT 1713.6200 957.9000 1715.2200 958.3800 ;
        RECT 1713.6200 963.3400 1715.2200 963.8200 ;
        RECT 1703.8800 957.9000 1705.4800 958.3800 ;
        RECT 1703.8800 963.3400 1705.4800 963.8200 ;
        RECT 1713.6200 941.5800 1715.2200 942.0600 ;
        RECT 1713.6200 947.0200 1715.2200 947.5000 ;
        RECT 1713.6200 952.4600 1715.2200 952.9400 ;
        RECT 1703.8800 941.5800 1705.4800 942.0600 ;
        RECT 1703.8800 947.0200 1705.4800 947.5000 ;
        RECT 1703.8800 952.4600 1705.4800 952.9400 ;
        RECT 1713.6200 930.7000 1715.2200 931.1800 ;
        RECT 1713.6200 936.1400 1715.2200 936.6200 ;
        RECT 1703.8800 930.7000 1705.4800 931.1800 ;
        RECT 1703.8800 936.1400 1705.4800 936.6200 ;
        RECT 1658.8800 968.7800 1660.4800 969.2600 ;
        RECT 1658.8800 974.2200 1660.4800 974.7000 ;
        RECT 1658.8800 979.6600 1660.4800 980.1400 ;
        RECT 1658.8800 957.9000 1660.4800 958.3800 ;
        RECT 1658.8800 963.3400 1660.4800 963.8200 ;
        RECT 1658.8800 941.5800 1660.4800 942.0600 ;
        RECT 1658.8800 947.0200 1660.4800 947.5000 ;
        RECT 1658.8800 952.4600 1660.4800 952.9400 ;
        RECT 1658.8800 930.7000 1660.4800 931.1800 ;
        RECT 1658.8800 936.1400 1660.4800 936.6200 ;
        RECT 1713.6200 914.3800 1715.2200 914.8600 ;
        RECT 1713.6200 919.8200 1715.2200 920.3000 ;
        RECT 1713.6200 925.2600 1715.2200 925.7400 ;
        RECT 1703.8800 914.3800 1705.4800 914.8600 ;
        RECT 1703.8800 919.8200 1705.4800 920.3000 ;
        RECT 1703.8800 925.2600 1705.4800 925.7400 ;
        RECT 1713.6200 903.5000 1715.2200 903.9800 ;
        RECT 1713.6200 908.9400 1715.2200 909.4200 ;
        RECT 1703.8800 903.5000 1705.4800 903.9800 ;
        RECT 1703.8800 908.9400 1705.4800 909.4200 ;
        RECT 1713.6200 887.1800 1715.2200 887.6600 ;
        RECT 1713.6200 892.6200 1715.2200 893.1000 ;
        RECT 1713.6200 898.0600 1715.2200 898.5400 ;
        RECT 1703.8800 887.1800 1705.4800 887.6600 ;
        RECT 1703.8800 892.6200 1705.4800 893.1000 ;
        RECT 1703.8800 898.0600 1705.4800 898.5400 ;
        RECT 1703.8800 881.7400 1705.4800 882.2200 ;
        RECT 1713.6200 881.7400 1715.2200 882.2200 ;
        RECT 1658.8800 914.3800 1660.4800 914.8600 ;
        RECT 1658.8800 919.8200 1660.4800 920.3000 ;
        RECT 1658.8800 925.2600 1660.4800 925.7400 ;
        RECT 1658.8800 903.5000 1660.4800 903.9800 ;
        RECT 1658.8800 908.9400 1660.4800 909.4200 ;
        RECT 1658.8800 887.1800 1660.4800 887.6600 ;
        RECT 1658.8800 892.6200 1660.4800 893.1000 ;
        RECT 1658.8800 898.0600 1660.4800 898.5400 ;
        RECT 1658.8800 881.7400 1660.4800 882.2200 ;
        RECT 1613.8800 968.7800 1615.4800 969.2600 ;
        RECT 1613.8800 974.2200 1615.4800 974.7000 ;
        RECT 1613.8800 979.6600 1615.4800 980.1400 ;
        RECT 1613.8800 957.9000 1615.4800 958.3800 ;
        RECT 1613.8800 963.3400 1615.4800 963.8200 ;
        RECT 1568.8800 968.7800 1570.4800 969.2600 ;
        RECT 1568.8800 974.2200 1570.4800 974.7000 ;
        RECT 1568.8800 979.6600 1570.4800 980.1400 ;
        RECT 1568.8800 957.9000 1570.4800 958.3800 ;
        RECT 1568.8800 963.3400 1570.4800 963.8200 ;
        RECT 1613.8800 941.5800 1615.4800 942.0600 ;
        RECT 1613.8800 947.0200 1615.4800 947.5000 ;
        RECT 1613.8800 952.4600 1615.4800 952.9400 ;
        RECT 1613.8800 930.7000 1615.4800 931.1800 ;
        RECT 1613.8800 936.1400 1615.4800 936.6200 ;
        RECT 1568.8800 941.5800 1570.4800 942.0600 ;
        RECT 1568.8800 947.0200 1570.4800 947.5000 ;
        RECT 1568.8800 952.4600 1570.4800 952.9400 ;
        RECT 1568.8800 930.7000 1570.4800 931.1800 ;
        RECT 1568.8800 936.1400 1570.4800 936.6200 ;
        RECT 1523.8800 968.7800 1525.4800 969.2600 ;
        RECT 1523.8800 974.2200 1525.4800 974.7000 ;
        RECT 1523.8800 979.6600 1525.4800 980.1400 ;
        RECT 1516.1200 968.7800 1517.7200 969.2600 ;
        RECT 1516.1200 974.2200 1517.7200 974.7000 ;
        RECT 1516.1200 979.6600 1517.7200 980.1400 ;
        RECT 1523.8800 957.9000 1525.4800 958.3800 ;
        RECT 1523.8800 963.3400 1525.4800 963.8200 ;
        RECT 1516.1200 957.9000 1517.7200 958.3800 ;
        RECT 1516.1200 963.3400 1517.7200 963.8200 ;
        RECT 1523.8800 941.5800 1525.4800 942.0600 ;
        RECT 1523.8800 947.0200 1525.4800 947.5000 ;
        RECT 1523.8800 952.4600 1525.4800 952.9400 ;
        RECT 1516.1200 941.5800 1517.7200 942.0600 ;
        RECT 1516.1200 947.0200 1517.7200 947.5000 ;
        RECT 1516.1200 952.4600 1517.7200 952.9400 ;
        RECT 1523.8800 930.7000 1525.4800 931.1800 ;
        RECT 1523.8800 936.1400 1525.4800 936.6200 ;
        RECT 1516.1200 930.7000 1517.7200 931.1800 ;
        RECT 1516.1200 936.1400 1517.7200 936.6200 ;
        RECT 1613.8800 914.3800 1615.4800 914.8600 ;
        RECT 1613.8800 919.8200 1615.4800 920.3000 ;
        RECT 1613.8800 925.2600 1615.4800 925.7400 ;
        RECT 1613.8800 903.5000 1615.4800 903.9800 ;
        RECT 1613.8800 908.9400 1615.4800 909.4200 ;
        RECT 1568.8800 914.3800 1570.4800 914.8600 ;
        RECT 1568.8800 919.8200 1570.4800 920.3000 ;
        RECT 1568.8800 925.2600 1570.4800 925.7400 ;
        RECT 1568.8800 903.5000 1570.4800 903.9800 ;
        RECT 1568.8800 908.9400 1570.4800 909.4200 ;
        RECT 1613.8800 887.1800 1615.4800 887.6600 ;
        RECT 1613.8800 892.6200 1615.4800 893.1000 ;
        RECT 1613.8800 898.0600 1615.4800 898.5400 ;
        RECT 1613.8800 881.7400 1615.4800 882.2200 ;
        RECT 1568.8800 887.1800 1570.4800 887.6600 ;
        RECT 1568.8800 892.6200 1570.4800 893.1000 ;
        RECT 1568.8800 898.0600 1570.4800 898.5400 ;
        RECT 1568.8800 881.7400 1570.4800 882.2200 ;
        RECT 1523.8800 914.3800 1525.4800 914.8600 ;
        RECT 1523.8800 919.8200 1525.4800 920.3000 ;
        RECT 1523.8800 925.2600 1525.4800 925.7400 ;
        RECT 1516.1200 914.3800 1517.7200 914.8600 ;
        RECT 1516.1200 919.8200 1517.7200 920.3000 ;
        RECT 1516.1200 925.2600 1517.7200 925.7400 ;
        RECT 1523.8800 903.5000 1525.4800 903.9800 ;
        RECT 1523.8800 908.9400 1525.4800 909.4200 ;
        RECT 1516.1200 903.5000 1517.7200 903.9800 ;
        RECT 1516.1200 908.9400 1517.7200 909.4200 ;
        RECT 1523.8800 887.1800 1525.4800 887.6600 ;
        RECT 1523.8800 892.6200 1525.4800 893.1000 ;
        RECT 1523.8800 898.0600 1525.4800 898.5400 ;
        RECT 1516.1200 887.1800 1517.7200 887.6600 ;
        RECT 1516.1200 892.6200 1517.7200 893.1000 ;
        RECT 1516.1200 898.0600 1517.7200 898.5400 ;
        RECT 1516.1200 881.7400 1517.7200 882.2200 ;
        RECT 1523.8800 881.7400 1525.4800 882.2200 ;
        RECT 1510.5600 1084.0500 1720.7800 1085.6500 ;
        RECT 1510.5600 877.5500 1720.7800 879.1500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 872.1200 1517.7200 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 1090.1600 1517.7200 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 872.1200 1715.2200 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 1090.1600 1715.2200 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 877.5500 1512.1600 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 877.5500 1720.7800 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 1084.0500 1512.1600 1085.6500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 1084.0500 1720.7800 1085.6500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 647.9100 1705.4800 856.0100 ;
        RECT 1658.8800 647.9100 1660.4800 856.0100 ;
        RECT 1613.8800 647.9100 1615.4800 856.0100 ;
        RECT 1568.8800 647.9100 1570.4800 856.0100 ;
        RECT 1523.8800 647.9100 1525.4800 856.0100 ;
        RECT 1713.6200 642.4800 1715.2200 862.1200 ;
        RECT 1516.1200 642.4800 1517.7200 862.1200 ;
      LAYER met3 ;
        RECT 1713.6200 837.0600 1715.2200 837.5400 ;
        RECT 1713.6200 842.5000 1715.2200 842.9800 ;
        RECT 1703.8800 837.0600 1705.4800 837.5400 ;
        RECT 1703.8800 842.5000 1705.4800 842.9800 ;
        RECT 1703.8800 847.9400 1705.4800 848.4200 ;
        RECT 1713.6200 847.9400 1715.2200 848.4200 ;
        RECT 1713.6200 826.1800 1715.2200 826.6600 ;
        RECT 1713.6200 831.6200 1715.2200 832.1000 ;
        RECT 1703.8800 826.1800 1705.4800 826.6600 ;
        RECT 1703.8800 831.6200 1705.4800 832.1000 ;
        RECT 1713.6200 809.8600 1715.2200 810.3400 ;
        RECT 1713.6200 815.3000 1715.2200 815.7800 ;
        RECT 1703.8800 809.8600 1705.4800 810.3400 ;
        RECT 1703.8800 815.3000 1705.4800 815.7800 ;
        RECT 1703.8800 820.7400 1705.4800 821.2200 ;
        RECT 1713.6200 820.7400 1715.2200 821.2200 ;
        RECT 1658.8800 837.0600 1660.4800 837.5400 ;
        RECT 1658.8800 842.5000 1660.4800 842.9800 ;
        RECT 1658.8800 847.9400 1660.4800 848.4200 ;
        RECT 1658.8800 826.1800 1660.4800 826.6600 ;
        RECT 1658.8800 831.6200 1660.4800 832.1000 ;
        RECT 1658.8800 809.8600 1660.4800 810.3400 ;
        RECT 1658.8800 815.3000 1660.4800 815.7800 ;
        RECT 1658.8800 820.7400 1660.4800 821.2200 ;
        RECT 1713.6200 793.5400 1715.2200 794.0200 ;
        RECT 1713.6200 798.9800 1715.2200 799.4600 ;
        RECT 1713.6200 804.4200 1715.2200 804.9000 ;
        RECT 1703.8800 793.5400 1705.4800 794.0200 ;
        RECT 1703.8800 798.9800 1705.4800 799.4600 ;
        RECT 1703.8800 804.4200 1705.4800 804.9000 ;
        RECT 1713.6200 782.6600 1715.2200 783.1400 ;
        RECT 1713.6200 788.1000 1715.2200 788.5800 ;
        RECT 1703.8800 782.6600 1705.4800 783.1400 ;
        RECT 1703.8800 788.1000 1705.4800 788.5800 ;
        RECT 1713.6200 766.3400 1715.2200 766.8200 ;
        RECT 1713.6200 771.7800 1715.2200 772.2600 ;
        RECT 1713.6200 777.2200 1715.2200 777.7000 ;
        RECT 1703.8800 766.3400 1705.4800 766.8200 ;
        RECT 1703.8800 771.7800 1705.4800 772.2600 ;
        RECT 1703.8800 777.2200 1705.4800 777.7000 ;
        RECT 1713.6200 755.4600 1715.2200 755.9400 ;
        RECT 1713.6200 760.9000 1715.2200 761.3800 ;
        RECT 1703.8800 755.4600 1705.4800 755.9400 ;
        RECT 1703.8800 760.9000 1705.4800 761.3800 ;
        RECT 1658.8800 793.5400 1660.4800 794.0200 ;
        RECT 1658.8800 798.9800 1660.4800 799.4600 ;
        RECT 1658.8800 804.4200 1660.4800 804.9000 ;
        RECT 1658.8800 782.6600 1660.4800 783.1400 ;
        RECT 1658.8800 788.1000 1660.4800 788.5800 ;
        RECT 1658.8800 766.3400 1660.4800 766.8200 ;
        RECT 1658.8800 771.7800 1660.4800 772.2600 ;
        RECT 1658.8800 777.2200 1660.4800 777.7000 ;
        RECT 1658.8800 755.4600 1660.4800 755.9400 ;
        RECT 1658.8800 760.9000 1660.4800 761.3800 ;
        RECT 1613.8800 837.0600 1615.4800 837.5400 ;
        RECT 1613.8800 842.5000 1615.4800 842.9800 ;
        RECT 1613.8800 847.9400 1615.4800 848.4200 ;
        RECT 1568.8800 837.0600 1570.4800 837.5400 ;
        RECT 1568.8800 842.5000 1570.4800 842.9800 ;
        RECT 1568.8800 847.9400 1570.4800 848.4200 ;
        RECT 1613.8800 826.1800 1615.4800 826.6600 ;
        RECT 1613.8800 831.6200 1615.4800 832.1000 ;
        RECT 1613.8800 809.8600 1615.4800 810.3400 ;
        RECT 1613.8800 815.3000 1615.4800 815.7800 ;
        RECT 1613.8800 820.7400 1615.4800 821.2200 ;
        RECT 1568.8800 826.1800 1570.4800 826.6600 ;
        RECT 1568.8800 831.6200 1570.4800 832.1000 ;
        RECT 1568.8800 809.8600 1570.4800 810.3400 ;
        RECT 1568.8800 815.3000 1570.4800 815.7800 ;
        RECT 1568.8800 820.7400 1570.4800 821.2200 ;
        RECT 1523.8800 837.0600 1525.4800 837.5400 ;
        RECT 1523.8800 842.5000 1525.4800 842.9800 ;
        RECT 1516.1200 837.0600 1517.7200 837.5400 ;
        RECT 1516.1200 842.5000 1517.7200 842.9800 ;
        RECT 1516.1200 847.9400 1517.7200 848.4200 ;
        RECT 1523.8800 847.9400 1525.4800 848.4200 ;
        RECT 1523.8800 826.1800 1525.4800 826.6600 ;
        RECT 1523.8800 831.6200 1525.4800 832.1000 ;
        RECT 1516.1200 826.1800 1517.7200 826.6600 ;
        RECT 1516.1200 831.6200 1517.7200 832.1000 ;
        RECT 1523.8800 809.8600 1525.4800 810.3400 ;
        RECT 1523.8800 815.3000 1525.4800 815.7800 ;
        RECT 1516.1200 809.8600 1517.7200 810.3400 ;
        RECT 1516.1200 815.3000 1517.7200 815.7800 ;
        RECT 1516.1200 820.7400 1517.7200 821.2200 ;
        RECT 1523.8800 820.7400 1525.4800 821.2200 ;
        RECT 1613.8800 793.5400 1615.4800 794.0200 ;
        RECT 1613.8800 798.9800 1615.4800 799.4600 ;
        RECT 1613.8800 804.4200 1615.4800 804.9000 ;
        RECT 1613.8800 782.6600 1615.4800 783.1400 ;
        RECT 1613.8800 788.1000 1615.4800 788.5800 ;
        RECT 1568.8800 793.5400 1570.4800 794.0200 ;
        RECT 1568.8800 798.9800 1570.4800 799.4600 ;
        RECT 1568.8800 804.4200 1570.4800 804.9000 ;
        RECT 1568.8800 782.6600 1570.4800 783.1400 ;
        RECT 1568.8800 788.1000 1570.4800 788.5800 ;
        RECT 1613.8800 766.3400 1615.4800 766.8200 ;
        RECT 1613.8800 771.7800 1615.4800 772.2600 ;
        RECT 1613.8800 777.2200 1615.4800 777.7000 ;
        RECT 1613.8800 755.4600 1615.4800 755.9400 ;
        RECT 1613.8800 760.9000 1615.4800 761.3800 ;
        RECT 1568.8800 766.3400 1570.4800 766.8200 ;
        RECT 1568.8800 771.7800 1570.4800 772.2600 ;
        RECT 1568.8800 777.2200 1570.4800 777.7000 ;
        RECT 1568.8800 755.4600 1570.4800 755.9400 ;
        RECT 1568.8800 760.9000 1570.4800 761.3800 ;
        RECT 1523.8800 793.5400 1525.4800 794.0200 ;
        RECT 1523.8800 798.9800 1525.4800 799.4600 ;
        RECT 1523.8800 804.4200 1525.4800 804.9000 ;
        RECT 1516.1200 793.5400 1517.7200 794.0200 ;
        RECT 1516.1200 798.9800 1517.7200 799.4600 ;
        RECT 1516.1200 804.4200 1517.7200 804.9000 ;
        RECT 1523.8800 782.6600 1525.4800 783.1400 ;
        RECT 1523.8800 788.1000 1525.4800 788.5800 ;
        RECT 1516.1200 782.6600 1517.7200 783.1400 ;
        RECT 1516.1200 788.1000 1517.7200 788.5800 ;
        RECT 1523.8800 766.3400 1525.4800 766.8200 ;
        RECT 1523.8800 771.7800 1525.4800 772.2600 ;
        RECT 1523.8800 777.2200 1525.4800 777.7000 ;
        RECT 1516.1200 766.3400 1517.7200 766.8200 ;
        RECT 1516.1200 771.7800 1517.7200 772.2600 ;
        RECT 1516.1200 777.2200 1517.7200 777.7000 ;
        RECT 1523.8800 755.4600 1525.4800 755.9400 ;
        RECT 1523.8800 760.9000 1525.4800 761.3800 ;
        RECT 1516.1200 755.4600 1517.7200 755.9400 ;
        RECT 1516.1200 760.9000 1517.7200 761.3800 ;
        RECT 1713.6200 739.1400 1715.2200 739.6200 ;
        RECT 1713.6200 744.5800 1715.2200 745.0600 ;
        RECT 1713.6200 750.0200 1715.2200 750.5000 ;
        RECT 1703.8800 739.1400 1705.4800 739.6200 ;
        RECT 1703.8800 744.5800 1705.4800 745.0600 ;
        RECT 1703.8800 750.0200 1705.4800 750.5000 ;
        RECT 1713.6200 728.2600 1715.2200 728.7400 ;
        RECT 1713.6200 733.7000 1715.2200 734.1800 ;
        RECT 1703.8800 728.2600 1705.4800 728.7400 ;
        RECT 1703.8800 733.7000 1705.4800 734.1800 ;
        RECT 1713.6200 711.9400 1715.2200 712.4200 ;
        RECT 1713.6200 717.3800 1715.2200 717.8600 ;
        RECT 1713.6200 722.8200 1715.2200 723.3000 ;
        RECT 1703.8800 711.9400 1705.4800 712.4200 ;
        RECT 1703.8800 717.3800 1705.4800 717.8600 ;
        RECT 1703.8800 722.8200 1705.4800 723.3000 ;
        RECT 1713.6200 701.0600 1715.2200 701.5400 ;
        RECT 1713.6200 706.5000 1715.2200 706.9800 ;
        RECT 1703.8800 701.0600 1705.4800 701.5400 ;
        RECT 1703.8800 706.5000 1705.4800 706.9800 ;
        RECT 1658.8800 739.1400 1660.4800 739.6200 ;
        RECT 1658.8800 744.5800 1660.4800 745.0600 ;
        RECT 1658.8800 750.0200 1660.4800 750.5000 ;
        RECT 1658.8800 728.2600 1660.4800 728.7400 ;
        RECT 1658.8800 733.7000 1660.4800 734.1800 ;
        RECT 1658.8800 711.9400 1660.4800 712.4200 ;
        RECT 1658.8800 717.3800 1660.4800 717.8600 ;
        RECT 1658.8800 722.8200 1660.4800 723.3000 ;
        RECT 1658.8800 701.0600 1660.4800 701.5400 ;
        RECT 1658.8800 706.5000 1660.4800 706.9800 ;
        RECT 1713.6200 684.7400 1715.2200 685.2200 ;
        RECT 1713.6200 690.1800 1715.2200 690.6600 ;
        RECT 1713.6200 695.6200 1715.2200 696.1000 ;
        RECT 1703.8800 684.7400 1705.4800 685.2200 ;
        RECT 1703.8800 690.1800 1705.4800 690.6600 ;
        RECT 1703.8800 695.6200 1705.4800 696.1000 ;
        RECT 1713.6200 673.8600 1715.2200 674.3400 ;
        RECT 1713.6200 679.3000 1715.2200 679.7800 ;
        RECT 1703.8800 673.8600 1705.4800 674.3400 ;
        RECT 1703.8800 679.3000 1705.4800 679.7800 ;
        RECT 1713.6200 657.5400 1715.2200 658.0200 ;
        RECT 1713.6200 662.9800 1715.2200 663.4600 ;
        RECT 1713.6200 668.4200 1715.2200 668.9000 ;
        RECT 1703.8800 657.5400 1705.4800 658.0200 ;
        RECT 1703.8800 662.9800 1705.4800 663.4600 ;
        RECT 1703.8800 668.4200 1705.4800 668.9000 ;
        RECT 1703.8800 652.1000 1705.4800 652.5800 ;
        RECT 1713.6200 652.1000 1715.2200 652.5800 ;
        RECT 1658.8800 684.7400 1660.4800 685.2200 ;
        RECT 1658.8800 690.1800 1660.4800 690.6600 ;
        RECT 1658.8800 695.6200 1660.4800 696.1000 ;
        RECT 1658.8800 673.8600 1660.4800 674.3400 ;
        RECT 1658.8800 679.3000 1660.4800 679.7800 ;
        RECT 1658.8800 657.5400 1660.4800 658.0200 ;
        RECT 1658.8800 662.9800 1660.4800 663.4600 ;
        RECT 1658.8800 668.4200 1660.4800 668.9000 ;
        RECT 1658.8800 652.1000 1660.4800 652.5800 ;
        RECT 1613.8800 739.1400 1615.4800 739.6200 ;
        RECT 1613.8800 744.5800 1615.4800 745.0600 ;
        RECT 1613.8800 750.0200 1615.4800 750.5000 ;
        RECT 1613.8800 728.2600 1615.4800 728.7400 ;
        RECT 1613.8800 733.7000 1615.4800 734.1800 ;
        RECT 1568.8800 739.1400 1570.4800 739.6200 ;
        RECT 1568.8800 744.5800 1570.4800 745.0600 ;
        RECT 1568.8800 750.0200 1570.4800 750.5000 ;
        RECT 1568.8800 728.2600 1570.4800 728.7400 ;
        RECT 1568.8800 733.7000 1570.4800 734.1800 ;
        RECT 1613.8800 711.9400 1615.4800 712.4200 ;
        RECT 1613.8800 717.3800 1615.4800 717.8600 ;
        RECT 1613.8800 722.8200 1615.4800 723.3000 ;
        RECT 1613.8800 701.0600 1615.4800 701.5400 ;
        RECT 1613.8800 706.5000 1615.4800 706.9800 ;
        RECT 1568.8800 711.9400 1570.4800 712.4200 ;
        RECT 1568.8800 717.3800 1570.4800 717.8600 ;
        RECT 1568.8800 722.8200 1570.4800 723.3000 ;
        RECT 1568.8800 701.0600 1570.4800 701.5400 ;
        RECT 1568.8800 706.5000 1570.4800 706.9800 ;
        RECT 1523.8800 739.1400 1525.4800 739.6200 ;
        RECT 1523.8800 744.5800 1525.4800 745.0600 ;
        RECT 1523.8800 750.0200 1525.4800 750.5000 ;
        RECT 1516.1200 739.1400 1517.7200 739.6200 ;
        RECT 1516.1200 744.5800 1517.7200 745.0600 ;
        RECT 1516.1200 750.0200 1517.7200 750.5000 ;
        RECT 1523.8800 728.2600 1525.4800 728.7400 ;
        RECT 1523.8800 733.7000 1525.4800 734.1800 ;
        RECT 1516.1200 728.2600 1517.7200 728.7400 ;
        RECT 1516.1200 733.7000 1517.7200 734.1800 ;
        RECT 1523.8800 711.9400 1525.4800 712.4200 ;
        RECT 1523.8800 717.3800 1525.4800 717.8600 ;
        RECT 1523.8800 722.8200 1525.4800 723.3000 ;
        RECT 1516.1200 711.9400 1517.7200 712.4200 ;
        RECT 1516.1200 717.3800 1517.7200 717.8600 ;
        RECT 1516.1200 722.8200 1517.7200 723.3000 ;
        RECT 1523.8800 701.0600 1525.4800 701.5400 ;
        RECT 1523.8800 706.5000 1525.4800 706.9800 ;
        RECT 1516.1200 701.0600 1517.7200 701.5400 ;
        RECT 1516.1200 706.5000 1517.7200 706.9800 ;
        RECT 1613.8800 684.7400 1615.4800 685.2200 ;
        RECT 1613.8800 690.1800 1615.4800 690.6600 ;
        RECT 1613.8800 695.6200 1615.4800 696.1000 ;
        RECT 1613.8800 673.8600 1615.4800 674.3400 ;
        RECT 1613.8800 679.3000 1615.4800 679.7800 ;
        RECT 1568.8800 684.7400 1570.4800 685.2200 ;
        RECT 1568.8800 690.1800 1570.4800 690.6600 ;
        RECT 1568.8800 695.6200 1570.4800 696.1000 ;
        RECT 1568.8800 673.8600 1570.4800 674.3400 ;
        RECT 1568.8800 679.3000 1570.4800 679.7800 ;
        RECT 1613.8800 657.5400 1615.4800 658.0200 ;
        RECT 1613.8800 662.9800 1615.4800 663.4600 ;
        RECT 1613.8800 668.4200 1615.4800 668.9000 ;
        RECT 1613.8800 652.1000 1615.4800 652.5800 ;
        RECT 1568.8800 657.5400 1570.4800 658.0200 ;
        RECT 1568.8800 662.9800 1570.4800 663.4600 ;
        RECT 1568.8800 668.4200 1570.4800 668.9000 ;
        RECT 1568.8800 652.1000 1570.4800 652.5800 ;
        RECT 1523.8800 684.7400 1525.4800 685.2200 ;
        RECT 1523.8800 690.1800 1525.4800 690.6600 ;
        RECT 1523.8800 695.6200 1525.4800 696.1000 ;
        RECT 1516.1200 684.7400 1517.7200 685.2200 ;
        RECT 1516.1200 690.1800 1517.7200 690.6600 ;
        RECT 1516.1200 695.6200 1517.7200 696.1000 ;
        RECT 1523.8800 673.8600 1525.4800 674.3400 ;
        RECT 1523.8800 679.3000 1525.4800 679.7800 ;
        RECT 1516.1200 673.8600 1517.7200 674.3400 ;
        RECT 1516.1200 679.3000 1517.7200 679.7800 ;
        RECT 1523.8800 657.5400 1525.4800 658.0200 ;
        RECT 1523.8800 662.9800 1525.4800 663.4600 ;
        RECT 1523.8800 668.4200 1525.4800 668.9000 ;
        RECT 1516.1200 657.5400 1517.7200 658.0200 ;
        RECT 1516.1200 662.9800 1517.7200 663.4600 ;
        RECT 1516.1200 668.4200 1517.7200 668.9000 ;
        RECT 1516.1200 652.1000 1517.7200 652.5800 ;
        RECT 1523.8800 652.1000 1525.4800 652.5800 ;
        RECT 1510.5600 854.4100 1720.7800 856.0100 ;
        RECT 1510.5600 647.9100 1720.7800 649.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 642.4800 1517.7200 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 860.5200 1517.7200 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 642.4800 1715.2200 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 860.5200 1715.2200 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 647.9100 1512.1600 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 647.9100 1720.7800 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 854.4100 1512.1600 856.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 854.4100 1720.7800 856.0100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1703.8800 418.2700 1705.4800 626.3700 ;
        RECT 1658.8800 418.2700 1660.4800 626.3700 ;
        RECT 1613.8800 418.2700 1615.4800 626.3700 ;
        RECT 1568.8800 418.2700 1570.4800 626.3700 ;
        RECT 1523.8800 418.2700 1525.4800 626.3700 ;
        RECT 1713.6200 412.8400 1715.2200 632.4800 ;
        RECT 1516.1200 412.8400 1517.7200 632.4800 ;
      LAYER met3 ;
        RECT 1713.6200 607.4200 1715.2200 607.9000 ;
        RECT 1713.6200 612.8600 1715.2200 613.3400 ;
        RECT 1703.8800 607.4200 1705.4800 607.9000 ;
        RECT 1703.8800 612.8600 1705.4800 613.3400 ;
        RECT 1703.8800 618.3000 1705.4800 618.7800 ;
        RECT 1713.6200 618.3000 1715.2200 618.7800 ;
        RECT 1713.6200 596.5400 1715.2200 597.0200 ;
        RECT 1713.6200 601.9800 1715.2200 602.4600 ;
        RECT 1703.8800 596.5400 1705.4800 597.0200 ;
        RECT 1703.8800 601.9800 1705.4800 602.4600 ;
        RECT 1713.6200 580.2200 1715.2200 580.7000 ;
        RECT 1713.6200 585.6600 1715.2200 586.1400 ;
        RECT 1703.8800 580.2200 1705.4800 580.7000 ;
        RECT 1703.8800 585.6600 1705.4800 586.1400 ;
        RECT 1703.8800 591.1000 1705.4800 591.5800 ;
        RECT 1713.6200 591.1000 1715.2200 591.5800 ;
        RECT 1658.8800 607.4200 1660.4800 607.9000 ;
        RECT 1658.8800 612.8600 1660.4800 613.3400 ;
        RECT 1658.8800 618.3000 1660.4800 618.7800 ;
        RECT 1658.8800 596.5400 1660.4800 597.0200 ;
        RECT 1658.8800 601.9800 1660.4800 602.4600 ;
        RECT 1658.8800 580.2200 1660.4800 580.7000 ;
        RECT 1658.8800 585.6600 1660.4800 586.1400 ;
        RECT 1658.8800 591.1000 1660.4800 591.5800 ;
        RECT 1713.6200 563.9000 1715.2200 564.3800 ;
        RECT 1713.6200 569.3400 1715.2200 569.8200 ;
        RECT 1713.6200 574.7800 1715.2200 575.2600 ;
        RECT 1703.8800 563.9000 1705.4800 564.3800 ;
        RECT 1703.8800 569.3400 1705.4800 569.8200 ;
        RECT 1703.8800 574.7800 1705.4800 575.2600 ;
        RECT 1713.6200 553.0200 1715.2200 553.5000 ;
        RECT 1713.6200 558.4600 1715.2200 558.9400 ;
        RECT 1703.8800 553.0200 1705.4800 553.5000 ;
        RECT 1703.8800 558.4600 1705.4800 558.9400 ;
        RECT 1713.6200 536.7000 1715.2200 537.1800 ;
        RECT 1713.6200 542.1400 1715.2200 542.6200 ;
        RECT 1713.6200 547.5800 1715.2200 548.0600 ;
        RECT 1703.8800 536.7000 1705.4800 537.1800 ;
        RECT 1703.8800 542.1400 1705.4800 542.6200 ;
        RECT 1703.8800 547.5800 1705.4800 548.0600 ;
        RECT 1713.6200 525.8200 1715.2200 526.3000 ;
        RECT 1713.6200 531.2600 1715.2200 531.7400 ;
        RECT 1703.8800 525.8200 1705.4800 526.3000 ;
        RECT 1703.8800 531.2600 1705.4800 531.7400 ;
        RECT 1658.8800 563.9000 1660.4800 564.3800 ;
        RECT 1658.8800 569.3400 1660.4800 569.8200 ;
        RECT 1658.8800 574.7800 1660.4800 575.2600 ;
        RECT 1658.8800 553.0200 1660.4800 553.5000 ;
        RECT 1658.8800 558.4600 1660.4800 558.9400 ;
        RECT 1658.8800 536.7000 1660.4800 537.1800 ;
        RECT 1658.8800 542.1400 1660.4800 542.6200 ;
        RECT 1658.8800 547.5800 1660.4800 548.0600 ;
        RECT 1658.8800 525.8200 1660.4800 526.3000 ;
        RECT 1658.8800 531.2600 1660.4800 531.7400 ;
        RECT 1613.8800 607.4200 1615.4800 607.9000 ;
        RECT 1613.8800 612.8600 1615.4800 613.3400 ;
        RECT 1613.8800 618.3000 1615.4800 618.7800 ;
        RECT 1568.8800 607.4200 1570.4800 607.9000 ;
        RECT 1568.8800 612.8600 1570.4800 613.3400 ;
        RECT 1568.8800 618.3000 1570.4800 618.7800 ;
        RECT 1613.8800 596.5400 1615.4800 597.0200 ;
        RECT 1613.8800 601.9800 1615.4800 602.4600 ;
        RECT 1613.8800 580.2200 1615.4800 580.7000 ;
        RECT 1613.8800 585.6600 1615.4800 586.1400 ;
        RECT 1613.8800 591.1000 1615.4800 591.5800 ;
        RECT 1568.8800 596.5400 1570.4800 597.0200 ;
        RECT 1568.8800 601.9800 1570.4800 602.4600 ;
        RECT 1568.8800 580.2200 1570.4800 580.7000 ;
        RECT 1568.8800 585.6600 1570.4800 586.1400 ;
        RECT 1568.8800 591.1000 1570.4800 591.5800 ;
        RECT 1523.8800 607.4200 1525.4800 607.9000 ;
        RECT 1523.8800 612.8600 1525.4800 613.3400 ;
        RECT 1516.1200 607.4200 1517.7200 607.9000 ;
        RECT 1516.1200 612.8600 1517.7200 613.3400 ;
        RECT 1516.1200 618.3000 1517.7200 618.7800 ;
        RECT 1523.8800 618.3000 1525.4800 618.7800 ;
        RECT 1523.8800 596.5400 1525.4800 597.0200 ;
        RECT 1523.8800 601.9800 1525.4800 602.4600 ;
        RECT 1516.1200 596.5400 1517.7200 597.0200 ;
        RECT 1516.1200 601.9800 1517.7200 602.4600 ;
        RECT 1523.8800 580.2200 1525.4800 580.7000 ;
        RECT 1523.8800 585.6600 1525.4800 586.1400 ;
        RECT 1516.1200 580.2200 1517.7200 580.7000 ;
        RECT 1516.1200 585.6600 1517.7200 586.1400 ;
        RECT 1516.1200 591.1000 1517.7200 591.5800 ;
        RECT 1523.8800 591.1000 1525.4800 591.5800 ;
        RECT 1613.8800 563.9000 1615.4800 564.3800 ;
        RECT 1613.8800 569.3400 1615.4800 569.8200 ;
        RECT 1613.8800 574.7800 1615.4800 575.2600 ;
        RECT 1613.8800 553.0200 1615.4800 553.5000 ;
        RECT 1613.8800 558.4600 1615.4800 558.9400 ;
        RECT 1568.8800 563.9000 1570.4800 564.3800 ;
        RECT 1568.8800 569.3400 1570.4800 569.8200 ;
        RECT 1568.8800 574.7800 1570.4800 575.2600 ;
        RECT 1568.8800 553.0200 1570.4800 553.5000 ;
        RECT 1568.8800 558.4600 1570.4800 558.9400 ;
        RECT 1613.8800 536.7000 1615.4800 537.1800 ;
        RECT 1613.8800 542.1400 1615.4800 542.6200 ;
        RECT 1613.8800 547.5800 1615.4800 548.0600 ;
        RECT 1613.8800 525.8200 1615.4800 526.3000 ;
        RECT 1613.8800 531.2600 1615.4800 531.7400 ;
        RECT 1568.8800 536.7000 1570.4800 537.1800 ;
        RECT 1568.8800 542.1400 1570.4800 542.6200 ;
        RECT 1568.8800 547.5800 1570.4800 548.0600 ;
        RECT 1568.8800 525.8200 1570.4800 526.3000 ;
        RECT 1568.8800 531.2600 1570.4800 531.7400 ;
        RECT 1523.8800 563.9000 1525.4800 564.3800 ;
        RECT 1523.8800 569.3400 1525.4800 569.8200 ;
        RECT 1523.8800 574.7800 1525.4800 575.2600 ;
        RECT 1516.1200 563.9000 1517.7200 564.3800 ;
        RECT 1516.1200 569.3400 1517.7200 569.8200 ;
        RECT 1516.1200 574.7800 1517.7200 575.2600 ;
        RECT 1523.8800 553.0200 1525.4800 553.5000 ;
        RECT 1523.8800 558.4600 1525.4800 558.9400 ;
        RECT 1516.1200 553.0200 1517.7200 553.5000 ;
        RECT 1516.1200 558.4600 1517.7200 558.9400 ;
        RECT 1523.8800 536.7000 1525.4800 537.1800 ;
        RECT 1523.8800 542.1400 1525.4800 542.6200 ;
        RECT 1523.8800 547.5800 1525.4800 548.0600 ;
        RECT 1516.1200 536.7000 1517.7200 537.1800 ;
        RECT 1516.1200 542.1400 1517.7200 542.6200 ;
        RECT 1516.1200 547.5800 1517.7200 548.0600 ;
        RECT 1523.8800 525.8200 1525.4800 526.3000 ;
        RECT 1523.8800 531.2600 1525.4800 531.7400 ;
        RECT 1516.1200 525.8200 1517.7200 526.3000 ;
        RECT 1516.1200 531.2600 1517.7200 531.7400 ;
        RECT 1713.6200 509.5000 1715.2200 509.9800 ;
        RECT 1713.6200 514.9400 1715.2200 515.4200 ;
        RECT 1713.6200 520.3800 1715.2200 520.8600 ;
        RECT 1703.8800 509.5000 1705.4800 509.9800 ;
        RECT 1703.8800 514.9400 1705.4800 515.4200 ;
        RECT 1703.8800 520.3800 1705.4800 520.8600 ;
        RECT 1713.6200 498.6200 1715.2200 499.1000 ;
        RECT 1713.6200 504.0600 1715.2200 504.5400 ;
        RECT 1703.8800 498.6200 1705.4800 499.1000 ;
        RECT 1703.8800 504.0600 1705.4800 504.5400 ;
        RECT 1713.6200 482.3000 1715.2200 482.7800 ;
        RECT 1713.6200 487.7400 1715.2200 488.2200 ;
        RECT 1713.6200 493.1800 1715.2200 493.6600 ;
        RECT 1703.8800 482.3000 1705.4800 482.7800 ;
        RECT 1703.8800 487.7400 1705.4800 488.2200 ;
        RECT 1703.8800 493.1800 1705.4800 493.6600 ;
        RECT 1713.6200 471.4200 1715.2200 471.9000 ;
        RECT 1713.6200 476.8600 1715.2200 477.3400 ;
        RECT 1703.8800 471.4200 1705.4800 471.9000 ;
        RECT 1703.8800 476.8600 1705.4800 477.3400 ;
        RECT 1658.8800 509.5000 1660.4800 509.9800 ;
        RECT 1658.8800 514.9400 1660.4800 515.4200 ;
        RECT 1658.8800 520.3800 1660.4800 520.8600 ;
        RECT 1658.8800 498.6200 1660.4800 499.1000 ;
        RECT 1658.8800 504.0600 1660.4800 504.5400 ;
        RECT 1658.8800 482.3000 1660.4800 482.7800 ;
        RECT 1658.8800 487.7400 1660.4800 488.2200 ;
        RECT 1658.8800 493.1800 1660.4800 493.6600 ;
        RECT 1658.8800 471.4200 1660.4800 471.9000 ;
        RECT 1658.8800 476.8600 1660.4800 477.3400 ;
        RECT 1713.6200 455.1000 1715.2200 455.5800 ;
        RECT 1713.6200 460.5400 1715.2200 461.0200 ;
        RECT 1713.6200 465.9800 1715.2200 466.4600 ;
        RECT 1703.8800 455.1000 1705.4800 455.5800 ;
        RECT 1703.8800 460.5400 1705.4800 461.0200 ;
        RECT 1703.8800 465.9800 1705.4800 466.4600 ;
        RECT 1713.6200 444.2200 1715.2200 444.7000 ;
        RECT 1713.6200 449.6600 1715.2200 450.1400 ;
        RECT 1703.8800 444.2200 1705.4800 444.7000 ;
        RECT 1703.8800 449.6600 1705.4800 450.1400 ;
        RECT 1713.6200 427.9000 1715.2200 428.3800 ;
        RECT 1713.6200 433.3400 1715.2200 433.8200 ;
        RECT 1713.6200 438.7800 1715.2200 439.2600 ;
        RECT 1703.8800 427.9000 1705.4800 428.3800 ;
        RECT 1703.8800 433.3400 1705.4800 433.8200 ;
        RECT 1703.8800 438.7800 1705.4800 439.2600 ;
        RECT 1703.8800 422.4600 1705.4800 422.9400 ;
        RECT 1713.6200 422.4600 1715.2200 422.9400 ;
        RECT 1658.8800 455.1000 1660.4800 455.5800 ;
        RECT 1658.8800 460.5400 1660.4800 461.0200 ;
        RECT 1658.8800 465.9800 1660.4800 466.4600 ;
        RECT 1658.8800 444.2200 1660.4800 444.7000 ;
        RECT 1658.8800 449.6600 1660.4800 450.1400 ;
        RECT 1658.8800 427.9000 1660.4800 428.3800 ;
        RECT 1658.8800 433.3400 1660.4800 433.8200 ;
        RECT 1658.8800 438.7800 1660.4800 439.2600 ;
        RECT 1658.8800 422.4600 1660.4800 422.9400 ;
        RECT 1613.8800 509.5000 1615.4800 509.9800 ;
        RECT 1613.8800 514.9400 1615.4800 515.4200 ;
        RECT 1613.8800 520.3800 1615.4800 520.8600 ;
        RECT 1613.8800 498.6200 1615.4800 499.1000 ;
        RECT 1613.8800 504.0600 1615.4800 504.5400 ;
        RECT 1568.8800 509.5000 1570.4800 509.9800 ;
        RECT 1568.8800 514.9400 1570.4800 515.4200 ;
        RECT 1568.8800 520.3800 1570.4800 520.8600 ;
        RECT 1568.8800 498.6200 1570.4800 499.1000 ;
        RECT 1568.8800 504.0600 1570.4800 504.5400 ;
        RECT 1613.8800 482.3000 1615.4800 482.7800 ;
        RECT 1613.8800 487.7400 1615.4800 488.2200 ;
        RECT 1613.8800 493.1800 1615.4800 493.6600 ;
        RECT 1613.8800 471.4200 1615.4800 471.9000 ;
        RECT 1613.8800 476.8600 1615.4800 477.3400 ;
        RECT 1568.8800 482.3000 1570.4800 482.7800 ;
        RECT 1568.8800 487.7400 1570.4800 488.2200 ;
        RECT 1568.8800 493.1800 1570.4800 493.6600 ;
        RECT 1568.8800 471.4200 1570.4800 471.9000 ;
        RECT 1568.8800 476.8600 1570.4800 477.3400 ;
        RECT 1523.8800 509.5000 1525.4800 509.9800 ;
        RECT 1523.8800 514.9400 1525.4800 515.4200 ;
        RECT 1523.8800 520.3800 1525.4800 520.8600 ;
        RECT 1516.1200 509.5000 1517.7200 509.9800 ;
        RECT 1516.1200 514.9400 1517.7200 515.4200 ;
        RECT 1516.1200 520.3800 1517.7200 520.8600 ;
        RECT 1523.8800 498.6200 1525.4800 499.1000 ;
        RECT 1523.8800 504.0600 1525.4800 504.5400 ;
        RECT 1516.1200 498.6200 1517.7200 499.1000 ;
        RECT 1516.1200 504.0600 1517.7200 504.5400 ;
        RECT 1523.8800 482.3000 1525.4800 482.7800 ;
        RECT 1523.8800 487.7400 1525.4800 488.2200 ;
        RECT 1523.8800 493.1800 1525.4800 493.6600 ;
        RECT 1516.1200 482.3000 1517.7200 482.7800 ;
        RECT 1516.1200 487.7400 1517.7200 488.2200 ;
        RECT 1516.1200 493.1800 1517.7200 493.6600 ;
        RECT 1523.8800 471.4200 1525.4800 471.9000 ;
        RECT 1523.8800 476.8600 1525.4800 477.3400 ;
        RECT 1516.1200 471.4200 1517.7200 471.9000 ;
        RECT 1516.1200 476.8600 1517.7200 477.3400 ;
        RECT 1613.8800 455.1000 1615.4800 455.5800 ;
        RECT 1613.8800 460.5400 1615.4800 461.0200 ;
        RECT 1613.8800 465.9800 1615.4800 466.4600 ;
        RECT 1613.8800 444.2200 1615.4800 444.7000 ;
        RECT 1613.8800 449.6600 1615.4800 450.1400 ;
        RECT 1568.8800 455.1000 1570.4800 455.5800 ;
        RECT 1568.8800 460.5400 1570.4800 461.0200 ;
        RECT 1568.8800 465.9800 1570.4800 466.4600 ;
        RECT 1568.8800 444.2200 1570.4800 444.7000 ;
        RECT 1568.8800 449.6600 1570.4800 450.1400 ;
        RECT 1613.8800 427.9000 1615.4800 428.3800 ;
        RECT 1613.8800 433.3400 1615.4800 433.8200 ;
        RECT 1613.8800 438.7800 1615.4800 439.2600 ;
        RECT 1613.8800 422.4600 1615.4800 422.9400 ;
        RECT 1568.8800 427.9000 1570.4800 428.3800 ;
        RECT 1568.8800 433.3400 1570.4800 433.8200 ;
        RECT 1568.8800 438.7800 1570.4800 439.2600 ;
        RECT 1568.8800 422.4600 1570.4800 422.9400 ;
        RECT 1523.8800 455.1000 1525.4800 455.5800 ;
        RECT 1523.8800 460.5400 1525.4800 461.0200 ;
        RECT 1523.8800 465.9800 1525.4800 466.4600 ;
        RECT 1516.1200 455.1000 1517.7200 455.5800 ;
        RECT 1516.1200 460.5400 1517.7200 461.0200 ;
        RECT 1516.1200 465.9800 1517.7200 466.4600 ;
        RECT 1523.8800 444.2200 1525.4800 444.7000 ;
        RECT 1523.8800 449.6600 1525.4800 450.1400 ;
        RECT 1516.1200 444.2200 1517.7200 444.7000 ;
        RECT 1516.1200 449.6600 1517.7200 450.1400 ;
        RECT 1523.8800 427.9000 1525.4800 428.3800 ;
        RECT 1523.8800 433.3400 1525.4800 433.8200 ;
        RECT 1523.8800 438.7800 1525.4800 439.2600 ;
        RECT 1516.1200 427.9000 1517.7200 428.3800 ;
        RECT 1516.1200 433.3400 1517.7200 433.8200 ;
        RECT 1516.1200 438.7800 1517.7200 439.2600 ;
        RECT 1516.1200 422.4600 1517.7200 422.9400 ;
        RECT 1523.8800 422.4600 1525.4800 422.9400 ;
        RECT 1510.5600 624.7700 1720.7800 626.3700 ;
        RECT 1510.5600 418.2700 1720.7800 419.8700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 412.8400 1517.7200 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.1200 630.8800 1517.7200 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 412.8400 1715.2200 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1713.6200 630.8800 1715.2200 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 418.2700 1512.1600 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 418.2700 1720.7800 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1510.5600 624.7700 1512.1600 626.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1719.1800 624.7700 1720.7800 626.3700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 1736.2400 2479.6000 1737.8400 2509.8600 ;
        RECT 1933.9400 2479.6000 1935.5400 2509.8600 ;
      LAYER met3 ;
        RECT 1933.9400 2497.3800 1935.5400 2497.8600 ;
        RECT 1736.2400 2497.3800 1737.8400 2497.8600 ;
        RECT 1933.9400 2491.9400 1935.5400 2492.4200 ;
        RECT 1933.9400 2486.5000 1935.5400 2486.9800 ;
        RECT 1736.2400 2491.9400 1737.8400 2492.4200 ;
        RECT 1736.2400 2486.5000 1737.8400 2486.9800 ;
        RECT 1730.7800 2503.1000 1941.0000 2504.7000 ;
        RECT 1730.7800 2483.5700 1941.0000 2485.1700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.2400 2479.6000 1737.8400 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.2400 2508.2600 1737.8400 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.9400 2479.6000 1935.5400 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.9400 2508.2600 1935.5400 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2483.5700 1732.3800 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2483.5700 1941.0000 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2503.1000 1732.3800 2504.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2503.1000 1941.0000 2504.7000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 188.6300 1925.7000 396.7300 ;
        RECT 1879.1000 188.6300 1880.7000 396.7300 ;
        RECT 1834.1000 188.6300 1835.7000 396.7300 ;
        RECT 1789.1000 188.6300 1790.7000 396.7300 ;
        RECT 1744.1000 188.6300 1745.7000 396.7300 ;
        RECT 1933.8400 183.2000 1935.4400 402.8400 ;
        RECT 1736.3400 183.2000 1737.9400 402.8400 ;
      LAYER met3 ;
        RECT 1933.8400 377.7800 1935.4400 378.2600 ;
        RECT 1933.8400 383.2200 1935.4400 383.7000 ;
        RECT 1924.1000 377.7800 1925.7000 378.2600 ;
        RECT 1924.1000 383.2200 1925.7000 383.7000 ;
        RECT 1924.1000 388.6600 1925.7000 389.1400 ;
        RECT 1933.8400 388.6600 1935.4400 389.1400 ;
        RECT 1933.8400 366.9000 1935.4400 367.3800 ;
        RECT 1933.8400 372.3400 1935.4400 372.8200 ;
        RECT 1924.1000 366.9000 1925.7000 367.3800 ;
        RECT 1924.1000 372.3400 1925.7000 372.8200 ;
        RECT 1933.8400 350.5800 1935.4400 351.0600 ;
        RECT 1933.8400 356.0200 1935.4400 356.5000 ;
        RECT 1924.1000 350.5800 1925.7000 351.0600 ;
        RECT 1924.1000 356.0200 1925.7000 356.5000 ;
        RECT 1924.1000 361.4600 1925.7000 361.9400 ;
        RECT 1933.8400 361.4600 1935.4400 361.9400 ;
        RECT 1879.1000 377.7800 1880.7000 378.2600 ;
        RECT 1879.1000 383.2200 1880.7000 383.7000 ;
        RECT 1879.1000 388.6600 1880.7000 389.1400 ;
        RECT 1879.1000 366.9000 1880.7000 367.3800 ;
        RECT 1879.1000 372.3400 1880.7000 372.8200 ;
        RECT 1879.1000 350.5800 1880.7000 351.0600 ;
        RECT 1879.1000 356.0200 1880.7000 356.5000 ;
        RECT 1879.1000 361.4600 1880.7000 361.9400 ;
        RECT 1933.8400 334.2600 1935.4400 334.7400 ;
        RECT 1933.8400 339.7000 1935.4400 340.1800 ;
        RECT 1933.8400 345.1400 1935.4400 345.6200 ;
        RECT 1924.1000 334.2600 1925.7000 334.7400 ;
        RECT 1924.1000 339.7000 1925.7000 340.1800 ;
        RECT 1924.1000 345.1400 1925.7000 345.6200 ;
        RECT 1933.8400 323.3800 1935.4400 323.8600 ;
        RECT 1933.8400 328.8200 1935.4400 329.3000 ;
        RECT 1924.1000 323.3800 1925.7000 323.8600 ;
        RECT 1924.1000 328.8200 1925.7000 329.3000 ;
        RECT 1933.8400 307.0600 1935.4400 307.5400 ;
        RECT 1933.8400 312.5000 1935.4400 312.9800 ;
        RECT 1933.8400 317.9400 1935.4400 318.4200 ;
        RECT 1924.1000 307.0600 1925.7000 307.5400 ;
        RECT 1924.1000 312.5000 1925.7000 312.9800 ;
        RECT 1924.1000 317.9400 1925.7000 318.4200 ;
        RECT 1933.8400 296.1800 1935.4400 296.6600 ;
        RECT 1933.8400 301.6200 1935.4400 302.1000 ;
        RECT 1924.1000 296.1800 1925.7000 296.6600 ;
        RECT 1924.1000 301.6200 1925.7000 302.1000 ;
        RECT 1879.1000 334.2600 1880.7000 334.7400 ;
        RECT 1879.1000 339.7000 1880.7000 340.1800 ;
        RECT 1879.1000 345.1400 1880.7000 345.6200 ;
        RECT 1879.1000 323.3800 1880.7000 323.8600 ;
        RECT 1879.1000 328.8200 1880.7000 329.3000 ;
        RECT 1879.1000 307.0600 1880.7000 307.5400 ;
        RECT 1879.1000 312.5000 1880.7000 312.9800 ;
        RECT 1879.1000 317.9400 1880.7000 318.4200 ;
        RECT 1879.1000 296.1800 1880.7000 296.6600 ;
        RECT 1879.1000 301.6200 1880.7000 302.1000 ;
        RECT 1834.1000 377.7800 1835.7000 378.2600 ;
        RECT 1834.1000 383.2200 1835.7000 383.7000 ;
        RECT 1834.1000 388.6600 1835.7000 389.1400 ;
        RECT 1789.1000 377.7800 1790.7000 378.2600 ;
        RECT 1789.1000 383.2200 1790.7000 383.7000 ;
        RECT 1789.1000 388.6600 1790.7000 389.1400 ;
        RECT 1834.1000 366.9000 1835.7000 367.3800 ;
        RECT 1834.1000 372.3400 1835.7000 372.8200 ;
        RECT 1834.1000 350.5800 1835.7000 351.0600 ;
        RECT 1834.1000 356.0200 1835.7000 356.5000 ;
        RECT 1834.1000 361.4600 1835.7000 361.9400 ;
        RECT 1789.1000 366.9000 1790.7000 367.3800 ;
        RECT 1789.1000 372.3400 1790.7000 372.8200 ;
        RECT 1789.1000 350.5800 1790.7000 351.0600 ;
        RECT 1789.1000 356.0200 1790.7000 356.5000 ;
        RECT 1789.1000 361.4600 1790.7000 361.9400 ;
        RECT 1744.1000 377.7800 1745.7000 378.2600 ;
        RECT 1744.1000 383.2200 1745.7000 383.7000 ;
        RECT 1736.3400 377.7800 1737.9400 378.2600 ;
        RECT 1736.3400 383.2200 1737.9400 383.7000 ;
        RECT 1736.3400 388.6600 1737.9400 389.1400 ;
        RECT 1744.1000 388.6600 1745.7000 389.1400 ;
        RECT 1744.1000 366.9000 1745.7000 367.3800 ;
        RECT 1744.1000 372.3400 1745.7000 372.8200 ;
        RECT 1736.3400 366.9000 1737.9400 367.3800 ;
        RECT 1736.3400 372.3400 1737.9400 372.8200 ;
        RECT 1744.1000 350.5800 1745.7000 351.0600 ;
        RECT 1744.1000 356.0200 1745.7000 356.5000 ;
        RECT 1736.3400 350.5800 1737.9400 351.0600 ;
        RECT 1736.3400 356.0200 1737.9400 356.5000 ;
        RECT 1736.3400 361.4600 1737.9400 361.9400 ;
        RECT 1744.1000 361.4600 1745.7000 361.9400 ;
        RECT 1834.1000 334.2600 1835.7000 334.7400 ;
        RECT 1834.1000 339.7000 1835.7000 340.1800 ;
        RECT 1834.1000 345.1400 1835.7000 345.6200 ;
        RECT 1834.1000 323.3800 1835.7000 323.8600 ;
        RECT 1834.1000 328.8200 1835.7000 329.3000 ;
        RECT 1789.1000 334.2600 1790.7000 334.7400 ;
        RECT 1789.1000 339.7000 1790.7000 340.1800 ;
        RECT 1789.1000 345.1400 1790.7000 345.6200 ;
        RECT 1789.1000 323.3800 1790.7000 323.8600 ;
        RECT 1789.1000 328.8200 1790.7000 329.3000 ;
        RECT 1834.1000 307.0600 1835.7000 307.5400 ;
        RECT 1834.1000 312.5000 1835.7000 312.9800 ;
        RECT 1834.1000 317.9400 1835.7000 318.4200 ;
        RECT 1834.1000 296.1800 1835.7000 296.6600 ;
        RECT 1834.1000 301.6200 1835.7000 302.1000 ;
        RECT 1789.1000 307.0600 1790.7000 307.5400 ;
        RECT 1789.1000 312.5000 1790.7000 312.9800 ;
        RECT 1789.1000 317.9400 1790.7000 318.4200 ;
        RECT 1789.1000 296.1800 1790.7000 296.6600 ;
        RECT 1789.1000 301.6200 1790.7000 302.1000 ;
        RECT 1744.1000 334.2600 1745.7000 334.7400 ;
        RECT 1744.1000 339.7000 1745.7000 340.1800 ;
        RECT 1744.1000 345.1400 1745.7000 345.6200 ;
        RECT 1736.3400 334.2600 1737.9400 334.7400 ;
        RECT 1736.3400 339.7000 1737.9400 340.1800 ;
        RECT 1736.3400 345.1400 1737.9400 345.6200 ;
        RECT 1744.1000 323.3800 1745.7000 323.8600 ;
        RECT 1744.1000 328.8200 1745.7000 329.3000 ;
        RECT 1736.3400 323.3800 1737.9400 323.8600 ;
        RECT 1736.3400 328.8200 1737.9400 329.3000 ;
        RECT 1744.1000 307.0600 1745.7000 307.5400 ;
        RECT 1744.1000 312.5000 1745.7000 312.9800 ;
        RECT 1744.1000 317.9400 1745.7000 318.4200 ;
        RECT 1736.3400 307.0600 1737.9400 307.5400 ;
        RECT 1736.3400 312.5000 1737.9400 312.9800 ;
        RECT 1736.3400 317.9400 1737.9400 318.4200 ;
        RECT 1744.1000 296.1800 1745.7000 296.6600 ;
        RECT 1744.1000 301.6200 1745.7000 302.1000 ;
        RECT 1736.3400 296.1800 1737.9400 296.6600 ;
        RECT 1736.3400 301.6200 1737.9400 302.1000 ;
        RECT 1933.8400 279.8600 1935.4400 280.3400 ;
        RECT 1933.8400 285.3000 1935.4400 285.7800 ;
        RECT 1933.8400 290.7400 1935.4400 291.2200 ;
        RECT 1924.1000 279.8600 1925.7000 280.3400 ;
        RECT 1924.1000 285.3000 1925.7000 285.7800 ;
        RECT 1924.1000 290.7400 1925.7000 291.2200 ;
        RECT 1933.8400 268.9800 1935.4400 269.4600 ;
        RECT 1933.8400 274.4200 1935.4400 274.9000 ;
        RECT 1924.1000 268.9800 1925.7000 269.4600 ;
        RECT 1924.1000 274.4200 1925.7000 274.9000 ;
        RECT 1933.8400 252.6600 1935.4400 253.1400 ;
        RECT 1933.8400 258.1000 1935.4400 258.5800 ;
        RECT 1933.8400 263.5400 1935.4400 264.0200 ;
        RECT 1924.1000 252.6600 1925.7000 253.1400 ;
        RECT 1924.1000 258.1000 1925.7000 258.5800 ;
        RECT 1924.1000 263.5400 1925.7000 264.0200 ;
        RECT 1933.8400 241.7800 1935.4400 242.2600 ;
        RECT 1933.8400 247.2200 1935.4400 247.7000 ;
        RECT 1924.1000 241.7800 1925.7000 242.2600 ;
        RECT 1924.1000 247.2200 1925.7000 247.7000 ;
        RECT 1879.1000 279.8600 1880.7000 280.3400 ;
        RECT 1879.1000 285.3000 1880.7000 285.7800 ;
        RECT 1879.1000 290.7400 1880.7000 291.2200 ;
        RECT 1879.1000 268.9800 1880.7000 269.4600 ;
        RECT 1879.1000 274.4200 1880.7000 274.9000 ;
        RECT 1879.1000 252.6600 1880.7000 253.1400 ;
        RECT 1879.1000 258.1000 1880.7000 258.5800 ;
        RECT 1879.1000 263.5400 1880.7000 264.0200 ;
        RECT 1879.1000 241.7800 1880.7000 242.2600 ;
        RECT 1879.1000 247.2200 1880.7000 247.7000 ;
        RECT 1933.8400 225.4600 1935.4400 225.9400 ;
        RECT 1933.8400 230.9000 1935.4400 231.3800 ;
        RECT 1933.8400 236.3400 1935.4400 236.8200 ;
        RECT 1924.1000 225.4600 1925.7000 225.9400 ;
        RECT 1924.1000 230.9000 1925.7000 231.3800 ;
        RECT 1924.1000 236.3400 1925.7000 236.8200 ;
        RECT 1933.8400 214.5800 1935.4400 215.0600 ;
        RECT 1933.8400 220.0200 1935.4400 220.5000 ;
        RECT 1924.1000 214.5800 1925.7000 215.0600 ;
        RECT 1924.1000 220.0200 1925.7000 220.5000 ;
        RECT 1933.8400 198.2600 1935.4400 198.7400 ;
        RECT 1933.8400 203.7000 1935.4400 204.1800 ;
        RECT 1933.8400 209.1400 1935.4400 209.6200 ;
        RECT 1924.1000 198.2600 1925.7000 198.7400 ;
        RECT 1924.1000 203.7000 1925.7000 204.1800 ;
        RECT 1924.1000 209.1400 1925.7000 209.6200 ;
        RECT 1924.1000 192.8200 1925.7000 193.3000 ;
        RECT 1933.8400 192.8200 1935.4400 193.3000 ;
        RECT 1879.1000 225.4600 1880.7000 225.9400 ;
        RECT 1879.1000 230.9000 1880.7000 231.3800 ;
        RECT 1879.1000 236.3400 1880.7000 236.8200 ;
        RECT 1879.1000 214.5800 1880.7000 215.0600 ;
        RECT 1879.1000 220.0200 1880.7000 220.5000 ;
        RECT 1879.1000 198.2600 1880.7000 198.7400 ;
        RECT 1879.1000 203.7000 1880.7000 204.1800 ;
        RECT 1879.1000 209.1400 1880.7000 209.6200 ;
        RECT 1879.1000 192.8200 1880.7000 193.3000 ;
        RECT 1834.1000 279.8600 1835.7000 280.3400 ;
        RECT 1834.1000 285.3000 1835.7000 285.7800 ;
        RECT 1834.1000 290.7400 1835.7000 291.2200 ;
        RECT 1834.1000 268.9800 1835.7000 269.4600 ;
        RECT 1834.1000 274.4200 1835.7000 274.9000 ;
        RECT 1789.1000 279.8600 1790.7000 280.3400 ;
        RECT 1789.1000 285.3000 1790.7000 285.7800 ;
        RECT 1789.1000 290.7400 1790.7000 291.2200 ;
        RECT 1789.1000 268.9800 1790.7000 269.4600 ;
        RECT 1789.1000 274.4200 1790.7000 274.9000 ;
        RECT 1834.1000 252.6600 1835.7000 253.1400 ;
        RECT 1834.1000 258.1000 1835.7000 258.5800 ;
        RECT 1834.1000 263.5400 1835.7000 264.0200 ;
        RECT 1834.1000 241.7800 1835.7000 242.2600 ;
        RECT 1834.1000 247.2200 1835.7000 247.7000 ;
        RECT 1789.1000 252.6600 1790.7000 253.1400 ;
        RECT 1789.1000 258.1000 1790.7000 258.5800 ;
        RECT 1789.1000 263.5400 1790.7000 264.0200 ;
        RECT 1789.1000 241.7800 1790.7000 242.2600 ;
        RECT 1789.1000 247.2200 1790.7000 247.7000 ;
        RECT 1744.1000 279.8600 1745.7000 280.3400 ;
        RECT 1744.1000 285.3000 1745.7000 285.7800 ;
        RECT 1744.1000 290.7400 1745.7000 291.2200 ;
        RECT 1736.3400 279.8600 1737.9400 280.3400 ;
        RECT 1736.3400 285.3000 1737.9400 285.7800 ;
        RECT 1736.3400 290.7400 1737.9400 291.2200 ;
        RECT 1744.1000 268.9800 1745.7000 269.4600 ;
        RECT 1744.1000 274.4200 1745.7000 274.9000 ;
        RECT 1736.3400 268.9800 1737.9400 269.4600 ;
        RECT 1736.3400 274.4200 1737.9400 274.9000 ;
        RECT 1744.1000 252.6600 1745.7000 253.1400 ;
        RECT 1744.1000 258.1000 1745.7000 258.5800 ;
        RECT 1744.1000 263.5400 1745.7000 264.0200 ;
        RECT 1736.3400 252.6600 1737.9400 253.1400 ;
        RECT 1736.3400 258.1000 1737.9400 258.5800 ;
        RECT 1736.3400 263.5400 1737.9400 264.0200 ;
        RECT 1744.1000 241.7800 1745.7000 242.2600 ;
        RECT 1744.1000 247.2200 1745.7000 247.7000 ;
        RECT 1736.3400 241.7800 1737.9400 242.2600 ;
        RECT 1736.3400 247.2200 1737.9400 247.7000 ;
        RECT 1834.1000 225.4600 1835.7000 225.9400 ;
        RECT 1834.1000 230.9000 1835.7000 231.3800 ;
        RECT 1834.1000 236.3400 1835.7000 236.8200 ;
        RECT 1834.1000 214.5800 1835.7000 215.0600 ;
        RECT 1834.1000 220.0200 1835.7000 220.5000 ;
        RECT 1789.1000 225.4600 1790.7000 225.9400 ;
        RECT 1789.1000 230.9000 1790.7000 231.3800 ;
        RECT 1789.1000 236.3400 1790.7000 236.8200 ;
        RECT 1789.1000 214.5800 1790.7000 215.0600 ;
        RECT 1789.1000 220.0200 1790.7000 220.5000 ;
        RECT 1834.1000 198.2600 1835.7000 198.7400 ;
        RECT 1834.1000 203.7000 1835.7000 204.1800 ;
        RECT 1834.1000 209.1400 1835.7000 209.6200 ;
        RECT 1834.1000 192.8200 1835.7000 193.3000 ;
        RECT 1789.1000 198.2600 1790.7000 198.7400 ;
        RECT 1789.1000 203.7000 1790.7000 204.1800 ;
        RECT 1789.1000 209.1400 1790.7000 209.6200 ;
        RECT 1789.1000 192.8200 1790.7000 193.3000 ;
        RECT 1744.1000 225.4600 1745.7000 225.9400 ;
        RECT 1744.1000 230.9000 1745.7000 231.3800 ;
        RECT 1744.1000 236.3400 1745.7000 236.8200 ;
        RECT 1736.3400 225.4600 1737.9400 225.9400 ;
        RECT 1736.3400 230.9000 1737.9400 231.3800 ;
        RECT 1736.3400 236.3400 1737.9400 236.8200 ;
        RECT 1744.1000 214.5800 1745.7000 215.0600 ;
        RECT 1744.1000 220.0200 1745.7000 220.5000 ;
        RECT 1736.3400 214.5800 1737.9400 215.0600 ;
        RECT 1736.3400 220.0200 1737.9400 220.5000 ;
        RECT 1744.1000 198.2600 1745.7000 198.7400 ;
        RECT 1744.1000 203.7000 1745.7000 204.1800 ;
        RECT 1744.1000 209.1400 1745.7000 209.6200 ;
        RECT 1736.3400 198.2600 1737.9400 198.7400 ;
        RECT 1736.3400 203.7000 1737.9400 204.1800 ;
        RECT 1736.3400 209.1400 1737.9400 209.6200 ;
        RECT 1736.3400 192.8200 1737.9400 193.3000 ;
        RECT 1744.1000 192.8200 1745.7000 193.3000 ;
        RECT 1730.7800 395.1300 1941.0000 396.7300 ;
        RECT 1730.7800 188.6300 1941.0000 190.2300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 183.2000 1737.9400 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 401.2400 1737.9400 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 183.2000 1935.4400 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 401.2400 1935.4400 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 188.6300 1732.3800 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 188.6300 1941.0000 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 395.1300 1732.3800 396.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 395.1300 1941.0000 396.7300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 1736.2400 142.9400 1737.8400 173.2000 ;
        RECT 1933.9400 142.9400 1935.5400 173.2000 ;
      LAYER met3 ;
        RECT 1933.9400 160.7200 1935.5400 161.2000 ;
        RECT 1736.2400 160.7200 1737.8400 161.2000 ;
        RECT 1933.9400 155.2800 1935.5400 155.7600 ;
        RECT 1933.9400 149.8400 1935.5400 150.3200 ;
        RECT 1736.2400 155.2800 1737.8400 155.7600 ;
        RECT 1736.2400 149.8400 1737.8400 150.3200 ;
        RECT 1730.7800 166.4400 1941.0000 168.0400 ;
        RECT 1730.7800 146.9100 1941.0000 148.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.2400 142.9400 1737.8400 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.2400 171.6000 1737.8400 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.9400 142.9400 1935.5400 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.9400 171.6000 1935.5400 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 146.9100 1732.3800 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 146.9100 1941.0000 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 166.4400 1732.3800 168.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 166.4400 1941.0000 168.0400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 2255.3900 1925.7000 2463.4900 ;
        RECT 1879.1000 2255.3900 1880.7000 2463.4900 ;
        RECT 1834.1000 2255.3900 1835.7000 2463.4900 ;
        RECT 1789.1000 2255.3900 1790.7000 2463.4900 ;
        RECT 1744.1000 2255.3900 1745.7000 2463.4900 ;
        RECT 1933.8400 2249.9600 1935.4400 2469.6000 ;
        RECT 1736.3400 2249.9600 1737.9400 2469.6000 ;
      LAYER met3 ;
        RECT 1933.8400 2444.5400 1935.4400 2445.0200 ;
        RECT 1933.8400 2449.9800 1935.4400 2450.4600 ;
        RECT 1924.1000 2444.5400 1925.7000 2445.0200 ;
        RECT 1924.1000 2449.9800 1925.7000 2450.4600 ;
        RECT 1924.1000 2455.4200 1925.7000 2455.9000 ;
        RECT 1933.8400 2455.4200 1935.4400 2455.9000 ;
        RECT 1933.8400 2433.6600 1935.4400 2434.1400 ;
        RECT 1933.8400 2439.1000 1935.4400 2439.5800 ;
        RECT 1924.1000 2433.6600 1925.7000 2434.1400 ;
        RECT 1924.1000 2439.1000 1925.7000 2439.5800 ;
        RECT 1933.8400 2417.3400 1935.4400 2417.8200 ;
        RECT 1933.8400 2422.7800 1935.4400 2423.2600 ;
        RECT 1924.1000 2417.3400 1925.7000 2417.8200 ;
        RECT 1924.1000 2422.7800 1925.7000 2423.2600 ;
        RECT 1924.1000 2428.2200 1925.7000 2428.7000 ;
        RECT 1933.8400 2428.2200 1935.4400 2428.7000 ;
        RECT 1879.1000 2444.5400 1880.7000 2445.0200 ;
        RECT 1879.1000 2449.9800 1880.7000 2450.4600 ;
        RECT 1879.1000 2455.4200 1880.7000 2455.9000 ;
        RECT 1879.1000 2433.6600 1880.7000 2434.1400 ;
        RECT 1879.1000 2439.1000 1880.7000 2439.5800 ;
        RECT 1879.1000 2417.3400 1880.7000 2417.8200 ;
        RECT 1879.1000 2422.7800 1880.7000 2423.2600 ;
        RECT 1879.1000 2428.2200 1880.7000 2428.7000 ;
        RECT 1933.8400 2401.0200 1935.4400 2401.5000 ;
        RECT 1933.8400 2406.4600 1935.4400 2406.9400 ;
        RECT 1933.8400 2411.9000 1935.4400 2412.3800 ;
        RECT 1924.1000 2401.0200 1925.7000 2401.5000 ;
        RECT 1924.1000 2406.4600 1925.7000 2406.9400 ;
        RECT 1924.1000 2411.9000 1925.7000 2412.3800 ;
        RECT 1933.8400 2390.1400 1935.4400 2390.6200 ;
        RECT 1933.8400 2395.5800 1935.4400 2396.0600 ;
        RECT 1924.1000 2390.1400 1925.7000 2390.6200 ;
        RECT 1924.1000 2395.5800 1925.7000 2396.0600 ;
        RECT 1933.8400 2373.8200 1935.4400 2374.3000 ;
        RECT 1933.8400 2379.2600 1935.4400 2379.7400 ;
        RECT 1933.8400 2384.7000 1935.4400 2385.1800 ;
        RECT 1924.1000 2373.8200 1925.7000 2374.3000 ;
        RECT 1924.1000 2379.2600 1925.7000 2379.7400 ;
        RECT 1924.1000 2384.7000 1925.7000 2385.1800 ;
        RECT 1933.8400 2362.9400 1935.4400 2363.4200 ;
        RECT 1933.8400 2368.3800 1935.4400 2368.8600 ;
        RECT 1924.1000 2362.9400 1925.7000 2363.4200 ;
        RECT 1924.1000 2368.3800 1925.7000 2368.8600 ;
        RECT 1879.1000 2401.0200 1880.7000 2401.5000 ;
        RECT 1879.1000 2406.4600 1880.7000 2406.9400 ;
        RECT 1879.1000 2411.9000 1880.7000 2412.3800 ;
        RECT 1879.1000 2390.1400 1880.7000 2390.6200 ;
        RECT 1879.1000 2395.5800 1880.7000 2396.0600 ;
        RECT 1879.1000 2373.8200 1880.7000 2374.3000 ;
        RECT 1879.1000 2379.2600 1880.7000 2379.7400 ;
        RECT 1879.1000 2384.7000 1880.7000 2385.1800 ;
        RECT 1879.1000 2362.9400 1880.7000 2363.4200 ;
        RECT 1879.1000 2368.3800 1880.7000 2368.8600 ;
        RECT 1834.1000 2444.5400 1835.7000 2445.0200 ;
        RECT 1834.1000 2449.9800 1835.7000 2450.4600 ;
        RECT 1834.1000 2455.4200 1835.7000 2455.9000 ;
        RECT 1789.1000 2444.5400 1790.7000 2445.0200 ;
        RECT 1789.1000 2449.9800 1790.7000 2450.4600 ;
        RECT 1789.1000 2455.4200 1790.7000 2455.9000 ;
        RECT 1834.1000 2433.6600 1835.7000 2434.1400 ;
        RECT 1834.1000 2439.1000 1835.7000 2439.5800 ;
        RECT 1834.1000 2417.3400 1835.7000 2417.8200 ;
        RECT 1834.1000 2422.7800 1835.7000 2423.2600 ;
        RECT 1834.1000 2428.2200 1835.7000 2428.7000 ;
        RECT 1789.1000 2433.6600 1790.7000 2434.1400 ;
        RECT 1789.1000 2439.1000 1790.7000 2439.5800 ;
        RECT 1789.1000 2417.3400 1790.7000 2417.8200 ;
        RECT 1789.1000 2422.7800 1790.7000 2423.2600 ;
        RECT 1789.1000 2428.2200 1790.7000 2428.7000 ;
        RECT 1744.1000 2444.5400 1745.7000 2445.0200 ;
        RECT 1744.1000 2449.9800 1745.7000 2450.4600 ;
        RECT 1736.3400 2444.5400 1737.9400 2445.0200 ;
        RECT 1736.3400 2449.9800 1737.9400 2450.4600 ;
        RECT 1736.3400 2455.4200 1737.9400 2455.9000 ;
        RECT 1744.1000 2455.4200 1745.7000 2455.9000 ;
        RECT 1744.1000 2433.6600 1745.7000 2434.1400 ;
        RECT 1744.1000 2439.1000 1745.7000 2439.5800 ;
        RECT 1736.3400 2433.6600 1737.9400 2434.1400 ;
        RECT 1736.3400 2439.1000 1737.9400 2439.5800 ;
        RECT 1744.1000 2417.3400 1745.7000 2417.8200 ;
        RECT 1744.1000 2422.7800 1745.7000 2423.2600 ;
        RECT 1736.3400 2417.3400 1737.9400 2417.8200 ;
        RECT 1736.3400 2422.7800 1737.9400 2423.2600 ;
        RECT 1736.3400 2428.2200 1737.9400 2428.7000 ;
        RECT 1744.1000 2428.2200 1745.7000 2428.7000 ;
        RECT 1834.1000 2401.0200 1835.7000 2401.5000 ;
        RECT 1834.1000 2406.4600 1835.7000 2406.9400 ;
        RECT 1834.1000 2411.9000 1835.7000 2412.3800 ;
        RECT 1834.1000 2390.1400 1835.7000 2390.6200 ;
        RECT 1834.1000 2395.5800 1835.7000 2396.0600 ;
        RECT 1789.1000 2401.0200 1790.7000 2401.5000 ;
        RECT 1789.1000 2406.4600 1790.7000 2406.9400 ;
        RECT 1789.1000 2411.9000 1790.7000 2412.3800 ;
        RECT 1789.1000 2390.1400 1790.7000 2390.6200 ;
        RECT 1789.1000 2395.5800 1790.7000 2396.0600 ;
        RECT 1834.1000 2373.8200 1835.7000 2374.3000 ;
        RECT 1834.1000 2379.2600 1835.7000 2379.7400 ;
        RECT 1834.1000 2384.7000 1835.7000 2385.1800 ;
        RECT 1834.1000 2362.9400 1835.7000 2363.4200 ;
        RECT 1834.1000 2368.3800 1835.7000 2368.8600 ;
        RECT 1789.1000 2373.8200 1790.7000 2374.3000 ;
        RECT 1789.1000 2379.2600 1790.7000 2379.7400 ;
        RECT 1789.1000 2384.7000 1790.7000 2385.1800 ;
        RECT 1789.1000 2362.9400 1790.7000 2363.4200 ;
        RECT 1789.1000 2368.3800 1790.7000 2368.8600 ;
        RECT 1744.1000 2401.0200 1745.7000 2401.5000 ;
        RECT 1744.1000 2406.4600 1745.7000 2406.9400 ;
        RECT 1744.1000 2411.9000 1745.7000 2412.3800 ;
        RECT 1736.3400 2401.0200 1737.9400 2401.5000 ;
        RECT 1736.3400 2406.4600 1737.9400 2406.9400 ;
        RECT 1736.3400 2411.9000 1737.9400 2412.3800 ;
        RECT 1744.1000 2390.1400 1745.7000 2390.6200 ;
        RECT 1744.1000 2395.5800 1745.7000 2396.0600 ;
        RECT 1736.3400 2390.1400 1737.9400 2390.6200 ;
        RECT 1736.3400 2395.5800 1737.9400 2396.0600 ;
        RECT 1744.1000 2373.8200 1745.7000 2374.3000 ;
        RECT 1744.1000 2379.2600 1745.7000 2379.7400 ;
        RECT 1744.1000 2384.7000 1745.7000 2385.1800 ;
        RECT 1736.3400 2373.8200 1737.9400 2374.3000 ;
        RECT 1736.3400 2379.2600 1737.9400 2379.7400 ;
        RECT 1736.3400 2384.7000 1737.9400 2385.1800 ;
        RECT 1744.1000 2362.9400 1745.7000 2363.4200 ;
        RECT 1744.1000 2368.3800 1745.7000 2368.8600 ;
        RECT 1736.3400 2362.9400 1737.9400 2363.4200 ;
        RECT 1736.3400 2368.3800 1737.9400 2368.8600 ;
        RECT 1933.8400 2346.6200 1935.4400 2347.1000 ;
        RECT 1933.8400 2352.0600 1935.4400 2352.5400 ;
        RECT 1933.8400 2357.5000 1935.4400 2357.9800 ;
        RECT 1924.1000 2346.6200 1925.7000 2347.1000 ;
        RECT 1924.1000 2352.0600 1925.7000 2352.5400 ;
        RECT 1924.1000 2357.5000 1925.7000 2357.9800 ;
        RECT 1933.8400 2335.7400 1935.4400 2336.2200 ;
        RECT 1933.8400 2341.1800 1935.4400 2341.6600 ;
        RECT 1924.1000 2335.7400 1925.7000 2336.2200 ;
        RECT 1924.1000 2341.1800 1925.7000 2341.6600 ;
        RECT 1933.8400 2319.4200 1935.4400 2319.9000 ;
        RECT 1933.8400 2324.8600 1935.4400 2325.3400 ;
        RECT 1933.8400 2330.3000 1935.4400 2330.7800 ;
        RECT 1924.1000 2319.4200 1925.7000 2319.9000 ;
        RECT 1924.1000 2324.8600 1925.7000 2325.3400 ;
        RECT 1924.1000 2330.3000 1925.7000 2330.7800 ;
        RECT 1933.8400 2308.5400 1935.4400 2309.0200 ;
        RECT 1933.8400 2313.9800 1935.4400 2314.4600 ;
        RECT 1924.1000 2308.5400 1925.7000 2309.0200 ;
        RECT 1924.1000 2313.9800 1925.7000 2314.4600 ;
        RECT 1879.1000 2346.6200 1880.7000 2347.1000 ;
        RECT 1879.1000 2352.0600 1880.7000 2352.5400 ;
        RECT 1879.1000 2357.5000 1880.7000 2357.9800 ;
        RECT 1879.1000 2335.7400 1880.7000 2336.2200 ;
        RECT 1879.1000 2341.1800 1880.7000 2341.6600 ;
        RECT 1879.1000 2319.4200 1880.7000 2319.9000 ;
        RECT 1879.1000 2324.8600 1880.7000 2325.3400 ;
        RECT 1879.1000 2330.3000 1880.7000 2330.7800 ;
        RECT 1879.1000 2308.5400 1880.7000 2309.0200 ;
        RECT 1879.1000 2313.9800 1880.7000 2314.4600 ;
        RECT 1933.8400 2292.2200 1935.4400 2292.7000 ;
        RECT 1933.8400 2297.6600 1935.4400 2298.1400 ;
        RECT 1933.8400 2303.1000 1935.4400 2303.5800 ;
        RECT 1924.1000 2292.2200 1925.7000 2292.7000 ;
        RECT 1924.1000 2297.6600 1925.7000 2298.1400 ;
        RECT 1924.1000 2303.1000 1925.7000 2303.5800 ;
        RECT 1933.8400 2281.3400 1935.4400 2281.8200 ;
        RECT 1933.8400 2286.7800 1935.4400 2287.2600 ;
        RECT 1924.1000 2281.3400 1925.7000 2281.8200 ;
        RECT 1924.1000 2286.7800 1925.7000 2287.2600 ;
        RECT 1933.8400 2265.0200 1935.4400 2265.5000 ;
        RECT 1933.8400 2270.4600 1935.4400 2270.9400 ;
        RECT 1933.8400 2275.9000 1935.4400 2276.3800 ;
        RECT 1924.1000 2265.0200 1925.7000 2265.5000 ;
        RECT 1924.1000 2270.4600 1925.7000 2270.9400 ;
        RECT 1924.1000 2275.9000 1925.7000 2276.3800 ;
        RECT 1924.1000 2259.5800 1925.7000 2260.0600 ;
        RECT 1933.8400 2259.5800 1935.4400 2260.0600 ;
        RECT 1879.1000 2292.2200 1880.7000 2292.7000 ;
        RECT 1879.1000 2297.6600 1880.7000 2298.1400 ;
        RECT 1879.1000 2303.1000 1880.7000 2303.5800 ;
        RECT 1879.1000 2281.3400 1880.7000 2281.8200 ;
        RECT 1879.1000 2286.7800 1880.7000 2287.2600 ;
        RECT 1879.1000 2265.0200 1880.7000 2265.5000 ;
        RECT 1879.1000 2270.4600 1880.7000 2270.9400 ;
        RECT 1879.1000 2275.9000 1880.7000 2276.3800 ;
        RECT 1879.1000 2259.5800 1880.7000 2260.0600 ;
        RECT 1834.1000 2346.6200 1835.7000 2347.1000 ;
        RECT 1834.1000 2352.0600 1835.7000 2352.5400 ;
        RECT 1834.1000 2357.5000 1835.7000 2357.9800 ;
        RECT 1834.1000 2335.7400 1835.7000 2336.2200 ;
        RECT 1834.1000 2341.1800 1835.7000 2341.6600 ;
        RECT 1789.1000 2346.6200 1790.7000 2347.1000 ;
        RECT 1789.1000 2352.0600 1790.7000 2352.5400 ;
        RECT 1789.1000 2357.5000 1790.7000 2357.9800 ;
        RECT 1789.1000 2335.7400 1790.7000 2336.2200 ;
        RECT 1789.1000 2341.1800 1790.7000 2341.6600 ;
        RECT 1834.1000 2319.4200 1835.7000 2319.9000 ;
        RECT 1834.1000 2324.8600 1835.7000 2325.3400 ;
        RECT 1834.1000 2330.3000 1835.7000 2330.7800 ;
        RECT 1834.1000 2308.5400 1835.7000 2309.0200 ;
        RECT 1834.1000 2313.9800 1835.7000 2314.4600 ;
        RECT 1789.1000 2319.4200 1790.7000 2319.9000 ;
        RECT 1789.1000 2324.8600 1790.7000 2325.3400 ;
        RECT 1789.1000 2330.3000 1790.7000 2330.7800 ;
        RECT 1789.1000 2308.5400 1790.7000 2309.0200 ;
        RECT 1789.1000 2313.9800 1790.7000 2314.4600 ;
        RECT 1744.1000 2346.6200 1745.7000 2347.1000 ;
        RECT 1744.1000 2352.0600 1745.7000 2352.5400 ;
        RECT 1744.1000 2357.5000 1745.7000 2357.9800 ;
        RECT 1736.3400 2346.6200 1737.9400 2347.1000 ;
        RECT 1736.3400 2352.0600 1737.9400 2352.5400 ;
        RECT 1736.3400 2357.5000 1737.9400 2357.9800 ;
        RECT 1744.1000 2335.7400 1745.7000 2336.2200 ;
        RECT 1744.1000 2341.1800 1745.7000 2341.6600 ;
        RECT 1736.3400 2335.7400 1737.9400 2336.2200 ;
        RECT 1736.3400 2341.1800 1737.9400 2341.6600 ;
        RECT 1744.1000 2319.4200 1745.7000 2319.9000 ;
        RECT 1744.1000 2324.8600 1745.7000 2325.3400 ;
        RECT 1744.1000 2330.3000 1745.7000 2330.7800 ;
        RECT 1736.3400 2319.4200 1737.9400 2319.9000 ;
        RECT 1736.3400 2324.8600 1737.9400 2325.3400 ;
        RECT 1736.3400 2330.3000 1737.9400 2330.7800 ;
        RECT 1744.1000 2308.5400 1745.7000 2309.0200 ;
        RECT 1744.1000 2313.9800 1745.7000 2314.4600 ;
        RECT 1736.3400 2308.5400 1737.9400 2309.0200 ;
        RECT 1736.3400 2313.9800 1737.9400 2314.4600 ;
        RECT 1834.1000 2292.2200 1835.7000 2292.7000 ;
        RECT 1834.1000 2297.6600 1835.7000 2298.1400 ;
        RECT 1834.1000 2303.1000 1835.7000 2303.5800 ;
        RECT 1834.1000 2281.3400 1835.7000 2281.8200 ;
        RECT 1834.1000 2286.7800 1835.7000 2287.2600 ;
        RECT 1789.1000 2292.2200 1790.7000 2292.7000 ;
        RECT 1789.1000 2297.6600 1790.7000 2298.1400 ;
        RECT 1789.1000 2303.1000 1790.7000 2303.5800 ;
        RECT 1789.1000 2281.3400 1790.7000 2281.8200 ;
        RECT 1789.1000 2286.7800 1790.7000 2287.2600 ;
        RECT 1834.1000 2265.0200 1835.7000 2265.5000 ;
        RECT 1834.1000 2270.4600 1835.7000 2270.9400 ;
        RECT 1834.1000 2275.9000 1835.7000 2276.3800 ;
        RECT 1834.1000 2259.5800 1835.7000 2260.0600 ;
        RECT 1789.1000 2265.0200 1790.7000 2265.5000 ;
        RECT 1789.1000 2270.4600 1790.7000 2270.9400 ;
        RECT 1789.1000 2275.9000 1790.7000 2276.3800 ;
        RECT 1789.1000 2259.5800 1790.7000 2260.0600 ;
        RECT 1744.1000 2292.2200 1745.7000 2292.7000 ;
        RECT 1744.1000 2297.6600 1745.7000 2298.1400 ;
        RECT 1744.1000 2303.1000 1745.7000 2303.5800 ;
        RECT 1736.3400 2292.2200 1737.9400 2292.7000 ;
        RECT 1736.3400 2297.6600 1737.9400 2298.1400 ;
        RECT 1736.3400 2303.1000 1737.9400 2303.5800 ;
        RECT 1744.1000 2281.3400 1745.7000 2281.8200 ;
        RECT 1744.1000 2286.7800 1745.7000 2287.2600 ;
        RECT 1736.3400 2281.3400 1737.9400 2281.8200 ;
        RECT 1736.3400 2286.7800 1737.9400 2287.2600 ;
        RECT 1744.1000 2265.0200 1745.7000 2265.5000 ;
        RECT 1744.1000 2270.4600 1745.7000 2270.9400 ;
        RECT 1744.1000 2275.9000 1745.7000 2276.3800 ;
        RECT 1736.3400 2265.0200 1737.9400 2265.5000 ;
        RECT 1736.3400 2270.4600 1737.9400 2270.9400 ;
        RECT 1736.3400 2275.9000 1737.9400 2276.3800 ;
        RECT 1736.3400 2259.5800 1737.9400 2260.0600 ;
        RECT 1744.1000 2259.5800 1745.7000 2260.0600 ;
        RECT 1730.7800 2461.8900 1941.0000 2463.4900 ;
        RECT 1730.7800 2255.3900 1941.0000 2256.9900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 2249.9600 1737.9400 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 2468.0000 1737.9400 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 2249.9600 1935.4400 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 2468.0000 1935.4400 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2255.3900 1732.3800 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2255.3900 1941.0000 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2461.8900 1732.3800 2463.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2461.8900 1941.0000 2463.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 2025.7500 1925.7000 2233.8500 ;
        RECT 1879.1000 2025.7500 1880.7000 2233.8500 ;
        RECT 1834.1000 2025.7500 1835.7000 2233.8500 ;
        RECT 1789.1000 2025.7500 1790.7000 2233.8500 ;
        RECT 1744.1000 2025.7500 1745.7000 2233.8500 ;
        RECT 1933.8400 2020.3200 1935.4400 2239.9600 ;
        RECT 1736.3400 2020.3200 1737.9400 2239.9600 ;
      LAYER met3 ;
        RECT 1933.8400 2214.9000 1935.4400 2215.3800 ;
        RECT 1933.8400 2220.3400 1935.4400 2220.8200 ;
        RECT 1924.1000 2214.9000 1925.7000 2215.3800 ;
        RECT 1924.1000 2220.3400 1925.7000 2220.8200 ;
        RECT 1924.1000 2225.7800 1925.7000 2226.2600 ;
        RECT 1933.8400 2225.7800 1935.4400 2226.2600 ;
        RECT 1933.8400 2204.0200 1935.4400 2204.5000 ;
        RECT 1933.8400 2209.4600 1935.4400 2209.9400 ;
        RECT 1924.1000 2204.0200 1925.7000 2204.5000 ;
        RECT 1924.1000 2209.4600 1925.7000 2209.9400 ;
        RECT 1933.8400 2187.7000 1935.4400 2188.1800 ;
        RECT 1933.8400 2193.1400 1935.4400 2193.6200 ;
        RECT 1924.1000 2187.7000 1925.7000 2188.1800 ;
        RECT 1924.1000 2193.1400 1925.7000 2193.6200 ;
        RECT 1924.1000 2198.5800 1925.7000 2199.0600 ;
        RECT 1933.8400 2198.5800 1935.4400 2199.0600 ;
        RECT 1879.1000 2214.9000 1880.7000 2215.3800 ;
        RECT 1879.1000 2220.3400 1880.7000 2220.8200 ;
        RECT 1879.1000 2225.7800 1880.7000 2226.2600 ;
        RECT 1879.1000 2204.0200 1880.7000 2204.5000 ;
        RECT 1879.1000 2209.4600 1880.7000 2209.9400 ;
        RECT 1879.1000 2187.7000 1880.7000 2188.1800 ;
        RECT 1879.1000 2193.1400 1880.7000 2193.6200 ;
        RECT 1879.1000 2198.5800 1880.7000 2199.0600 ;
        RECT 1933.8400 2171.3800 1935.4400 2171.8600 ;
        RECT 1933.8400 2176.8200 1935.4400 2177.3000 ;
        RECT 1933.8400 2182.2600 1935.4400 2182.7400 ;
        RECT 1924.1000 2171.3800 1925.7000 2171.8600 ;
        RECT 1924.1000 2176.8200 1925.7000 2177.3000 ;
        RECT 1924.1000 2182.2600 1925.7000 2182.7400 ;
        RECT 1933.8400 2160.5000 1935.4400 2160.9800 ;
        RECT 1933.8400 2165.9400 1935.4400 2166.4200 ;
        RECT 1924.1000 2160.5000 1925.7000 2160.9800 ;
        RECT 1924.1000 2165.9400 1925.7000 2166.4200 ;
        RECT 1933.8400 2144.1800 1935.4400 2144.6600 ;
        RECT 1933.8400 2149.6200 1935.4400 2150.1000 ;
        RECT 1933.8400 2155.0600 1935.4400 2155.5400 ;
        RECT 1924.1000 2144.1800 1925.7000 2144.6600 ;
        RECT 1924.1000 2149.6200 1925.7000 2150.1000 ;
        RECT 1924.1000 2155.0600 1925.7000 2155.5400 ;
        RECT 1933.8400 2133.3000 1935.4400 2133.7800 ;
        RECT 1933.8400 2138.7400 1935.4400 2139.2200 ;
        RECT 1924.1000 2133.3000 1925.7000 2133.7800 ;
        RECT 1924.1000 2138.7400 1925.7000 2139.2200 ;
        RECT 1879.1000 2171.3800 1880.7000 2171.8600 ;
        RECT 1879.1000 2176.8200 1880.7000 2177.3000 ;
        RECT 1879.1000 2182.2600 1880.7000 2182.7400 ;
        RECT 1879.1000 2160.5000 1880.7000 2160.9800 ;
        RECT 1879.1000 2165.9400 1880.7000 2166.4200 ;
        RECT 1879.1000 2144.1800 1880.7000 2144.6600 ;
        RECT 1879.1000 2149.6200 1880.7000 2150.1000 ;
        RECT 1879.1000 2155.0600 1880.7000 2155.5400 ;
        RECT 1879.1000 2133.3000 1880.7000 2133.7800 ;
        RECT 1879.1000 2138.7400 1880.7000 2139.2200 ;
        RECT 1834.1000 2214.9000 1835.7000 2215.3800 ;
        RECT 1834.1000 2220.3400 1835.7000 2220.8200 ;
        RECT 1834.1000 2225.7800 1835.7000 2226.2600 ;
        RECT 1789.1000 2214.9000 1790.7000 2215.3800 ;
        RECT 1789.1000 2220.3400 1790.7000 2220.8200 ;
        RECT 1789.1000 2225.7800 1790.7000 2226.2600 ;
        RECT 1834.1000 2204.0200 1835.7000 2204.5000 ;
        RECT 1834.1000 2209.4600 1835.7000 2209.9400 ;
        RECT 1834.1000 2187.7000 1835.7000 2188.1800 ;
        RECT 1834.1000 2193.1400 1835.7000 2193.6200 ;
        RECT 1834.1000 2198.5800 1835.7000 2199.0600 ;
        RECT 1789.1000 2204.0200 1790.7000 2204.5000 ;
        RECT 1789.1000 2209.4600 1790.7000 2209.9400 ;
        RECT 1789.1000 2187.7000 1790.7000 2188.1800 ;
        RECT 1789.1000 2193.1400 1790.7000 2193.6200 ;
        RECT 1789.1000 2198.5800 1790.7000 2199.0600 ;
        RECT 1744.1000 2214.9000 1745.7000 2215.3800 ;
        RECT 1744.1000 2220.3400 1745.7000 2220.8200 ;
        RECT 1736.3400 2214.9000 1737.9400 2215.3800 ;
        RECT 1736.3400 2220.3400 1737.9400 2220.8200 ;
        RECT 1736.3400 2225.7800 1737.9400 2226.2600 ;
        RECT 1744.1000 2225.7800 1745.7000 2226.2600 ;
        RECT 1744.1000 2204.0200 1745.7000 2204.5000 ;
        RECT 1744.1000 2209.4600 1745.7000 2209.9400 ;
        RECT 1736.3400 2204.0200 1737.9400 2204.5000 ;
        RECT 1736.3400 2209.4600 1737.9400 2209.9400 ;
        RECT 1744.1000 2187.7000 1745.7000 2188.1800 ;
        RECT 1744.1000 2193.1400 1745.7000 2193.6200 ;
        RECT 1736.3400 2187.7000 1737.9400 2188.1800 ;
        RECT 1736.3400 2193.1400 1737.9400 2193.6200 ;
        RECT 1736.3400 2198.5800 1737.9400 2199.0600 ;
        RECT 1744.1000 2198.5800 1745.7000 2199.0600 ;
        RECT 1834.1000 2171.3800 1835.7000 2171.8600 ;
        RECT 1834.1000 2176.8200 1835.7000 2177.3000 ;
        RECT 1834.1000 2182.2600 1835.7000 2182.7400 ;
        RECT 1834.1000 2160.5000 1835.7000 2160.9800 ;
        RECT 1834.1000 2165.9400 1835.7000 2166.4200 ;
        RECT 1789.1000 2171.3800 1790.7000 2171.8600 ;
        RECT 1789.1000 2176.8200 1790.7000 2177.3000 ;
        RECT 1789.1000 2182.2600 1790.7000 2182.7400 ;
        RECT 1789.1000 2160.5000 1790.7000 2160.9800 ;
        RECT 1789.1000 2165.9400 1790.7000 2166.4200 ;
        RECT 1834.1000 2144.1800 1835.7000 2144.6600 ;
        RECT 1834.1000 2149.6200 1835.7000 2150.1000 ;
        RECT 1834.1000 2155.0600 1835.7000 2155.5400 ;
        RECT 1834.1000 2133.3000 1835.7000 2133.7800 ;
        RECT 1834.1000 2138.7400 1835.7000 2139.2200 ;
        RECT 1789.1000 2144.1800 1790.7000 2144.6600 ;
        RECT 1789.1000 2149.6200 1790.7000 2150.1000 ;
        RECT 1789.1000 2155.0600 1790.7000 2155.5400 ;
        RECT 1789.1000 2133.3000 1790.7000 2133.7800 ;
        RECT 1789.1000 2138.7400 1790.7000 2139.2200 ;
        RECT 1744.1000 2171.3800 1745.7000 2171.8600 ;
        RECT 1744.1000 2176.8200 1745.7000 2177.3000 ;
        RECT 1744.1000 2182.2600 1745.7000 2182.7400 ;
        RECT 1736.3400 2171.3800 1737.9400 2171.8600 ;
        RECT 1736.3400 2176.8200 1737.9400 2177.3000 ;
        RECT 1736.3400 2182.2600 1737.9400 2182.7400 ;
        RECT 1744.1000 2160.5000 1745.7000 2160.9800 ;
        RECT 1744.1000 2165.9400 1745.7000 2166.4200 ;
        RECT 1736.3400 2160.5000 1737.9400 2160.9800 ;
        RECT 1736.3400 2165.9400 1737.9400 2166.4200 ;
        RECT 1744.1000 2144.1800 1745.7000 2144.6600 ;
        RECT 1744.1000 2149.6200 1745.7000 2150.1000 ;
        RECT 1744.1000 2155.0600 1745.7000 2155.5400 ;
        RECT 1736.3400 2144.1800 1737.9400 2144.6600 ;
        RECT 1736.3400 2149.6200 1737.9400 2150.1000 ;
        RECT 1736.3400 2155.0600 1737.9400 2155.5400 ;
        RECT 1744.1000 2133.3000 1745.7000 2133.7800 ;
        RECT 1744.1000 2138.7400 1745.7000 2139.2200 ;
        RECT 1736.3400 2133.3000 1737.9400 2133.7800 ;
        RECT 1736.3400 2138.7400 1737.9400 2139.2200 ;
        RECT 1933.8400 2116.9800 1935.4400 2117.4600 ;
        RECT 1933.8400 2122.4200 1935.4400 2122.9000 ;
        RECT 1933.8400 2127.8600 1935.4400 2128.3400 ;
        RECT 1924.1000 2116.9800 1925.7000 2117.4600 ;
        RECT 1924.1000 2122.4200 1925.7000 2122.9000 ;
        RECT 1924.1000 2127.8600 1925.7000 2128.3400 ;
        RECT 1933.8400 2106.1000 1935.4400 2106.5800 ;
        RECT 1933.8400 2111.5400 1935.4400 2112.0200 ;
        RECT 1924.1000 2106.1000 1925.7000 2106.5800 ;
        RECT 1924.1000 2111.5400 1925.7000 2112.0200 ;
        RECT 1933.8400 2089.7800 1935.4400 2090.2600 ;
        RECT 1933.8400 2095.2200 1935.4400 2095.7000 ;
        RECT 1933.8400 2100.6600 1935.4400 2101.1400 ;
        RECT 1924.1000 2089.7800 1925.7000 2090.2600 ;
        RECT 1924.1000 2095.2200 1925.7000 2095.7000 ;
        RECT 1924.1000 2100.6600 1925.7000 2101.1400 ;
        RECT 1933.8400 2078.9000 1935.4400 2079.3800 ;
        RECT 1933.8400 2084.3400 1935.4400 2084.8200 ;
        RECT 1924.1000 2078.9000 1925.7000 2079.3800 ;
        RECT 1924.1000 2084.3400 1925.7000 2084.8200 ;
        RECT 1879.1000 2116.9800 1880.7000 2117.4600 ;
        RECT 1879.1000 2122.4200 1880.7000 2122.9000 ;
        RECT 1879.1000 2127.8600 1880.7000 2128.3400 ;
        RECT 1879.1000 2106.1000 1880.7000 2106.5800 ;
        RECT 1879.1000 2111.5400 1880.7000 2112.0200 ;
        RECT 1879.1000 2089.7800 1880.7000 2090.2600 ;
        RECT 1879.1000 2095.2200 1880.7000 2095.7000 ;
        RECT 1879.1000 2100.6600 1880.7000 2101.1400 ;
        RECT 1879.1000 2078.9000 1880.7000 2079.3800 ;
        RECT 1879.1000 2084.3400 1880.7000 2084.8200 ;
        RECT 1933.8400 2062.5800 1935.4400 2063.0600 ;
        RECT 1933.8400 2068.0200 1935.4400 2068.5000 ;
        RECT 1933.8400 2073.4600 1935.4400 2073.9400 ;
        RECT 1924.1000 2062.5800 1925.7000 2063.0600 ;
        RECT 1924.1000 2068.0200 1925.7000 2068.5000 ;
        RECT 1924.1000 2073.4600 1925.7000 2073.9400 ;
        RECT 1933.8400 2051.7000 1935.4400 2052.1800 ;
        RECT 1933.8400 2057.1400 1935.4400 2057.6200 ;
        RECT 1924.1000 2051.7000 1925.7000 2052.1800 ;
        RECT 1924.1000 2057.1400 1925.7000 2057.6200 ;
        RECT 1933.8400 2035.3800 1935.4400 2035.8600 ;
        RECT 1933.8400 2040.8200 1935.4400 2041.3000 ;
        RECT 1933.8400 2046.2600 1935.4400 2046.7400 ;
        RECT 1924.1000 2035.3800 1925.7000 2035.8600 ;
        RECT 1924.1000 2040.8200 1925.7000 2041.3000 ;
        RECT 1924.1000 2046.2600 1925.7000 2046.7400 ;
        RECT 1924.1000 2029.9400 1925.7000 2030.4200 ;
        RECT 1933.8400 2029.9400 1935.4400 2030.4200 ;
        RECT 1879.1000 2062.5800 1880.7000 2063.0600 ;
        RECT 1879.1000 2068.0200 1880.7000 2068.5000 ;
        RECT 1879.1000 2073.4600 1880.7000 2073.9400 ;
        RECT 1879.1000 2051.7000 1880.7000 2052.1800 ;
        RECT 1879.1000 2057.1400 1880.7000 2057.6200 ;
        RECT 1879.1000 2035.3800 1880.7000 2035.8600 ;
        RECT 1879.1000 2040.8200 1880.7000 2041.3000 ;
        RECT 1879.1000 2046.2600 1880.7000 2046.7400 ;
        RECT 1879.1000 2029.9400 1880.7000 2030.4200 ;
        RECT 1834.1000 2116.9800 1835.7000 2117.4600 ;
        RECT 1834.1000 2122.4200 1835.7000 2122.9000 ;
        RECT 1834.1000 2127.8600 1835.7000 2128.3400 ;
        RECT 1834.1000 2106.1000 1835.7000 2106.5800 ;
        RECT 1834.1000 2111.5400 1835.7000 2112.0200 ;
        RECT 1789.1000 2116.9800 1790.7000 2117.4600 ;
        RECT 1789.1000 2122.4200 1790.7000 2122.9000 ;
        RECT 1789.1000 2127.8600 1790.7000 2128.3400 ;
        RECT 1789.1000 2106.1000 1790.7000 2106.5800 ;
        RECT 1789.1000 2111.5400 1790.7000 2112.0200 ;
        RECT 1834.1000 2089.7800 1835.7000 2090.2600 ;
        RECT 1834.1000 2095.2200 1835.7000 2095.7000 ;
        RECT 1834.1000 2100.6600 1835.7000 2101.1400 ;
        RECT 1834.1000 2078.9000 1835.7000 2079.3800 ;
        RECT 1834.1000 2084.3400 1835.7000 2084.8200 ;
        RECT 1789.1000 2089.7800 1790.7000 2090.2600 ;
        RECT 1789.1000 2095.2200 1790.7000 2095.7000 ;
        RECT 1789.1000 2100.6600 1790.7000 2101.1400 ;
        RECT 1789.1000 2078.9000 1790.7000 2079.3800 ;
        RECT 1789.1000 2084.3400 1790.7000 2084.8200 ;
        RECT 1744.1000 2116.9800 1745.7000 2117.4600 ;
        RECT 1744.1000 2122.4200 1745.7000 2122.9000 ;
        RECT 1744.1000 2127.8600 1745.7000 2128.3400 ;
        RECT 1736.3400 2116.9800 1737.9400 2117.4600 ;
        RECT 1736.3400 2122.4200 1737.9400 2122.9000 ;
        RECT 1736.3400 2127.8600 1737.9400 2128.3400 ;
        RECT 1744.1000 2106.1000 1745.7000 2106.5800 ;
        RECT 1744.1000 2111.5400 1745.7000 2112.0200 ;
        RECT 1736.3400 2106.1000 1737.9400 2106.5800 ;
        RECT 1736.3400 2111.5400 1737.9400 2112.0200 ;
        RECT 1744.1000 2089.7800 1745.7000 2090.2600 ;
        RECT 1744.1000 2095.2200 1745.7000 2095.7000 ;
        RECT 1744.1000 2100.6600 1745.7000 2101.1400 ;
        RECT 1736.3400 2089.7800 1737.9400 2090.2600 ;
        RECT 1736.3400 2095.2200 1737.9400 2095.7000 ;
        RECT 1736.3400 2100.6600 1737.9400 2101.1400 ;
        RECT 1744.1000 2078.9000 1745.7000 2079.3800 ;
        RECT 1744.1000 2084.3400 1745.7000 2084.8200 ;
        RECT 1736.3400 2078.9000 1737.9400 2079.3800 ;
        RECT 1736.3400 2084.3400 1737.9400 2084.8200 ;
        RECT 1834.1000 2062.5800 1835.7000 2063.0600 ;
        RECT 1834.1000 2068.0200 1835.7000 2068.5000 ;
        RECT 1834.1000 2073.4600 1835.7000 2073.9400 ;
        RECT 1834.1000 2051.7000 1835.7000 2052.1800 ;
        RECT 1834.1000 2057.1400 1835.7000 2057.6200 ;
        RECT 1789.1000 2062.5800 1790.7000 2063.0600 ;
        RECT 1789.1000 2068.0200 1790.7000 2068.5000 ;
        RECT 1789.1000 2073.4600 1790.7000 2073.9400 ;
        RECT 1789.1000 2051.7000 1790.7000 2052.1800 ;
        RECT 1789.1000 2057.1400 1790.7000 2057.6200 ;
        RECT 1834.1000 2035.3800 1835.7000 2035.8600 ;
        RECT 1834.1000 2040.8200 1835.7000 2041.3000 ;
        RECT 1834.1000 2046.2600 1835.7000 2046.7400 ;
        RECT 1834.1000 2029.9400 1835.7000 2030.4200 ;
        RECT 1789.1000 2035.3800 1790.7000 2035.8600 ;
        RECT 1789.1000 2040.8200 1790.7000 2041.3000 ;
        RECT 1789.1000 2046.2600 1790.7000 2046.7400 ;
        RECT 1789.1000 2029.9400 1790.7000 2030.4200 ;
        RECT 1744.1000 2062.5800 1745.7000 2063.0600 ;
        RECT 1744.1000 2068.0200 1745.7000 2068.5000 ;
        RECT 1744.1000 2073.4600 1745.7000 2073.9400 ;
        RECT 1736.3400 2062.5800 1737.9400 2063.0600 ;
        RECT 1736.3400 2068.0200 1737.9400 2068.5000 ;
        RECT 1736.3400 2073.4600 1737.9400 2073.9400 ;
        RECT 1744.1000 2051.7000 1745.7000 2052.1800 ;
        RECT 1744.1000 2057.1400 1745.7000 2057.6200 ;
        RECT 1736.3400 2051.7000 1737.9400 2052.1800 ;
        RECT 1736.3400 2057.1400 1737.9400 2057.6200 ;
        RECT 1744.1000 2035.3800 1745.7000 2035.8600 ;
        RECT 1744.1000 2040.8200 1745.7000 2041.3000 ;
        RECT 1744.1000 2046.2600 1745.7000 2046.7400 ;
        RECT 1736.3400 2035.3800 1737.9400 2035.8600 ;
        RECT 1736.3400 2040.8200 1737.9400 2041.3000 ;
        RECT 1736.3400 2046.2600 1737.9400 2046.7400 ;
        RECT 1736.3400 2029.9400 1737.9400 2030.4200 ;
        RECT 1744.1000 2029.9400 1745.7000 2030.4200 ;
        RECT 1730.7800 2232.2500 1941.0000 2233.8500 ;
        RECT 1730.7800 2025.7500 1941.0000 2027.3500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 2020.3200 1737.9400 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 2238.3600 1737.9400 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 2020.3200 1935.4400 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 2238.3600 1935.4400 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2025.7500 1732.3800 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2025.7500 1941.0000 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2232.2500 1732.3800 2233.8500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2232.2500 1941.0000 2233.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 1796.1100 1925.7000 2004.2100 ;
        RECT 1879.1000 1796.1100 1880.7000 2004.2100 ;
        RECT 1834.1000 1796.1100 1835.7000 2004.2100 ;
        RECT 1789.1000 1796.1100 1790.7000 2004.2100 ;
        RECT 1744.1000 1796.1100 1745.7000 2004.2100 ;
        RECT 1933.8400 1790.6800 1935.4400 2010.3200 ;
        RECT 1736.3400 1790.6800 1737.9400 2010.3200 ;
      LAYER met3 ;
        RECT 1933.8400 1985.2600 1935.4400 1985.7400 ;
        RECT 1933.8400 1990.7000 1935.4400 1991.1800 ;
        RECT 1924.1000 1985.2600 1925.7000 1985.7400 ;
        RECT 1924.1000 1990.7000 1925.7000 1991.1800 ;
        RECT 1924.1000 1996.1400 1925.7000 1996.6200 ;
        RECT 1933.8400 1996.1400 1935.4400 1996.6200 ;
        RECT 1933.8400 1974.3800 1935.4400 1974.8600 ;
        RECT 1933.8400 1979.8200 1935.4400 1980.3000 ;
        RECT 1924.1000 1974.3800 1925.7000 1974.8600 ;
        RECT 1924.1000 1979.8200 1925.7000 1980.3000 ;
        RECT 1933.8400 1958.0600 1935.4400 1958.5400 ;
        RECT 1933.8400 1963.5000 1935.4400 1963.9800 ;
        RECT 1924.1000 1958.0600 1925.7000 1958.5400 ;
        RECT 1924.1000 1963.5000 1925.7000 1963.9800 ;
        RECT 1924.1000 1968.9400 1925.7000 1969.4200 ;
        RECT 1933.8400 1968.9400 1935.4400 1969.4200 ;
        RECT 1879.1000 1985.2600 1880.7000 1985.7400 ;
        RECT 1879.1000 1990.7000 1880.7000 1991.1800 ;
        RECT 1879.1000 1996.1400 1880.7000 1996.6200 ;
        RECT 1879.1000 1974.3800 1880.7000 1974.8600 ;
        RECT 1879.1000 1979.8200 1880.7000 1980.3000 ;
        RECT 1879.1000 1958.0600 1880.7000 1958.5400 ;
        RECT 1879.1000 1963.5000 1880.7000 1963.9800 ;
        RECT 1879.1000 1968.9400 1880.7000 1969.4200 ;
        RECT 1933.8400 1941.7400 1935.4400 1942.2200 ;
        RECT 1933.8400 1947.1800 1935.4400 1947.6600 ;
        RECT 1933.8400 1952.6200 1935.4400 1953.1000 ;
        RECT 1924.1000 1941.7400 1925.7000 1942.2200 ;
        RECT 1924.1000 1947.1800 1925.7000 1947.6600 ;
        RECT 1924.1000 1952.6200 1925.7000 1953.1000 ;
        RECT 1933.8400 1930.8600 1935.4400 1931.3400 ;
        RECT 1933.8400 1936.3000 1935.4400 1936.7800 ;
        RECT 1924.1000 1930.8600 1925.7000 1931.3400 ;
        RECT 1924.1000 1936.3000 1925.7000 1936.7800 ;
        RECT 1933.8400 1914.5400 1935.4400 1915.0200 ;
        RECT 1933.8400 1919.9800 1935.4400 1920.4600 ;
        RECT 1933.8400 1925.4200 1935.4400 1925.9000 ;
        RECT 1924.1000 1914.5400 1925.7000 1915.0200 ;
        RECT 1924.1000 1919.9800 1925.7000 1920.4600 ;
        RECT 1924.1000 1925.4200 1925.7000 1925.9000 ;
        RECT 1933.8400 1903.6600 1935.4400 1904.1400 ;
        RECT 1933.8400 1909.1000 1935.4400 1909.5800 ;
        RECT 1924.1000 1903.6600 1925.7000 1904.1400 ;
        RECT 1924.1000 1909.1000 1925.7000 1909.5800 ;
        RECT 1879.1000 1941.7400 1880.7000 1942.2200 ;
        RECT 1879.1000 1947.1800 1880.7000 1947.6600 ;
        RECT 1879.1000 1952.6200 1880.7000 1953.1000 ;
        RECT 1879.1000 1930.8600 1880.7000 1931.3400 ;
        RECT 1879.1000 1936.3000 1880.7000 1936.7800 ;
        RECT 1879.1000 1914.5400 1880.7000 1915.0200 ;
        RECT 1879.1000 1919.9800 1880.7000 1920.4600 ;
        RECT 1879.1000 1925.4200 1880.7000 1925.9000 ;
        RECT 1879.1000 1903.6600 1880.7000 1904.1400 ;
        RECT 1879.1000 1909.1000 1880.7000 1909.5800 ;
        RECT 1834.1000 1985.2600 1835.7000 1985.7400 ;
        RECT 1834.1000 1990.7000 1835.7000 1991.1800 ;
        RECT 1834.1000 1996.1400 1835.7000 1996.6200 ;
        RECT 1789.1000 1985.2600 1790.7000 1985.7400 ;
        RECT 1789.1000 1990.7000 1790.7000 1991.1800 ;
        RECT 1789.1000 1996.1400 1790.7000 1996.6200 ;
        RECT 1834.1000 1974.3800 1835.7000 1974.8600 ;
        RECT 1834.1000 1979.8200 1835.7000 1980.3000 ;
        RECT 1834.1000 1958.0600 1835.7000 1958.5400 ;
        RECT 1834.1000 1963.5000 1835.7000 1963.9800 ;
        RECT 1834.1000 1968.9400 1835.7000 1969.4200 ;
        RECT 1789.1000 1974.3800 1790.7000 1974.8600 ;
        RECT 1789.1000 1979.8200 1790.7000 1980.3000 ;
        RECT 1789.1000 1958.0600 1790.7000 1958.5400 ;
        RECT 1789.1000 1963.5000 1790.7000 1963.9800 ;
        RECT 1789.1000 1968.9400 1790.7000 1969.4200 ;
        RECT 1744.1000 1985.2600 1745.7000 1985.7400 ;
        RECT 1744.1000 1990.7000 1745.7000 1991.1800 ;
        RECT 1736.3400 1985.2600 1737.9400 1985.7400 ;
        RECT 1736.3400 1990.7000 1737.9400 1991.1800 ;
        RECT 1736.3400 1996.1400 1737.9400 1996.6200 ;
        RECT 1744.1000 1996.1400 1745.7000 1996.6200 ;
        RECT 1744.1000 1974.3800 1745.7000 1974.8600 ;
        RECT 1744.1000 1979.8200 1745.7000 1980.3000 ;
        RECT 1736.3400 1974.3800 1737.9400 1974.8600 ;
        RECT 1736.3400 1979.8200 1737.9400 1980.3000 ;
        RECT 1744.1000 1958.0600 1745.7000 1958.5400 ;
        RECT 1744.1000 1963.5000 1745.7000 1963.9800 ;
        RECT 1736.3400 1958.0600 1737.9400 1958.5400 ;
        RECT 1736.3400 1963.5000 1737.9400 1963.9800 ;
        RECT 1736.3400 1968.9400 1737.9400 1969.4200 ;
        RECT 1744.1000 1968.9400 1745.7000 1969.4200 ;
        RECT 1834.1000 1941.7400 1835.7000 1942.2200 ;
        RECT 1834.1000 1947.1800 1835.7000 1947.6600 ;
        RECT 1834.1000 1952.6200 1835.7000 1953.1000 ;
        RECT 1834.1000 1930.8600 1835.7000 1931.3400 ;
        RECT 1834.1000 1936.3000 1835.7000 1936.7800 ;
        RECT 1789.1000 1941.7400 1790.7000 1942.2200 ;
        RECT 1789.1000 1947.1800 1790.7000 1947.6600 ;
        RECT 1789.1000 1952.6200 1790.7000 1953.1000 ;
        RECT 1789.1000 1930.8600 1790.7000 1931.3400 ;
        RECT 1789.1000 1936.3000 1790.7000 1936.7800 ;
        RECT 1834.1000 1914.5400 1835.7000 1915.0200 ;
        RECT 1834.1000 1919.9800 1835.7000 1920.4600 ;
        RECT 1834.1000 1925.4200 1835.7000 1925.9000 ;
        RECT 1834.1000 1903.6600 1835.7000 1904.1400 ;
        RECT 1834.1000 1909.1000 1835.7000 1909.5800 ;
        RECT 1789.1000 1914.5400 1790.7000 1915.0200 ;
        RECT 1789.1000 1919.9800 1790.7000 1920.4600 ;
        RECT 1789.1000 1925.4200 1790.7000 1925.9000 ;
        RECT 1789.1000 1903.6600 1790.7000 1904.1400 ;
        RECT 1789.1000 1909.1000 1790.7000 1909.5800 ;
        RECT 1744.1000 1941.7400 1745.7000 1942.2200 ;
        RECT 1744.1000 1947.1800 1745.7000 1947.6600 ;
        RECT 1744.1000 1952.6200 1745.7000 1953.1000 ;
        RECT 1736.3400 1941.7400 1737.9400 1942.2200 ;
        RECT 1736.3400 1947.1800 1737.9400 1947.6600 ;
        RECT 1736.3400 1952.6200 1737.9400 1953.1000 ;
        RECT 1744.1000 1930.8600 1745.7000 1931.3400 ;
        RECT 1744.1000 1936.3000 1745.7000 1936.7800 ;
        RECT 1736.3400 1930.8600 1737.9400 1931.3400 ;
        RECT 1736.3400 1936.3000 1737.9400 1936.7800 ;
        RECT 1744.1000 1914.5400 1745.7000 1915.0200 ;
        RECT 1744.1000 1919.9800 1745.7000 1920.4600 ;
        RECT 1744.1000 1925.4200 1745.7000 1925.9000 ;
        RECT 1736.3400 1914.5400 1737.9400 1915.0200 ;
        RECT 1736.3400 1919.9800 1737.9400 1920.4600 ;
        RECT 1736.3400 1925.4200 1737.9400 1925.9000 ;
        RECT 1744.1000 1903.6600 1745.7000 1904.1400 ;
        RECT 1744.1000 1909.1000 1745.7000 1909.5800 ;
        RECT 1736.3400 1903.6600 1737.9400 1904.1400 ;
        RECT 1736.3400 1909.1000 1737.9400 1909.5800 ;
        RECT 1933.8400 1887.3400 1935.4400 1887.8200 ;
        RECT 1933.8400 1892.7800 1935.4400 1893.2600 ;
        RECT 1933.8400 1898.2200 1935.4400 1898.7000 ;
        RECT 1924.1000 1887.3400 1925.7000 1887.8200 ;
        RECT 1924.1000 1892.7800 1925.7000 1893.2600 ;
        RECT 1924.1000 1898.2200 1925.7000 1898.7000 ;
        RECT 1933.8400 1876.4600 1935.4400 1876.9400 ;
        RECT 1933.8400 1881.9000 1935.4400 1882.3800 ;
        RECT 1924.1000 1876.4600 1925.7000 1876.9400 ;
        RECT 1924.1000 1881.9000 1925.7000 1882.3800 ;
        RECT 1933.8400 1860.1400 1935.4400 1860.6200 ;
        RECT 1933.8400 1865.5800 1935.4400 1866.0600 ;
        RECT 1933.8400 1871.0200 1935.4400 1871.5000 ;
        RECT 1924.1000 1860.1400 1925.7000 1860.6200 ;
        RECT 1924.1000 1865.5800 1925.7000 1866.0600 ;
        RECT 1924.1000 1871.0200 1925.7000 1871.5000 ;
        RECT 1933.8400 1849.2600 1935.4400 1849.7400 ;
        RECT 1933.8400 1854.7000 1935.4400 1855.1800 ;
        RECT 1924.1000 1849.2600 1925.7000 1849.7400 ;
        RECT 1924.1000 1854.7000 1925.7000 1855.1800 ;
        RECT 1879.1000 1887.3400 1880.7000 1887.8200 ;
        RECT 1879.1000 1892.7800 1880.7000 1893.2600 ;
        RECT 1879.1000 1898.2200 1880.7000 1898.7000 ;
        RECT 1879.1000 1876.4600 1880.7000 1876.9400 ;
        RECT 1879.1000 1881.9000 1880.7000 1882.3800 ;
        RECT 1879.1000 1860.1400 1880.7000 1860.6200 ;
        RECT 1879.1000 1865.5800 1880.7000 1866.0600 ;
        RECT 1879.1000 1871.0200 1880.7000 1871.5000 ;
        RECT 1879.1000 1849.2600 1880.7000 1849.7400 ;
        RECT 1879.1000 1854.7000 1880.7000 1855.1800 ;
        RECT 1933.8400 1832.9400 1935.4400 1833.4200 ;
        RECT 1933.8400 1838.3800 1935.4400 1838.8600 ;
        RECT 1933.8400 1843.8200 1935.4400 1844.3000 ;
        RECT 1924.1000 1832.9400 1925.7000 1833.4200 ;
        RECT 1924.1000 1838.3800 1925.7000 1838.8600 ;
        RECT 1924.1000 1843.8200 1925.7000 1844.3000 ;
        RECT 1933.8400 1822.0600 1935.4400 1822.5400 ;
        RECT 1933.8400 1827.5000 1935.4400 1827.9800 ;
        RECT 1924.1000 1822.0600 1925.7000 1822.5400 ;
        RECT 1924.1000 1827.5000 1925.7000 1827.9800 ;
        RECT 1933.8400 1805.7400 1935.4400 1806.2200 ;
        RECT 1933.8400 1811.1800 1935.4400 1811.6600 ;
        RECT 1933.8400 1816.6200 1935.4400 1817.1000 ;
        RECT 1924.1000 1805.7400 1925.7000 1806.2200 ;
        RECT 1924.1000 1811.1800 1925.7000 1811.6600 ;
        RECT 1924.1000 1816.6200 1925.7000 1817.1000 ;
        RECT 1924.1000 1800.3000 1925.7000 1800.7800 ;
        RECT 1933.8400 1800.3000 1935.4400 1800.7800 ;
        RECT 1879.1000 1832.9400 1880.7000 1833.4200 ;
        RECT 1879.1000 1838.3800 1880.7000 1838.8600 ;
        RECT 1879.1000 1843.8200 1880.7000 1844.3000 ;
        RECT 1879.1000 1822.0600 1880.7000 1822.5400 ;
        RECT 1879.1000 1827.5000 1880.7000 1827.9800 ;
        RECT 1879.1000 1805.7400 1880.7000 1806.2200 ;
        RECT 1879.1000 1811.1800 1880.7000 1811.6600 ;
        RECT 1879.1000 1816.6200 1880.7000 1817.1000 ;
        RECT 1879.1000 1800.3000 1880.7000 1800.7800 ;
        RECT 1834.1000 1887.3400 1835.7000 1887.8200 ;
        RECT 1834.1000 1892.7800 1835.7000 1893.2600 ;
        RECT 1834.1000 1898.2200 1835.7000 1898.7000 ;
        RECT 1834.1000 1876.4600 1835.7000 1876.9400 ;
        RECT 1834.1000 1881.9000 1835.7000 1882.3800 ;
        RECT 1789.1000 1887.3400 1790.7000 1887.8200 ;
        RECT 1789.1000 1892.7800 1790.7000 1893.2600 ;
        RECT 1789.1000 1898.2200 1790.7000 1898.7000 ;
        RECT 1789.1000 1876.4600 1790.7000 1876.9400 ;
        RECT 1789.1000 1881.9000 1790.7000 1882.3800 ;
        RECT 1834.1000 1860.1400 1835.7000 1860.6200 ;
        RECT 1834.1000 1865.5800 1835.7000 1866.0600 ;
        RECT 1834.1000 1871.0200 1835.7000 1871.5000 ;
        RECT 1834.1000 1849.2600 1835.7000 1849.7400 ;
        RECT 1834.1000 1854.7000 1835.7000 1855.1800 ;
        RECT 1789.1000 1860.1400 1790.7000 1860.6200 ;
        RECT 1789.1000 1865.5800 1790.7000 1866.0600 ;
        RECT 1789.1000 1871.0200 1790.7000 1871.5000 ;
        RECT 1789.1000 1849.2600 1790.7000 1849.7400 ;
        RECT 1789.1000 1854.7000 1790.7000 1855.1800 ;
        RECT 1744.1000 1887.3400 1745.7000 1887.8200 ;
        RECT 1744.1000 1892.7800 1745.7000 1893.2600 ;
        RECT 1744.1000 1898.2200 1745.7000 1898.7000 ;
        RECT 1736.3400 1887.3400 1737.9400 1887.8200 ;
        RECT 1736.3400 1892.7800 1737.9400 1893.2600 ;
        RECT 1736.3400 1898.2200 1737.9400 1898.7000 ;
        RECT 1744.1000 1876.4600 1745.7000 1876.9400 ;
        RECT 1744.1000 1881.9000 1745.7000 1882.3800 ;
        RECT 1736.3400 1876.4600 1737.9400 1876.9400 ;
        RECT 1736.3400 1881.9000 1737.9400 1882.3800 ;
        RECT 1744.1000 1860.1400 1745.7000 1860.6200 ;
        RECT 1744.1000 1865.5800 1745.7000 1866.0600 ;
        RECT 1744.1000 1871.0200 1745.7000 1871.5000 ;
        RECT 1736.3400 1860.1400 1737.9400 1860.6200 ;
        RECT 1736.3400 1865.5800 1737.9400 1866.0600 ;
        RECT 1736.3400 1871.0200 1737.9400 1871.5000 ;
        RECT 1744.1000 1849.2600 1745.7000 1849.7400 ;
        RECT 1744.1000 1854.7000 1745.7000 1855.1800 ;
        RECT 1736.3400 1849.2600 1737.9400 1849.7400 ;
        RECT 1736.3400 1854.7000 1737.9400 1855.1800 ;
        RECT 1834.1000 1832.9400 1835.7000 1833.4200 ;
        RECT 1834.1000 1838.3800 1835.7000 1838.8600 ;
        RECT 1834.1000 1843.8200 1835.7000 1844.3000 ;
        RECT 1834.1000 1822.0600 1835.7000 1822.5400 ;
        RECT 1834.1000 1827.5000 1835.7000 1827.9800 ;
        RECT 1789.1000 1832.9400 1790.7000 1833.4200 ;
        RECT 1789.1000 1838.3800 1790.7000 1838.8600 ;
        RECT 1789.1000 1843.8200 1790.7000 1844.3000 ;
        RECT 1789.1000 1822.0600 1790.7000 1822.5400 ;
        RECT 1789.1000 1827.5000 1790.7000 1827.9800 ;
        RECT 1834.1000 1805.7400 1835.7000 1806.2200 ;
        RECT 1834.1000 1811.1800 1835.7000 1811.6600 ;
        RECT 1834.1000 1816.6200 1835.7000 1817.1000 ;
        RECT 1834.1000 1800.3000 1835.7000 1800.7800 ;
        RECT 1789.1000 1805.7400 1790.7000 1806.2200 ;
        RECT 1789.1000 1811.1800 1790.7000 1811.6600 ;
        RECT 1789.1000 1816.6200 1790.7000 1817.1000 ;
        RECT 1789.1000 1800.3000 1790.7000 1800.7800 ;
        RECT 1744.1000 1832.9400 1745.7000 1833.4200 ;
        RECT 1744.1000 1838.3800 1745.7000 1838.8600 ;
        RECT 1744.1000 1843.8200 1745.7000 1844.3000 ;
        RECT 1736.3400 1832.9400 1737.9400 1833.4200 ;
        RECT 1736.3400 1838.3800 1737.9400 1838.8600 ;
        RECT 1736.3400 1843.8200 1737.9400 1844.3000 ;
        RECT 1744.1000 1822.0600 1745.7000 1822.5400 ;
        RECT 1744.1000 1827.5000 1745.7000 1827.9800 ;
        RECT 1736.3400 1822.0600 1737.9400 1822.5400 ;
        RECT 1736.3400 1827.5000 1737.9400 1827.9800 ;
        RECT 1744.1000 1805.7400 1745.7000 1806.2200 ;
        RECT 1744.1000 1811.1800 1745.7000 1811.6600 ;
        RECT 1744.1000 1816.6200 1745.7000 1817.1000 ;
        RECT 1736.3400 1805.7400 1737.9400 1806.2200 ;
        RECT 1736.3400 1811.1800 1737.9400 1811.6600 ;
        RECT 1736.3400 1816.6200 1737.9400 1817.1000 ;
        RECT 1736.3400 1800.3000 1737.9400 1800.7800 ;
        RECT 1744.1000 1800.3000 1745.7000 1800.7800 ;
        RECT 1730.7800 2002.6100 1941.0000 2004.2100 ;
        RECT 1730.7800 1796.1100 1941.0000 1797.7100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1790.6800 1737.9400 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 2008.7200 1737.9400 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1790.6800 1935.4400 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 2008.7200 1935.4400 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1796.1100 1732.3800 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1796.1100 1941.0000 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 2002.6100 1732.3800 2004.2100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 2002.6100 1941.0000 2004.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 1566.4700 1925.7000 1774.5700 ;
        RECT 1879.1000 1566.4700 1880.7000 1774.5700 ;
        RECT 1834.1000 1566.4700 1835.7000 1774.5700 ;
        RECT 1789.1000 1566.4700 1790.7000 1774.5700 ;
        RECT 1744.1000 1566.4700 1745.7000 1774.5700 ;
        RECT 1933.8400 1561.0400 1935.4400 1780.6800 ;
        RECT 1736.3400 1561.0400 1737.9400 1780.6800 ;
      LAYER met3 ;
        RECT 1933.8400 1755.6200 1935.4400 1756.1000 ;
        RECT 1933.8400 1761.0600 1935.4400 1761.5400 ;
        RECT 1924.1000 1755.6200 1925.7000 1756.1000 ;
        RECT 1924.1000 1761.0600 1925.7000 1761.5400 ;
        RECT 1924.1000 1766.5000 1925.7000 1766.9800 ;
        RECT 1933.8400 1766.5000 1935.4400 1766.9800 ;
        RECT 1933.8400 1744.7400 1935.4400 1745.2200 ;
        RECT 1933.8400 1750.1800 1935.4400 1750.6600 ;
        RECT 1924.1000 1744.7400 1925.7000 1745.2200 ;
        RECT 1924.1000 1750.1800 1925.7000 1750.6600 ;
        RECT 1933.8400 1728.4200 1935.4400 1728.9000 ;
        RECT 1933.8400 1733.8600 1935.4400 1734.3400 ;
        RECT 1924.1000 1728.4200 1925.7000 1728.9000 ;
        RECT 1924.1000 1733.8600 1925.7000 1734.3400 ;
        RECT 1924.1000 1739.3000 1925.7000 1739.7800 ;
        RECT 1933.8400 1739.3000 1935.4400 1739.7800 ;
        RECT 1879.1000 1755.6200 1880.7000 1756.1000 ;
        RECT 1879.1000 1761.0600 1880.7000 1761.5400 ;
        RECT 1879.1000 1766.5000 1880.7000 1766.9800 ;
        RECT 1879.1000 1744.7400 1880.7000 1745.2200 ;
        RECT 1879.1000 1750.1800 1880.7000 1750.6600 ;
        RECT 1879.1000 1728.4200 1880.7000 1728.9000 ;
        RECT 1879.1000 1733.8600 1880.7000 1734.3400 ;
        RECT 1879.1000 1739.3000 1880.7000 1739.7800 ;
        RECT 1933.8400 1712.1000 1935.4400 1712.5800 ;
        RECT 1933.8400 1717.5400 1935.4400 1718.0200 ;
        RECT 1933.8400 1722.9800 1935.4400 1723.4600 ;
        RECT 1924.1000 1712.1000 1925.7000 1712.5800 ;
        RECT 1924.1000 1717.5400 1925.7000 1718.0200 ;
        RECT 1924.1000 1722.9800 1925.7000 1723.4600 ;
        RECT 1933.8400 1701.2200 1935.4400 1701.7000 ;
        RECT 1933.8400 1706.6600 1935.4400 1707.1400 ;
        RECT 1924.1000 1701.2200 1925.7000 1701.7000 ;
        RECT 1924.1000 1706.6600 1925.7000 1707.1400 ;
        RECT 1933.8400 1684.9000 1935.4400 1685.3800 ;
        RECT 1933.8400 1690.3400 1935.4400 1690.8200 ;
        RECT 1933.8400 1695.7800 1935.4400 1696.2600 ;
        RECT 1924.1000 1684.9000 1925.7000 1685.3800 ;
        RECT 1924.1000 1690.3400 1925.7000 1690.8200 ;
        RECT 1924.1000 1695.7800 1925.7000 1696.2600 ;
        RECT 1933.8400 1674.0200 1935.4400 1674.5000 ;
        RECT 1933.8400 1679.4600 1935.4400 1679.9400 ;
        RECT 1924.1000 1674.0200 1925.7000 1674.5000 ;
        RECT 1924.1000 1679.4600 1925.7000 1679.9400 ;
        RECT 1879.1000 1712.1000 1880.7000 1712.5800 ;
        RECT 1879.1000 1717.5400 1880.7000 1718.0200 ;
        RECT 1879.1000 1722.9800 1880.7000 1723.4600 ;
        RECT 1879.1000 1701.2200 1880.7000 1701.7000 ;
        RECT 1879.1000 1706.6600 1880.7000 1707.1400 ;
        RECT 1879.1000 1684.9000 1880.7000 1685.3800 ;
        RECT 1879.1000 1690.3400 1880.7000 1690.8200 ;
        RECT 1879.1000 1695.7800 1880.7000 1696.2600 ;
        RECT 1879.1000 1674.0200 1880.7000 1674.5000 ;
        RECT 1879.1000 1679.4600 1880.7000 1679.9400 ;
        RECT 1834.1000 1755.6200 1835.7000 1756.1000 ;
        RECT 1834.1000 1761.0600 1835.7000 1761.5400 ;
        RECT 1834.1000 1766.5000 1835.7000 1766.9800 ;
        RECT 1789.1000 1755.6200 1790.7000 1756.1000 ;
        RECT 1789.1000 1761.0600 1790.7000 1761.5400 ;
        RECT 1789.1000 1766.5000 1790.7000 1766.9800 ;
        RECT 1834.1000 1744.7400 1835.7000 1745.2200 ;
        RECT 1834.1000 1750.1800 1835.7000 1750.6600 ;
        RECT 1834.1000 1728.4200 1835.7000 1728.9000 ;
        RECT 1834.1000 1733.8600 1835.7000 1734.3400 ;
        RECT 1834.1000 1739.3000 1835.7000 1739.7800 ;
        RECT 1789.1000 1744.7400 1790.7000 1745.2200 ;
        RECT 1789.1000 1750.1800 1790.7000 1750.6600 ;
        RECT 1789.1000 1728.4200 1790.7000 1728.9000 ;
        RECT 1789.1000 1733.8600 1790.7000 1734.3400 ;
        RECT 1789.1000 1739.3000 1790.7000 1739.7800 ;
        RECT 1744.1000 1755.6200 1745.7000 1756.1000 ;
        RECT 1744.1000 1761.0600 1745.7000 1761.5400 ;
        RECT 1736.3400 1755.6200 1737.9400 1756.1000 ;
        RECT 1736.3400 1761.0600 1737.9400 1761.5400 ;
        RECT 1736.3400 1766.5000 1737.9400 1766.9800 ;
        RECT 1744.1000 1766.5000 1745.7000 1766.9800 ;
        RECT 1744.1000 1744.7400 1745.7000 1745.2200 ;
        RECT 1744.1000 1750.1800 1745.7000 1750.6600 ;
        RECT 1736.3400 1744.7400 1737.9400 1745.2200 ;
        RECT 1736.3400 1750.1800 1737.9400 1750.6600 ;
        RECT 1744.1000 1728.4200 1745.7000 1728.9000 ;
        RECT 1744.1000 1733.8600 1745.7000 1734.3400 ;
        RECT 1736.3400 1728.4200 1737.9400 1728.9000 ;
        RECT 1736.3400 1733.8600 1737.9400 1734.3400 ;
        RECT 1736.3400 1739.3000 1737.9400 1739.7800 ;
        RECT 1744.1000 1739.3000 1745.7000 1739.7800 ;
        RECT 1834.1000 1712.1000 1835.7000 1712.5800 ;
        RECT 1834.1000 1717.5400 1835.7000 1718.0200 ;
        RECT 1834.1000 1722.9800 1835.7000 1723.4600 ;
        RECT 1834.1000 1701.2200 1835.7000 1701.7000 ;
        RECT 1834.1000 1706.6600 1835.7000 1707.1400 ;
        RECT 1789.1000 1712.1000 1790.7000 1712.5800 ;
        RECT 1789.1000 1717.5400 1790.7000 1718.0200 ;
        RECT 1789.1000 1722.9800 1790.7000 1723.4600 ;
        RECT 1789.1000 1701.2200 1790.7000 1701.7000 ;
        RECT 1789.1000 1706.6600 1790.7000 1707.1400 ;
        RECT 1834.1000 1684.9000 1835.7000 1685.3800 ;
        RECT 1834.1000 1690.3400 1835.7000 1690.8200 ;
        RECT 1834.1000 1695.7800 1835.7000 1696.2600 ;
        RECT 1834.1000 1674.0200 1835.7000 1674.5000 ;
        RECT 1834.1000 1679.4600 1835.7000 1679.9400 ;
        RECT 1789.1000 1684.9000 1790.7000 1685.3800 ;
        RECT 1789.1000 1690.3400 1790.7000 1690.8200 ;
        RECT 1789.1000 1695.7800 1790.7000 1696.2600 ;
        RECT 1789.1000 1674.0200 1790.7000 1674.5000 ;
        RECT 1789.1000 1679.4600 1790.7000 1679.9400 ;
        RECT 1744.1000 1712.1000 1745.7000 1712.5800 ;
        RECT 1744.1000 1717.5400 1745.7000 1718.0200 ;
        RECT 1744.1000 1722.9800 1745.7000 1723.4600 ;
        RECT 1736.3400 1712.1000 1737.9400 1712.5800 ;
        RECT 1736.3400 1717.5400 1737.9400 1718.0200 ;
        RECT 1736.3400 1722.9800 1737.9400 1723.4600 ;
        RECT 1744.1000 1701.2200 1745.7000 1701.7000 ;
        RECT 1744.1000 1706.6600 1745.7000 1707.1400 ;
        RECT 1736.3400 1701.2200 1737.9400 1701.7000 ;
        RECT 1736.3400 1706.6600 1737.9400 1707.1400 ;
        RECT 1744.1000 1684.9000 1745.7000 1685.3800 ;
        RECT 1744.1000 1690.3400 1745.7000 1690.8200 ;
        RECT 1744.1000 1695.7800 1745.7000 1696.2600 ;
        RECT 1736.3400 1684.9000 1737.9400 1685.3800 ;
        RECT 1736.3400 1690.3400 1737.9400 1690.8200 ;
        RECT 1736.3400 1695.7800 1737.9400 1696.2600 ;
        RECT 1744.1000 1674.0200 1745.7000 1674.5000 ;
        RECT 1744.1000 1679.4600 1745.7000 1679.9400 ;
        RECT 1736.3400 1674.0200 1737.9400 1674.5000 ;
        RECT 1736.3400 1679.4600 1737.9400 1679.9400 ;
        RECT 1933.8400 1657.7000 1935.4400 1658.1800 ;
        RECT 1933.8400 1663.1400 1935.4400 1663.6200 ;
        RECT 1933.8400 1668.5800 1935.4400 1669.0600 ;
        RECT 1924.1000 1657.7000 1925.7000 1658.1800 ;
        RECT 1924.1000 1663.1400 1925.7000 1663.6200 ;
        RECT 1924.1000 1668.5800 1925.7000 1669.0600 ;
        RECT 1933.8400 1646.8200 1935.4400 1647.3000 ;
        RECT 1933.8400 1652.2600 1935.4400 1652.7400 ;
        RECT 1924.1000 1646.8200 1925.7000 1647.3000 ;
        RECT 1924.1000 1652.2600 1925.7000 1652.7400 ;
        RECT 1933.8400 1630.5000 1935.4400 1630.9800 ;
        RECT 1933.8400 1635.9400 1935.4400 1636.4200 ;
        RECT 1933.8400 1641.3800 1935.4400 1641.8600 ;
        RECT 1924.1000 1630.5000 1925.7000 1630.9800 ;
        RECT 1924.1000 1635.9400 1925.7000 1636.4200 ;
        RECT 1924.1000 1641.3800 1925.7000 1641.8600 ;
        RECT 1933.8400 1619.6200 1935.4400 1620.1000 ;
        RECT 1933.8400 1625.0600 1935.4400 1625.5400 ;
        RECT 1924.1000 1619.6200 1925.7000 1620.1000 ;
        RECT 1924.1000 1625.0600 1925.7000 1625.5400 ;
        RECT 1879.1000 1657.7000 1880.7000 1658.1800 ;
        RECT 1879.1000 1663.1400 1880.7000 1663.6200 ;
        RECT 1879.1000 1668.5800 1880.7000 1669.0600 ;
        RECT 1879.1000 1646.8200 1880.7000 1647.3000 ;
        RECT 1879.1000 1652.2600 1880.7000 1652.7400 ;
        RECT 1879.1000 1630.5000 1880.7000 1630.9800 ;
        RECT 1879.1000 1635.9400 1880.7000 1636.4200 ;
        RECT 1879.1000 1641.3800 1880.7000 1641.8600 ;
        RECT 1879.1000 1619.6200 1880.7000 1620.1000 ;
        RECT 1879.1000 1625.0600 1880.7000 1625.5400 ;
        RECT 1933.8400 1603.3000 1935.4400 1603.7800 ;
        RECT 1933.8400 1608.7400 1935.4400 1609.2200 ;
        RECT 1933.8400 1614.1800 1935.4400 1614.6600 ;
        RECT 1924.1000 1603.3000 1925.7000 1603.7800 ;
        RECT 1924.1000 1608.7400 1925.7000 1609.2200 ;
        RECT 1924.1000 1614.1800 1925.7000 1614.6600 ;
        RECT 1933.8400 1592.4200 1935.4400 1592.9000 ;
        RECT 1933.8400 1597.8600 1935.4400 1598.3400 ;
        RECT 1924.1000 1592.4200 1925.7000 1592.9000 ;
        RECT 1924.1000 1597.8600 1925.7000 1598.3400 ;
        RECT 1933.8400 1576.1000 1935.4400 1576.5800 ;
        RECT 1933.8400 1581.5400 1935.4400 1582.0200 ;
        RECT 1933.8400 1586.9800 1935.4400 1587.4600 ;
        RECT 1924.1000 1576.1000 1925.7000 1576.5800 ;
        RECT 1924.1000 1581.5400 1925.7000 1582.0200 ;
        RECT 1924.1000 1586.9800 1925.7000 1587.4600 ;
        RECT 1924.1000 1570.6600 1925.7000 1571.1400 ;
        RECT 1933.8400 1570.6600 1935.4400 1571.1400 ;
        RECT 1879.1000 1603.3000 1880.7000 1603.7800 ;
        RECT 1879.1000 1608.7400 1880.7000 1609.2200 ;
        RECT 1879.1000 1614.1800 1880.7000 1614.6600 ;
        RECT 1879.1000 1592.4200 1880.7000 1592.9000 ;
        RECT 1879.1000 1597.8600 1880.7000 1598.3400 ;
        RECT 1879.1000 1576.1000 1880.7000 1576.5800 ;
        RECT 1879.1000 1581.5400 1880.7000 1582.0200 ;
        RECT 1879.1000 1586.9800 1880.7000 1587.4600 ;
        RECT 1879.1000 1570.6600 1880.7000 1571.1400 ;
        RECT 1834.1000 1657.7000 1835.7000 1658.1800 ;
        RECT 1834.1000 1663.1400 1835.7000 1663.6200 ;
        RECT 1834.1000 1668.5800 1835.7000 1669.0600 ;
        RECT 1834.1000 1646.8200 1835.7000 1647.3000 ;
        RECT 1834.1000 1652.2600 1835.7000 1652.7400 ;
        RECT 1789.1000 1657.7000 1790.7000 1658.1800 ;
        RECT 1789.1000 1663.1400 1790.7000 1663.6200 ;
        RECT 1789.1000 1668.5800 1790.7000 1669.0600 ;
        RECT 1789.1000 1646.8200 1790.7000 1647.3000 ;
        RECT 1789.1000 1652.2600 1790.7000 1652.7400 ;
        RECT 1834.1000 1630.5000 1835.7000 1630.9800 ;
        RECT 1834.1000 1635.9400 1835.7000 1636.4200 ;
        RECT 1834.1000 1641.3800 1835.7000 1641.8600 ;
        RECT 1834.1000 1619.6200 1835.7000 1620.1000 ;
        RECT 1834.1000 1625.0600 1835.7000 1625.5400 ;
        RECT 1789.1000 1630.5000 1790.7000 1630.9800 ;
        RECT 1789.1000 1635.9400 1790.7000 1636.4200 ;
        RECT 1789.1000 1641.3800 1790.7000 1641.8600 ;
        RECT 1789.1000 1619.6200 1790.7000 1620.1000 ;
        RECT 1789.1000 1625.0600 1790.7000 1625.5400 ;
        RECT 1744.1000 1657.7000 1745.7000 1658.1800 ;
        RECT 1744.1000 1663.1400 1745.7000 1663.6200 ;
        RECT 1744.1000 1668.5800 1745.7000 1669.0600 ;
        RECT 1736.3400 1657.7000 1737.9400 1658.1800 ;
        RECT 1736.3400 1663.1400 1737.9400 1663.6200 ;
        RECT 1736.3400 1668.5800 1737.9400 1669.0600 ;
        RECT 1744.1000 1646.8200 1745.7000 1647.3000 ;
        RECT 1744.1000 1652.2600 1745.7000 1652.7400 ;
        RECT 1736.3400 1646.8200 1737.9400 1647.3000 ;
        RECT 1736.3400 1652.2600 1737.9400 1652.7400 ;
        RECT 1744.1000 1630.5000 1745.7000 1630.9800 ;
        RECT 1744.1000 1635.9400 1745.7000 1636.4200 ;
        RECT 1744.1000 1641.3800 1745.7000 1641.8600 ;
        RECT 1736.3400 1630.5000 1737.9400 1630.9800 ;
        RECT 1736.3400 1635.9400 1737.9400 1636.4200 ;
        RECT 1736.3400 1641.3800 1737.9400 1641.8600 ;
        RECT 1744.1000 1619.6200 1745.7000 1620.1000 ;
        RECT 1744.1000 1625.0600 1745.7000 1625.5400 ;
        RECT 1736.3400 1619.6200 1737.9400 1620.1000 ;
        RECT 1736.3400 1625.0600 1737.9400 1625.5400 ;
        RECT 1834.1000 1603.3000 1835.7000 1603.7800 ;
        RECT 1834.1000 1608.7400 1835.7000 1609.2200 ;
        RECT 1834.1000 1614.1800 1835.7000 1614.6600 ;
        RECT 1834.1000 1592.4200 1835.7000 1592.9000 ;
        RECT 1834.1000 1597.8600 1835.7000 1598.3400 ;
        RECT 1789.1000 1603.3000 1790.7000 1603.7800 ;
        RECT 1789.1000 1608.7400 1790.7000 1609.2200 ;
        RECT 1789.1000 1614.1800 1790.7000 1614.6600 ;
        RECT 1789.1000 1592.4200 1790.7000 1592.9000 ;
        RECT 1789.1000 1597.8600 1790.7000 1598.3400 ;
        RECT 1834.1000 1576.1000 1835.7000 1576.5800 ;
        RECT 1834.1000 1581.5400 1835.7000 1582.0200 ;
        RECT 1834.1000 1586.9800 1835.7000 1587.4600 ;
        RECT 1834.1000 1570.6600 1835.7000 1571.1400 ;
        RECT 1789.1000 1576.1000 1790.7000 1576.5800 ;
        RECT 1789.1000 1581.5400 1790.7000 1582.0200 ;
        RECT 1789.1000 1586.9800 1790.7000 1587.4600 ;
        RECT 1789.1000 1570.6600 1790.7000 1571.1400 ;
        RECT 1744.1000 1603.3000 1745.7000 1603.7800 ;
        RECT 1744.1000 1608.7400 1745.7000 1609.2200 ;
        RECT 1744.1000 1614.1800 1745.7000 1614.6600 ;
        RECT 1736.3400 1603.3000 1737.9400 1603.7800 ;
        RECT 1736.3400 1608.7400 1737.9400 1609.2200 ;
        RECT 1736.3400 1614.1800 1737.9400 1614.6600 ;
        RECT 1744.1000 1592.4200 1745.7000 1592.9000 ;
        RECT 1744.1000 1597.8600 1745.7000 1598.3400 ;
        RECT 1736.3400 1592.4200 1737.9400 1592.9000 ;
        RECT 1736.3400 1597.8600 1737.9400 1598.3400 ;
        RECT 1744.1000 1576.1000 1745.7000 1576.5800 ;
        RECT 1744.1000 1581.5400 1745.7000 1582.0200 ;
        RECT 1744.1000 1586.9800 1745.7000 1587.4600 ;
        RECT 1736.3400 1576.1000 1737.9400 1576.5800 ;
        RECT 1736.3400 1581.5400 1737.9400 1582.0200 ;
        RECT 1736.3400 1586.9800 1737.9400 1587.4600 ;
        RECT 1736.3400 1570.6600 1737.9400 1571.1400 ;
        RECT 1744.1000 1570.6600 1745.7000 1571.1400 ;
        RECT 1730.7800 1772.9700 1941.0000 1774.5700 ;
        RECT 1730.7800 1566.4700 1941.0000 1568.0700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1561.0400 1737.9400 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1779.0800 1737.9400 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1561.0400 1935.4400 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1779.0800 1935.4400 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1566.4700 1732.3800 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1566.4700 1941.0000 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1772.9700 1732.3800 1774.5700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1772.9700 1941.0000 1774.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 1336.8300 1925.7000 1544.9300 ;
        RECT 1879.1000 1336.8300 1880.7000 1544.9300 ;
        RECT 1834.1000 1336.8300 1835.7000 1544.9300 ;
        RECT 1789.1000 1336.8300 1790.7000 1544.9300 ;
        RECT 1744.1000 1336.8300 1745.7000 1544.9300 ;
        RECT 1933.8400 1331.4000 1935.4400 1551.0400 ;
        RECT 1736.3400 1331.4000 1737.9400 1551.0400 ;
      LAYER met3 ;
        RECT 1933.8400 1525.9800 1935.4400 1526.4600 ;
        RECT 1933.8400 1531.4200 1935.4400 1531.9000 ;
        RECT 1924.1000 1525.9800 1925.7000 1526.4600 ;
        RECT 1924.1000 1531.4200 1925.7000 1531.9000 ;
        RECT 1924.1000 1536.8600 1925.7000 1537.3400 ;
        RECT 1933.8400 1536.8600 1935.4400 1537.3400 ;
        RECT 1933.8400 1515.1000 1935.4400 1515.5800 ;
        RECT 1933.8400 1520.5400 1935.4400 1521.0200 ;
        RECT 1924.1000 1515.1000 1925.7000 1515.5800 ;
        RECT 1924.1000 1520.5400 1925.7000 1521.0200 ;
        RECT 1933.8400 1498.7800 1935.4400 1499.2600 ;
        RECT 1933.8400 1504.2200 1935.4400 1504.7000 ;
        RECT 1924.1000 1498.7800 1925.7000 1499.2600 ;
        RECT 1924.1000 1504.2200 1925.7000 1504.7000 ;
        RECT 1924.1000 1509.6600 1925.7000 1510.1400 ;
        RECT 1933.8400 1509.6600 1935.4400 1510.1400 ;
        RECT 1879.1000 1525.9800 1880.7000 1526.4600 ;
        RECT 1879.1000 1531.4200 1880.7000 1531.9000 ;
        RECT 1879.1000 1536.8600 1880.7000 1537.3400 ;
        RECT 1879.1000 1515.1000 1880.7000 1515.5800 ;
        RECT 1879.1000 1520.5400 1880.7000 1521.0200 ;
        RECT 1879.1000 1498.7800 1880.7000 1499.2600 ;
        RECT 1879.1000 1504.2200 1880.7000 1504.7000 ;
        RECT 1879.1000 1509.6600 1880.7000 1510.1400 ;
        RECT 1933.8400 1482.4600 1935.4400 1482.9400 ;
        RECT 1933.8400 1487.9000 1935.4400 1488.3800 ;
        RECT 1933.8400 1493.3400 1935.4400 1493.8200 ;
        RECT 1924.1000 1482.4600 1925.7000 1482.9400 ;
        RECT 1924.1000 1487.9000 1925.7000 1488.3800 ;
        RECT 1924.1000 1493.3400 1925.7000 1493.8200 ;
        RECT 1933.8400 1471.5800 1935.4400 1472.0600 ;
        RECT 1933.8400 1477.0200 1935.4400 1477.5000 ;
        RECT 1924.1000 1471.5800 1925.7000 1472.0600 ;
        RECT 1924.1000 1477.0200 1925.7000 1477.5000 ;
        RECT 1933.8400 1455.2600 1935.4400 1455.7400 ;
        RECT 1933.8400 1460.7000 1935.4400 1461.1800 ;
        RECT 1933.8400 1466.1400 1935.4400 1466.6200 ;
        RECT 1924.1000 1455.2600 1925.7000 1455.7400 ;
        RECT 1924.1000 1460.7000 1925.7000 1461.1800 ;
        RECT 1924.1000 1466.1400 1925.7000 1466.6200 ;
        RECT 1933.8400 1444.3800 1935.4400 1444.8600 ;
        RECT 1933.8400 1449.8200 1935.4400 1450.3000 ;
        RECT 1924.1000 1444.3800 1925.7000 1444.8600 ;
        RECT 1924.1000 1449.8200 1925.7000 1450.3000 ;
        RECT 1879.1000 1482.4600 1880.7000 1482.9400 ;
        RECT 1879.1000 1487.9000 1880.7000 1488.3800 ;
        RECT 1879.1000 1493.3400 1880.7000 1493.8200 ;
        RECT 1879.1000 1471.5800 1880.7000 1472.0600 ;
        RECT 1879.1000 1477.0200 1880.7000 1477.5000 ;
        RECT 1879.1000 1455.2600 1880.7000 1455.7400 ;
        RECT 1879.1000 1460.7000 1880.7000 1461.1800 ;
        RECT 1879.1000 1466.1400 1880.7000 1466.6200 ;
        RECT 1879.1000 1444.3800 1880.7000 1444.8600 ;
        RECT 1879.1000 1449.8200 1880.7000 1450.3000 ;
        RECT 1834.1000 1525.9800 1835.7000 1526.4600 ;
        RECT 1834.1000 1531.4200 1835.7000 1531.9000 ;
        RECT 1834.1000 1536.8600 1835.7000 1537.3400 ;
        RECT 1789.1000 1525.9800 1790.7000 1526.4600 ;
        RECT 1789.1000 1531.4200 1790.7000 1531.9000 ;
        RECT 1789.1000 1536.8600 1790.7000 1537.3400 ;
        RECT 1834.1000 1515.1000 1835.7000 1515.5800 ;
        RECT 1834.1000 1520.5400 1835.7000 1521.0200 ;
        RECT 1834.1000 1498.7800 1835.7000 1499.2600 ;
        RECT 1834.1000 1504.2200 1835.7000 1504.7000 ;
        RECT 1834.1000 1509.6600 1835.7000 1510.1400 ;
        RECT 1789.1000 1515.1000 1790.7000 1515.5800 ;
        RECT 1789.1000 1520.5400 1790.7000 1521.0200 ;
        RECT 1789.1000 1498.7800 1790.7000 1499.2600 ;
        RECT 1789.1000 1504.2200 1790.7000 1504.7000 ;
        RECT 1789.1000 1509.6600 1790.7000 1510.1400 ;
        RECT 1744.1000 1525.9800 1745.7000 1526.4600 ;
        RECT 1744.1000 1531.4200 1745.7000 1531.9000 ;
        RECT 1736.3400 1525.9800 1737.9400 1526.4600 ;
        RECT 1736.3400 1531.4200 1737.9400 1531.9000 ;
        RECT 1736.3400 1536.8600 1737.9400 1537.3400 ;
        RECT 1744.1000 1536.8600 1745.7000 1537.3400 ;
        RECT 1744.1000 1515.1000 1745.7000 1515.5800 ;
        RECT 1744.1000 1520.5400 1745.7000 1521.0200 ;
        RECT 1736.3400 1515.1000 1737.9400 1515.5800 ;
        RECT 1736.3400 1520.5400 1737.9400 1521.0200 ;
        RECT 1744.1000 1498.7800 1745.7000 1499.2600 ;
        RECT 1744.1000 1504.2200 1745.7000 1504.7000 ;
        RECT 1736.3400 1498.7800 1737.9400 1499.2600 ;
        RECT 1736.3400 1504.2200 1737.9400 1504.7000 ;
        RECT 1736.3400 1509.6600 1737.9400 1510.1400 ;
        RECT 1744.1000 1509.6600 1745.7000 1510.1400 ;
        RECT 1834.1000 1482.4600 1835.7000 1482.9400 ;
        RECT 1834.1000 1487.9000 1835.7000 1488.3800 ;
        RECT 1834.1000 1493.3400 1835.7000 1493.8200 ;
        RECT 1834.1000 1471.5800 1835.7000 1472.0600 ;
        RECT 1834.1000 1477.0200 1835.7000 1477.5000 ;
        RECT 1789.1000 1482.4600 1790.7000 1482.9400 ;
        RECT 1789.1000 1487.9000 1790.7000 1488.3800 ;
        RECT 1789.1000 1493.3400 1790.7000 1493.8200 ;
        RECT 1789.1000 1471.5800 1790.7000 1472.0600 ;
        RECT 1789.1000 1477.0200 1790.7000 1477.5000 ;
        RECT 1834.1000 1455.2600 1835.7000 1455.7400 ;
        RECT 1834.1000 1460.7000 1835.7000 1461.1800 ;
        RECT 1834.1000 1466.1400 1835.7000 1466.6200 ;
        RECT 1834.1000 1444.3800 1835.7000 1444.8600 ;
        RECT 1834.1000 1449.8200 1835.7000 1450.3000 ;
        RECT 1789.1000 1455.2600 1790.7000 1455.7400 ;
        RECT 1789.1000 1460.7000 1790.7000 1461.1800 ;
        RECT 1789.1000 1466.1400 1790.7000 1466.6200 ;
        RECT 1789.1000 1444.3800 1790.7000 1444.8600 ;
        RECT 1789.1000 1449.8200 1790.7000 1450.3000 ;
        RECT 1744.1000 1482.4600 1745.7000 1482.9400 ;
        RECT 1744.1000 1487.9000 1745.7000 1488.3800 ;
        RECT 1744.1000 1493.3400 1745.7000 1493.8200 ;
        RECT 1736.3400 1482.4600 1737.9400 1482.9400 ;
        RECT 1736.3400 1487.9000 1737.9400 1488.3800 ;
        RECT 1736.3400 1493.3400 1737.9400 1493.8200 ;
        RECT 1744.1000 1471.5800 1745.7000 1472.0600 ;
        RECT 1744.1000 1477.0200 1745.7000 1477.5000 ;
        RECT 1736.3400 1471.5800 1737.9400 1472.0600 ;
        RECT 1736.3400 1477.0200 1737.9400 1477.5000 ;
        RECT 1744.1000 1455.2600 1745.7000 1455.7400 ;
        RECT 1744.1000 1460.7000 1745.7000 1461.1800 ;
        RECT 1744.1000 1466.1400 1745.7000 1466.6200 ;
        RECT 1736.3400 1455.2600 1737.9400 1455.7400 ;
        RECT 1736.3400 1460.7000 1737.9400 1461.1800 ;
        RECT 1736.3400 1466.1400 1737.9400 1466.6200 ;
        RECT 1744.1000 1444.3800 1745.7000 1444.8600 ;
        RECT 1744.1000 1449.8200 1745.7000 1450.3000 ;
        RECT 1736.3400 1444.3800 1737.9400 1444.8600 ;
        RECT 1736.3400 1449.8200 1737.9400 1450.3000 ;
        RECT 1933.8400 1428.0600 1935.4400 1428.5400 ;
        RECT 1933.8400 1433.5000 1935.4400 1433.9800 ;
        RECT 1933.8400 1438.9400 1935.4400 1439.4200 ;
        RECT 1924.1000 1428.0600 1925.7000 1428.5400 ;
        RECT 1924.1000 1433.5000 1925.7000 1433.9800 ;
        RECT 1924.1000 1438.9400 1925.7000 1439.4200 ;
        RECT 1933.8400 1417.1800 1935.4400 1417.6600 ;
        RECT 1933.8400 1422.6200 1935.4400 1423.1000 ;
        RECT 1924.1000 1417.1800 1925.7000 1417.6600 ;
        RECT 1924.1000 1422.6200 1925.7000 1423.1000 ;
        RECT 1933.8400 1400.8600 1935.4400 1401.3400 ;
        RECT 1933.8400 1406.3000 1935.4400 1406.7800 ;
        RECT 1933.8400 1411.7400 1935.4400 1412.2200 ;
        RECT 1924.1000 1400.8600 1925.7000 1401.3400 ;
        RECT 1924.1000 1406.3000 1925.7000 1406.7800 ;
        RECT 1924.1000 1411.7400 1925.7000 1412.2200 ;
        RECT 1933.8400 1389.9800 1935.4400 1390.4600 ;
        RECT 1933.8400 1395.4200 1935.4400 1395.9000 ;
        RECT 1924.1000 1389.9800 1925.7000 1390.4600 ;
        RECT 1924.1000 1395.4200 1925.7000 1395.9000 ;
        RECT 1879.1000 1428.0600 1880.7000 1428.5400 ;
        RECT 1879.1000 1433.5000 1880.7000 1433.9800 ;
        RECT 1879.1000 1438.9400 1880.7000 1439.4200 ;
        RECT 1879.1000 1417.1800 1880.7000 1417.6600 ;
        RECT 1879.1000 1422.6200 1880.7000 1423.1000 ;
        RECT 1879.1000 1400.8600 1880.7000 1401.3400 ;
        RECT 1879.1000 1406.3000 1880.7000 1406.7800 ;
        RECT 1879.1000 1411.7400 1880.7000 1412.2200 ;
        RECT 1879.1000 1389.9800 1880.7000 1390.4600 ;
        RECT 1879.1000 1395.4200 1880.7000 1395.9000 ;
        RECT 1933.8400 1373.6600 1935.4400 1374.1400 ;
        RECT 1933.8400 1379.1000 1935.4400 1379.5800 ;
        RECT 1933.8400 1384.5400 1935.4400 1385.0200 ;
        RECT 1924.1000 1373.6600 1925.7000 1374.1400 ;
        RECT 1924.1000 1379.1000 1925.7000 1379.5800 ;
        RECT 1924.1000 1384.5400 1925.7000 1385.0200 ;
        RECT 1933.8400 1362.7800 1935.4400 1363.2600 ;
        RECT 1933.8400 1368.2200 1935.4400 1368.7000 ;
        RECT 1924.1000 1362.7800 1925.7000 1363.2600 ;
        RECT 1924.1000 1368.2200 1925.7000 1368.7000 ;
        RECT 1933.8400 1346.4600 1935.4400 1346.9400 ;
        RECT 1933.8400 1351.9000 1935.4400 1352.3800 ;
        RECT 1933.8400 1357.3400 1935.4400 1357.8200 ;
        RECT 1924.1000 1346.4600 1925.7000 1346.9400 ;
        RECT 1924.1000 1351.9000 1925.7000 1352.3800 ;
        RECT 1924.1000 1357.3400 1925.7000 1357.8200 ;
        RECT 1924.1000 1341.0200 1925.7000 1341.5000 ;
        RECT 1933.8400 1341.0200 1935.4400 1341.5000 ;
        RECT 1879.1000 1373.6600 1880.7000 1374.1400 ;
        RECT 1879.1000 1379.1000 1880.7000 1379.5800 ;
        RECT 1879.1000 1384.5400 1880.7000 1385.0200 ;
        RECT 1879.1000 1362.7800 1880.7000 1363.2600 ;
        RECT 1879.1000 1368.2200 1880.7000 1368.7000 ;
        RECT 1879.1000 1346.4600 1880.7000 1346.9400 ;
        RECT 1879.1000 1351.9000 1880.7000 1352.3800 ;
        RECT 1879.1000 1357.3400 1880.7000 1357.8200 ;
        RECT 1879.1000 1341.0200 1880.7000 1341.5000 ;
        RECT 1834.1000 1428.0600 1835.7000 1428.5400 ;
        RECT 1834.1000 1433.5000 1835.7000 1433.9800 ;
        RECT 1834.1000 1438.9400 1835.7000 1439.4200 ;
        RECT 1834.1000 1417.1800 1835.7000 1417.6600 ;
        RECT 1834.1000 1422.6200 1835.7000 1423.1000 ;
        RECT 1789.1000 1428.0600 1790.7000 1428.5400 ;
        RECT 1789.1000 1433.5000 1790.7000 1433.9800 ;
        RECT 1789.1000 1438.9400 1790.7000 1439.4200 ;
        RECT 1789.1000 1417.1800 1790.7000 1417.6600 ;
        RECT 1789.1000 1422.6200 1790.7000 1423.1000 ;
        RECT 1834.1000 1400.8600 1835.7000 1401.3400 ;
        RECT 1834.1000 1406.3000 1835.7000 1406.7800 ;
        RECT 1834.1000 1411.7400 1835.7000 1412.2200 ;
        RECT 1834.1000 1389.9800 1835.7000 1390.4600 ;
        RECT 1834.1000 1395.4200 1835.7000 1395.9000 ;
        RECT 1789.1000 1400.8600 1790.7000 1401.3400 ;
        RECT 1789.1000 1406.3000 1790.7000 1406.7800 ;
        RECT 1789.1000 1411.7400 1790.7000 1412.2200 ;
        RECT 1789.1000 1389.9800 1790.7000 1390.4600 ;
        RECT 1789.1000 1395.4200 1790.7000 1395.9000 ;
        RECT 1744.1000 1428.0600 1745.7000 1428.5400 ;
        RECT 1744.1000 1433.5000 1745.7000 1433.9800 ;
        RECT 1744.1000 1438.9400 1745.7000 1439.4200 ;
        RECT 1736.3400 1428.0600 1737.9400 1428.5400 ;
        RECT 1736.3400 1433.5000 1737.9400 1433.9800 ;
        RECT 1736.3400 1438.9400 1737.9400 1439.4200 ;
        RECT 1744.1000 1417.1800 1745.7000 1417.6600 ;
        RECT 1744.1000 1422.6200 1745.7000 1423.1000 ;
        RECT 1736.3400 1417.1800 1737.9400 1417.6600 ;
        RECT 1736.3400 1422.6200 1737.9400 1423.1000 ;
        RECT 1744.1000 1400.8600 1745.7000 1401.3400 ;
        RECT 1744.1000 1406.3000 1745.7000 1406.7800 ;
        RECT 1744.1000 1411.7400 1745.7000 1412.2200 ;
        RECT 1736.3400 1400.8600 1737.9400 1401.3400 ;
        RECT 1736.3400 1406.3000 1737.9400 1406.7800 ;
        RECT 1736.3400 1411.7400 1737.9400 1412.2200 ;
        RECT 1744.1000 1389.9800 1745.7000 1390.4600 ;
        RECT 1744.1000 1395.4200 1745.7000 1395.9000 ;
        RECT 1736.3400 1389.9800 1737.9400 1390.4600 ;
        RECT 1736.3400 1395.4200 1737.9400 1395.9000 ;
        RECT 1834.1000 1373.6600 1835.7000 1374.1400 ;
        RECT 1834.1000 1379.1000 1835.7000 1379.5800 ;
        RECT 1834.1000 1384.5400 1835.7000 1385.0200 ;
        RECT 1834.1000 1362.7800 1835.7000 1363.2600 ;
        RECT 1834.1000 1368.2200 1835.7000 1368.7000 ;
        RECT 1789.1000 1373.6600 1790.7000 1374.1400 ;
        RECT 1789.1000 1379.1000 1790.7000 1379.5800 ;
        RECT 1789.1000 1384.5400 1790.7000 1385.0200 ;
        RECT 1789.1000 1362.7800 1790.7000 1363.2600 ;
        RECT 1789.1000 1368.2200 1790.7000 1368.7000 ;
        RECT 1834.1000 1346.4600 1835.7000 1346.9400 ;
        RECT 1834.1000 1351.9000 1835.7000 1352.3800 ;
        RECT 1834.1000 1357.3400 1835.7000 1357.8200 ;
        RECT 1834.1000 1341.0200 1835.7000 1341.5000 ;
        RECT 1789.1000 1346.4600 1790.7000 1346.9400 ;
        RECT 1789.1000 1351.9000 1790.7000 1352.3800 ;
        RECT 1789.1000 1357.3400 1790.7000 1357.8200 ;
        RECT 1789.1000 1341.0200 1790.7000 1341.5000 ;
        RECT 1744.1000 1373.6600 1745.7000 1374.1400 ;
        RECT 1744.1000 1379.1000 1745.7000 1379.5800 ;
        RECT 1744.1000 1384.5400 1745.7000 1385.0200 ;
        RECT 1736.3400 1373.6600 1737.9400 1374.1400 ;
        RECT 1736.3400 1379.1000 1737.9400 1379.5800 ;
        RECT 1736.3400 1384.5400 1737.9400 1385.0200 ;
        RECT 1744.1000 1362.7800 1745.7000 1363.2600 ;
        RECT 1744.1000 1368.2200 1745.7000 1368.7000 ;
        RECT 1736.3400 1362.7800 1737.9400 1363.2600 ;
        RECT 1736.3400 1368.2200 1737.9400 1368.7000 ;
        RECT 1744.1000 1346.4600 1745.7000 1346.9400 ;
        RECT 1744.1000 1351.9000 1745.7000 1352.3800 ;
        RECT 1744.1000 1357.3400 1745.7000 1357.8200 ;
        RECT 1736.3400 1346.4600 1737.9400 1346.9400 ;
        RECT 1736.3400 1351.9000 1737.9400 1352.3800 ;
        RECT 1736.3400 1357.3400 1737.9400 1357.8200 ;
        RECT 1736.3400 1341.0200 1737.9400 1341.5000 ;
        RECT 1744.1000 1341.0200 1745.7000 1341.5000 ;
        RECT 1730.7800 1543.3300 1941.0000 1544.9300 ;
        RECT 1730.7800 1336.8300 1941.0000 1338.4300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1331.4000 1737.9400 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1549.4400 1737.9400 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1331.4000 1935.4400 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1549.4400 1935.4400 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1336.8300 1732.3800 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1336.8300 1941.0000 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1543.3300 1732.3800 1544.9300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1543.3300 1941.0000 1544.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 1107.1900 1925.7000 1315.2900 ;
        RECT 1879.1000 1107.1900 1880.7000 1315.2900 ;
        RECT 1834.1000 1107.1900 1835.7000 1315.2900 ;
        RECT 1789.1000 1107.1900 1790.7000 1315.2900 ;
        RECT 1744.1000 1107.1900 1745.7000 1315.2900 ;
        RECT 1933.8400 1101.7600 1935.4400 1321.4000 ;
        RECT 1736.3400 1101.7600 1737.9400 1321.4000 ;
      LAYER met3 ;
        RECT 1933.8400 1296.3400 1935.4400 1296.8200 ;
        RECT 1933.8400 1301.7800 1935.4400 1302.2600 ;
        RECT 1924.1000 1296.3400 1925.7000 1296.8200 ;
        RECT 1924.1000 1301.7800 1925.7000 1302.2600 ;
        RECT 1924.1000 1307.2200 1925.7000 1307.7000 ;
        RECT 1933.8400 1307.2200 1935.4400 1307.7000 ;
        RECT 1933.8400 1285.4600 1935.4400 1285.9400 ;
        RECT 1933.8400 1290.9000 1935.4400 1291.3800 ;
        RECT 1924.1000 1285.4600 1925.7000 1285.9400 ;
        RECT 1924.1000 1290.9000 1925.7000 1291.3800 ;
        RECT 1933.8400 1269.1400 1935.4400 1269.6200 ;
        RECT 1933.8400 1274.5800 1935.4400 1275.0600 ;
        RECT 1924.1000 1269.1400 1925.7000 1269.6200 ;
        RECT 1924.1000 1274.5800 1925.7000 1275.0600 ;
        RECT 1924.1000 1280.0200 1925.7000 1280.5000 ;
        RECT 1933.8400 1280.0200 1935.4400 1280.5000 ;
        RECT 1879.1000 1296.3400 1880.7000 1296.8200 ;
        RECT 1879.1000 1301.7800 1880.7000 1302.2600 ;
        RECT 1879.1000 1307.2200 1880.7000 1307.7000 ;
        RECT 1879.1000 1285.4600 1880.7000 1285.9400 ;
        RECT 1879.1000 1290.9000 1880.7000 1291.3800 ;
        RECT 1879.1000 1269.1400 1880.7000 1269.6200 ;
        RECT 1879.1000 1274.5800 1880.7000 1275.0600 ;
        RECT 1879.1000 1280.0200 1880.7000 1280.5000 ;
        RECT 1933.8400 1252.8200 1935.4400 1253.3000 ;
        RECT 1933.8400 1258.2600 1935.4400 1258.7400 ;
        RECT 1933.8400 1263.7000 1935.4400 1264.1800 ;
        RECT 1924.1000 1252.8200 1925.7000 1253.3000 ;
        RECT 1924.1000 1258.2600 1925.7000 1258.7400 ;
        RECT 1924.1000 1263.7000 1925.7000 1264.1800 ;
        RECT 1933.8400 1241.9400 1935.4400 1242.4200 ;
        RECT 1933.8400 1247.3800 1935.4400 1247.8600 ;
        RECT 1924.1000 1241.9400 1925.7000 1242.4200 ;
        RECT 1924.1000 1247.3800 1925.7000 1247.8600 ;
        RECT 1933.8400 1225.6200 1935.4400 1226.1000 ;
        RECT 1933.8400 1231.0600 1935.4400 1231.5400 ;
        RECT 1933.8400 1236.5000 1935.4400 1236.9800 ;
        RECT 1924.1000 1225.6200 1925.7000 1226.1000 ;
        RECT 1924.1000 1231.0600 1925.7000 1231.5400 ;
        RECT 1924.1000 1236.5000 1925.7000 1236.9800 ;
        RECT 1933.8400 1214.7400 1935.4400 1215.2200 ;
        RECT 1933.8400 1220.1800 1935.4400 1220.6600 ;
        RECT 1924.1000 1214.7400 1925.7000 1215.2200 ;
        RECT 1924.1000 1220.1800 1925.7000 1220.6600 ;
        RECT 1879.1000 1252.8200 1880.7000 1253.3000 ;
        RECT 1879.1000 1258.2600 1880.7000 1258.7400 ;
        RECT 1879.1000 1263.7000 1880.7000 1264.1800 ;
        RECT 1879.1000 1241.9400 1880.7000 1242.4200 ;
        RECT 1879.1000 1247.3800 1880.7000 1247.8600 ;
        RECT 1879.1000 1225.6200 1880.7000 1226.1000 ;
        RECT 1879.1000 1231.0600 1880.7000 1231.5400 ;
        RECT 1879.1000 1236.5000 1880.7000 1236.9800 ;
        RECT 1879.1000 1214.7400 1880.7000 1215.2200 ;
        RECT 1879.1000 1220.1800 1880.7000 1220.6600 ;
        RECT 1834.1000 1296.3400 1835.7000 1296.8200 ;
        RECT 1834.1000 1301.7800 1835.7000 1302.2600 ;
        RECT 1834.1000 1307.2200 1835.7000 1307.7000 ;
        RECT 1789.1000 1296.3400 1790.7000 1296.8200 ;
        RECT 1789.1000 1301.7800 1790.7000 1302.2600 ;
        RECT 1789.1000 1307.2200 1790.7000 1307.7000 ;
        RECT 1834.1000 1285.4600 1835.7000 1285.9400 ;
        RECT 1834.1000 1290.9000 1835.7000 1291.3800 ;
        RECT 1834.1000 1269.1400 1835.7000 1269.6200 ;
        RECT 1834.1000 1274.5800 1835.7000 1275.0600 ;
        RECT 1834.1000 1280.0200 1835.7000 1280.5000 ;
        RECT 1789.1000 1285.4600 1790.7000 1285.9400 ;
        RECT 1789.1000 1290.9000 1790.7000 1291.3800 ;
        RECT 1789.1000 1269.1400 1790.7000 1269.6200 ;
        RECT 1789.1000 1274.5800 1790.7000 1275.0600 ;
        RECT 1789.1000 1280.0200 1790.7000 1280.5000 ;
        RECT 1744.1000 1296.3400 1745.7000 1296.8200 ;
        RECT 1744.1000 1301.7800 1745.7000 1302.2600 ;
        RECT 1736.3400 1296.3400 1737.9400 1296.8200 ;
        RECT 1736.3400 1301.7800 1737.9400 1302.2600 ;
        RECT 1736.3400 1307.2200 1737.9400 1307.7000 ;
        RECT 1744.1000 1307.2200 1745.7000 1307.7000 ;
        RECT 1744.1000 1285.4600 1745.7000 1285.9400 ;
        RECT 1744.1000 1290.9000 1745.7000 1291.3800 ;
        RECT 1736.3400 1285.4600 1737.9400 1285.9400 ;
        RECT 1736.3400 1290.9000 1737.9400 1291.3800 ;
        RECT 1744.1000 1269.1400 1745.7000 1269.6200 ;
        RECT 1744.1000 1274.5800 1745.7000 1275.0600 ;
        RECT 1736.3400 1269.1400 1737.9400 1269.6200 ;
        RECT 1736.3400 1274.5800 1737.9400 1275.0600 ;
        RECT 1736.3400 1280.0200 1737.9400 1280.5000 ;
        RECT 1744.1000 1280.0200 1745.7000 1280.5000 ;
        RECT 1834.1000 1252.8200 1835.7000 1253.3000 ;
        RECT 1834.1000 1258.2600 1835.7000 1258.7400 ;
        RECT 1834.1000 1263.7000 1835.7000 1264.1800 ;
        RECT 1834.1000 1241.9400 1835.7000 1242.4200 ;
        RECT 1834.1000 1247.3800 1835.7000 1247.8600 ;
        RECT 1789.1000 1252.8200 1790.7000 1253.3000 ;
        RECT 1789.1000 1258.2600 1790.7000 1258.7400 ;
        RECT 1789.1000 1263.7000 1790.7000 1264.1800 ;
        RECT 1789.1000 1241.9400 1790.7000 1242.4200 ;
        RECT 1789.1000 1247.3800 1790.7000 1247.8600 ;
        RECT 1834.1000 1225.6200 1835.7000 1226.1000 ;
        RECT 1834.1000 1231.0600 1835.7000 1231.5400 ;
        RECT 1834.1000 1236.5000 1835.7000 1236.9800 ;
        RECT 1834.1000 1214.7400 1835.7000 1215.2200 ;
        RECT 1834.1000 1220.1800 1835.7000 1220.6600 ;
        RECT 1789.1000 1225.6200 1790.7000 1226.1000 ;
        RECT 1789.1000 1231.0600 1790.7000 1231.5400 ;
        RECT 1789.1000 1236.5000 1790.7000 1236.9800 ;
        RECT 1789.1000 1214.7400 1790.7000 1215.2200 ;
        RECT 1789.1000 1220.1800 1790.7000 1220.6600 ;
        RECT 1744.1000 1252.8200 1745.7000 1253.3000 ;
        RECT 1744.1000 1258.2600 1745.7000 1258.7400 ;
        RECT 1744.1000 1263.7000 1745.7000 1264.1800 ;
        RECT 1736.3400 1252.8200 1737.9400 1253.3000 ;
        RECT 1736.3400 1258.2600 1737.9400 1258.7400 ;
        RECT 1736.3400 1263.7000 1737.9400 1264.1800 ;
        RECT 1744.1000 1241.9400 1745.7000 1242.4200 ;
        RECT 1744.1000 1247.3800 1745.7000 1247.8600 ;
        RECT 1736.3400 1241.9400 1737.9400 1242.4200 ;
        RECT 1736.3400 1247.3800 1737.9400 1247.8600 ;
        RECT 1744.1000 1225.6200 1745.7000 1226.1000 ;
        RECT 1744.1000 1231.0600 1745.7000 1231.5400 ;
        RECT 1744.1000 1236.5000 1745.7000 1236.9800 ;
        RECT 1736.3400 1225.6200 1737.9400 1226.1000 ;
        RECT 1736.3400 1231.0600 1737.9400 1231.5400 ;
        RECT 1736.3400 1236.5000 1737.9400 1236.9800 ;
        RECT 1744.1000 1214.7400 1745.7000 1215.2200 ;
        RECT 1744.1000 1220.1800 1745.7000 1220.6600 ;
        RECT 1736.3400 1214.7400 1737.9400 1215.2200 ;
        RECT 1736.3400 1220.1800 1737.9400 1220.6600 ;
        RECT 1933.8400 1198.4200 1935.4400 1198.9000 ;
        RECT 1933.8400 1203.8600 1935.4400 1204.3400 ;
        RECT 1933.8400 1209.3000 1935.4400 1209.7800 ;
        RECT 1924.1000 1198.4200 1925.7000 1198.9000 ;
        RECT 1924.1000 1203.8600 1925.7000 1204.3400 ;
        RECT 1924.1000 1209.3000 1925.7000 1209.7800 ;
        RECT 1933.8400 1187.5400 1935.4400 1188.0200 ;
        RECT 1933.8400 1192.9800 1935.4400 1193.4600 ;
        RECT 1924.1000 1187.5400 1925.7000 1188.0200 ;
        RECT 1924.1000 1192.9800 1925.7000 1193.4600 ;
        RECT 1933.8400 1171.2200 1935.4400 1171.7000 ;
        RECT 1933.8400 1176.6600 1935.4400 1177.1400 ;
        RECT 1933.8400 1182.1000 1935.4400 1182.5800 ;
        RECT 1924.1000 1171.2200 1925.7000 1171.7000 ;
        RECT 1924.1000 1176.6600 1925.7000 1177.1400 ;
        RECT 1924.1000 1182.1000 1925.7000 1182.5800 ;
        RECT 1933.8400 1160.3400 1935.4400 1160.8200 ;
        RECT 1933.8400 1165.7800 1935.4400 1166.2600 ;
        RECT 1924.1000 1160.3400 1925.7000 1160.8200 ;
        RECT 1924.1000 1165.7800 1925.7000 1166.2600 ;
        RECT 1879.1000 1198.4200 1880.7000 1198.9000 ;
        RECT 1879.1000 1203.8600 1880.7000 1204.3400 ;
        RECT 1879.1000 1209.3000 1880.7000 1209.7800 ;
        RECT 1879.1000 1187.5400 1880.7000 1188.0200 ;
        RECT 1879.1000 1192.9800 1880.7000 1193.4600 ;
        RECT 1879.1000 1171.2200 1880.7000 1171.7000 ;
        RECT 1879.1000 1176.6600 1880.7000 1177.1400 ;
        RECT 1879.1000 1182.1000 1880.7000 1182.5800 ;
        RECT 1879.1000 1160.3400 1880.7000 1160.8200 ;
        RECT 1879.1000 1165.7800 1880.7000 1166.2600 ;
        RECT 1933.8400 1144.0200 1935.4400 1144.5000 ;
        RECT 1933.8400 1149.4600 1935.4400 1149.9400 ;
        RECT 1933.8400 1154.9000 1935.4400 1155.3800 ;
        RECT 1924.1000 1144.0200 1925.7000 1144.5000 ;
        RECT 1924.1000 1149.4600 1925.7000 1149.9400 ;
        RECT 1924.1000 1154.9000 1925.7000 1155.3800 ;
        RECT 1933.8400 1133.1400 1935.4400 1133.6200 ;
        RECT 1933.8400 1138.5800 1935.4400 1139.0600 ;
        RECT 1924.1000 1133.1400 1925.7000 1133.6200 ;
        RECT 1924.1000 1138.5800 1925.7000 1139.0600 ;
        RECT 1933.8400 1116.8200 1935.4400 1117.3000 ;
        RECT 1933.8400 1122.2600 1935.4400 1122.7400 ;
        RECT 1933.8400 1127.7000 1935.4400 1128.1800 ;
        RECT 1924.1000 1116.8200 1925.7000 1117.3000 ;
        RECT 1924.1000 1122.2600 1925.7000 1122.7400 ;
        RECT 1924.1000 1127.7000 1925.7000 1128.1800 ;
        RECT 1924.1000 1111.3800 1925.7000 1111.8600 ;
        RECT 1933.8400 1111.3800 1935.4400 1111.8600 ;
        RECT 1879.1000 1144.0200 1880.7000 1144.5000 ;
        RECT 1879.1000 1149.4600 1880.7000 1149.9400 ;
        RECT 1879.1000 1154.9000 1880.7000 1155.3800 ;
        RECT 1879.1000 1133.1400 1880.7000 1133.6200 ;
        RECT 1879.1000 1138.5800 1880.7000 1139.0600 ;
        RECT 1879.1000 1116.8200 1880.7000 1117.3000 ;
        RECT 1879.1000 1122.2600 1880.7000 1122.7400 ;
        RECT 1879.1000 1127.7000 1880.7000 1128.1800 ;
        RECT 1879.1000 1111.3800 1880.7000 1111.8600 ;
        RECT 1834.1000 1198.4200 1835.7000 1198.9000 ;
        RECT 1834.1000 1203.8600 1835.7000 1204.3400 ;
        RECT 1834.1000 1209.3000 1835.7000 1209.7800 ;
        RECT 1834.1000 1187.5400 1835.7000 1188.0200 ;
        RECT 1834.1000 1192.9800 1835.7000 1193.4600 ;
        RECT 1789.1000 1198.4200 1790.7000 1198.9000 ;
        RECT 1789.1000 1203.8600 1790.7000 1204.3400 ;
        RECT 1789.1000 1209.3000 1790.7000 1209.7800 ;
        RECT 1789.1000 1187.5400 1790.7000 1188.0200 ;
        RECT 1789.1000 1192.9800 1790.7000 1193.4600 ;
        RECT 1834.1000 1171.2200 1835.7000 1171.7000 ;
        RECT 1834.1000 1176.6600 1835.7000 1177.1400 ;
        RECT 1834.1000 1182.1000 1835.7000 1182.5800 ;
        RECT 1834.1000 1160.3400 1835.7000 1160.8200 ;
        RECT 1834.1000 1165.7800 1835.7000 1166.2600 ;
        RECT 1789.1000 1171.2200 1790.7000 1171.7000 ;
        RECT 1789.1000 1176.6600 1790.7000 1177.1400 ;
        RECT 1789.1000 1182.1000 1790.7000 1182.5800 ;
        RECT 1789.1000 1160.3400 1790.7000 1160.8200 ;
        RECT 1789.1000 1165.7800 1790.7000 1166.2600 ;
        RECT 1744.1000 1198.4200 1745.7000 1198.9000 ;
        RECT 1744.1000 1203.8600 1745.7000 1204.3400 ;
        RECT 1744.1000 1209.3000 1745.7000 1209.7800 ;
        RECT 1736.3400 1198.4200 1737.9400 1198.9000 ;
        RECT 1736.3400 1203.8600 1737.9400 1204.3400 ;
        RECT 1736.3400 1209.3000 1737.9400 1209.7800 ;
        RECT 1744.1000 1187.5400 1745.7000 1188.0200 ;
        RECT 1744.1000 1192.9800 1745.7000 1193.4600 ;
        RECT 1736.3400 1187.5400 1737.9400 1188.0200 ;
        RECT 1736.3400 1192.9800 1737.9400 1193.4600 ;
        RECT 1744.1000 1171.2200 1745.7000 1171.7000 ;
        RECT 1744.1000 1176.6600 1745.7000 1177.1400 ;
        RECT 1744.1000 1182.1000 1745.7000 1182.5800 ;
        RECT 1736.3400 1171.2200 1737.9400 1171.7000 ;
        RECT 1736.3400 1176.6600 1737.9400 1177.1400 ;
        RECT 1736.3400 1182.1000 1737.9400 1182.5800 ;
        RECT 1744.1000 1160.3400 1745.7000 1160.8200 ;
        RECT 1744.1000 1165.7800 1745.7000 1166.2600 ;
        RECT 1736.3400 1160.3400 1737.9400 1160.8200 ;
        RECT 1736.3400 1165.7800 1737.9400 1166.2600 ;
        RECT 1834.1000 1144.0200 1835.7000 1144.5000 ;
        RECT 1834.1000 1149.4600 1835.7000 1149.9400 ;
        RECT 1834.1000 1154.9000 1835.7000 1155.3800 ;
        RECT 1834.1000 1133.1400 1835.7000 1133.6200 ;
        RECT 1834.1000 1138.5800 1835.7000 1139.0600 ;
        RECT 1789.1000 1144.0200 1790.7000 1144.5000 ;
        RECT 1789.1000 1149.4600 1790.7000 1149.9400 ;
        RECT 1789.1000 1154.9000 1790.7000 1155.3800 ;
        RECT 1789.1000 1133.1400 1790.7000 1133.6200 ;
        RECT 1789.1000 1138.5800 1790.7000 1139.0600 ;
        RECT 1834.1000 1116.8200 1835.7000 1117.3000 ;
        RECT 1834.1000 1122.2600 1835.7000 1122.7400 ;
        RECT 1834.1000 1127.7000 1835.7000 1128.1800 ;
        RECT 1834.1000 1111.3800 1835.7000 1111.8600 ;
        RECT 1789.1000 1116.8200 1790.7000 1117.3000 ;
        RECT 1789.1000 1122.2600 1790.7000 1122.7400 ;
        RECT 1789.1000 1127.7000 1790.7000 1128.1800 ;
        RECT 1789.1000 1111.3800 1790.7000 1111.8600 ;
        RECT 1744.1000 1144.0200 1745.7000 1144.5000 ;
        RECT 1744.1000 1149.4600 1745.7000 1149.9400 ;
        RECT 1744.1000 1154.9000 1745.7000 1155.3800 ;
        RECT 1736.3400 1144.0200 1737.9400 1144.5000 ;
        RECT 1736.3400 1149.4600 1737.9400 1149.9400 ;
        RECT 1736.3400 1154.9000 1737.9400 1155.3800 ;
        RECT 1744.1000 1133.1400 1745.7000 1133.6200 ;
        RECT 1744.1000 1138.5800 1745.7000 1139.0600 ;
        RECT 1736.3400 1133.1400 1737.9400 1133.6200 ;
        RECT 1736.3400 1138.5800 1737.9400 1139.0600 ;
        RECT 1744.1000 1116.8200 1745.7000 1117.3000 ;
        RECT 1744.1000 1122.2600 1745.7000 1122.7400 ;
        RECT 1744.1000 1127.7000 1745.7000 1128.1800 ;
        RECT 1736.3400 1116.8200 1737.9400 1117.3000 ;
        RECT 1736.3400 1122.2600 1737.9400 1122.7400 ;
        RECT 1736.3400 1127.7000 1737.9400 1128.1800 ;
        RECT 1736.3400 1111.3800 1737.9400 1111.8600 ;
        RECT 1744.1000 1111.3800 1745.7000 1111.8600 ;
        RECT 1730.7800 1313.6900 1941.0000 1315.2900 ;
        RECT 1730.7800 1107.1900 1941.0000 1108.7900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1101.7600 1737.9400 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1319.8000 1737.9400 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1101.7600 1935.4400 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1319.8000 1935.4400 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1107.1900 1732.3800 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1107.1900 1941.0000 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1313.6900 1732.3800 1315.2900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1313.6900 1941.0000 1315.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 877.5500 1925.7000 1085.6500 ;
        RECT 1879.1000 877.5500 1880.7000 1085.6500 ;
        RECT 1834.1000 877.5500 1835.7000 1085.6500 ;
        RECT 1789.1000 877.5500 1790.7000 1085.6500 ;
        RECT 1744.1000 877.5500 1745.7000 1085.6500 ;
        RECT 1933.8400 872.1200 1935.4400 1091.7600 ;
        RECT 1736.3400 872.1200 1737.9400 1091.7600 ;
      LAYER met3 ;
        RECT 1933.8400 1066.7000 1935.4400 1067.1800 ;
        RECT 1933.8400 1072.1400 1935.4400 1072.6200 ;
        RECT 1924.1000 1066.7000 1925.7000 1067.1800 ;
        RECT 1924.1000 1072.1400 1925.7000 1072.6200 ;
        RECT 1924.1000 1077.5800 1925.7000 1078.0600 ;
        RECT 1933.8400 1077.5800 1935.4400 1078.0600 ;
        RECT 1933.8400 1055.8200 1935.4400 1056.3000 ;
        RECT 1933.8400 1061.2600 1935.4400 1061.7400 ;
        RECT 1924.1000 1055.8200 1925.7000 1056.3000 ;
        RECT 1924.1000 1061.2600 1925.7000 1061.7400 ;
        RECT 1933.8400 1039.5000 1935.4400 1039.9800 ;
        RECT 1933.8400 1044.9400 1935.4400 1045.4200 ;
        RECT 1924.1000 1039.5000 1925.7000 1039.9800 ;
        RECT 1924.1000 1044.9400 1925.7000 1045.4200 ;
        RECT 1924.1000 1050.3800 1925.7000 1050.8600 ;
        RECT 1933.8400 1050.3800 1935.4400 1050.8600 ;
        RECT 1879.1000 1066.7000 1880.7000 1067.1800 ;
        RECT 1879.1000 1072.1400 1880.7000 1072.6200 ;
        RECT 1879.1000 1077.5800 1880.7000 1078.0600 ;
        RECT 1879.1000 1055.8200 1880.7000 1056.3000 ;
        RECT 1879.1000 1061.2600 1880.7000 1061.7400 ;
        RECT 1879.1000 1039.5000 1880.7000 1039.9800 ;
        RECT 1879.1000 1044.9400 1880.7000 1045.4200 ;
        RECT 1879.1000 1050.3800 1880.7000 1050.8600 ;
        RECT 1933.8400 1023.1800 1935.4400 1023.6600 ;
        RECT 1933.8400 1028.6200 1935.4400 1029.1000 ;
        RECT 1933.8400 1034.0600 1935.4400 1034.5400 ;
        RECT 1924.1000 1023.1800 1925.7000 1023.6600 ;
        RECT 1924.1000 1028.6200 1925.7000 1029.1000 ;
        RECT 1924.1000 1034.0600 1925.7000 1034.5400 ;
        RECT 1933.8400 1012.3000 1935.4400 1012.7800 ;
        RECT 1933.8400 1017.7400 1935.4400 1018.2200 ;
        RECT 1924.1000 1012.3000 1925.7000 1012.7800 ;
        RECT 1924.1000 1017.7400 1925.7000 1018.2200 ;
        RECT 1933.8400 995.9800 1935.4400 996.4600 ;
        RECT 1933.8400 1001.4200 1935.4400 1001.9000 ;
        RECT 1933.8400 1006.8600 1935.4400 1007.3400 ;
        RECT 1924.1000 995.9800 1925.7000 996.4600 ;
        RECT 1924.1000 1001.4200 1925.7000 1001.9000 ;
        RECT 1924.1000 1006.8600 1925.7000 1007.3400 ;
        RECT 1933.8400 985.1000 1935.4400 985.5800 ;
        RECT 1933.8400 990.5400 1935.4400 991.0200 ;
        RECT 1924.1000 985.1000 1925.7000 985.5800 ;
        RECT 1924.1000 990.5400 1925.7000 991.0200 ;
        RECT 1879.1000 1023.1800 1880.7000 1023.6600 ;
        RECT 1879.1000 1028.6200 1880.7000 1029.1000 ;
        RECT 1879.1000 1034.0600 1880.7000 1034.5400 ;
        RECT 1879.1000 1012.3000 1880.7000 1012.7800 ;
        RECT 1879.1000 1017.7400 1880.7000 1018.2200 ;
        RECT 1879.1000 995.9800 1880.7000 996.4600 ;
        RECT 1879.1000 1001.4200 1880.7000 1001.9000 ;
        RECT 1879.1000 1006.8600 1880.7000 1007.3400 ;
        RECT 1879.1000 985.1000 1880.7000 985.5800 ;
        RECT 1879.1000 990.5400 1880.7000 991.0200 ;
        RECT 1834.1000 1066.7000 1835.7000 1067.1800 ;
        RECT 1834.1000 1072.1400 1835.7000 1072.6200 ;
        RECT 1834.1000 1077.5800 1835.7000 1078.0600 ;
        RECT 1789.1000 1066.7000 1790.7000 1067.1800 ;
        RECT 1789.1000 1072.1400 1790.7000 1072.6200 ;
        RECT 1789.1000 1077.5800 1790.7000 1078.0600 ;
        RECT 1834.1000 1055.8200 1835.7000 1056.3000 ;
        RECT 1834.1000 1061.2600 1835.7000 1061.7400 ;
        RECT 1834.1000 1039.5000 1835.7000 1039.9800 ;
        RECT 1834.1000 1044.9400 1835.7000 1045.4200 ;
        RECT 1834.1000 1050.3800 1835.7000 1050.8600 ;
        RECT 1789.1000 1055.8200 1790.7000 1056.3000 ;
        RECT 1789.1000 1061.2600 1790.7000 1061.7400 ;
        RECT 1789.1000 1039.5000 1790.7000 1039.9800 ;
        RECT 1789.1000 1044.9400 1790.7000 1045.4200 ;
        RECT 1789.1000 1050.3800 1790.7000 1050.8600 ;
        RECT 1744.1000 1066.7000 1745.7000 1067.1800 ;
        RECT 1744.1000 1072.1400 1745.7000 1072.6200 ;
        RECT 1736.3400 1066.7000 1737.9400 1067.1800 ;
        RECT 1736.3400 1072.1400 1737.9400 1072.6200 ;
        RECT 1736.3400 1077.5800 1737.9400 1078.0600 ;
        RECT 1744.1000 1077.5800 1745.7000 1078.0600 ;
        RECT 1744.1000 1055.8200 1745.7000 1056.3000 ;
        RECT 1744.1000 1061.2600 1745.7000 1061.7400 ;
        RECT 1736.3400 1055.8200 1737.9400 1056.3000 ;
        RECT 1736.3400 1061.2600 1737.9400 1061.7400 ;
        RECT 1744.1000 1039.5000 1745.7000 1039.9800 ;
        RECT 1744.1000 1044.9400 1745.7000 1045.4200 ;
        RECT 1736.3400 1039.5000 1737.9400 1039.9800 ;
        RECT 1736.3400 1044.9400 1737.9400 1045.4200 ;
        RECT 1736.3400 1050.3800 1737.9400 1050.8600 ;
        RECT 1744.1000 1050.3800 1745.7000 1050.8600 ;
        RECT 1834.1000 1023.1800 1835.7000 1023.6600 ;
        RECT 1834.1000 1028.6200 1835.7000 1029.1000 ;
        RECT 1834.1000 1034.0600 1835.7000 1034.5400 ;
        RECT 1834.1000 1012.3000 1835.7000 1012.7800 ;
        RECT 1834.1000 1017.7400 1835.7000 1018.2200 ;
        RECT 1789.1000 1023.1800 1790.7000 1023.6600 ;
        RECT 1789.1000 1028.6200 1790.7000 1029.1000 ;
        RECT 1789.1000 1034.0600 1790.7000 1034.5400 ;
        RECT 1789.1000 1012.3000 1790.7000 1012.7800 ;
        RECT 1789.1000 1017.7400 1790.7000 1018.2200 ;
        RECT 1834.1000 995.9800 1835.7000 996.4600 ;
        RECT 1834.1000 1001.4200 1835.7000 1001.9000 ;
        RECT 1834.1000 1006.8600 1835.7000 1007.3400 ;
        RECT 1834.1000 985.1000 1835.7000 985.5800 ;
        RECT 1834.1000 990.5400 1835.7000 991.0200 ;
        RECT 1789.1000 995.9800 1790.7000 996.4600 ;
        RECT 1789.1000 1001.4200 1790.7000 1001.9000 ;
        RECT 1789.1000 1006.8600 1790.7000 1007.3400 ;
        RECT 1789.1000 985.1000 1790.7000 985.5800 ;
        RECT 1789.1000 990.5400 1790.7000 991.0200 ;
        RECT 1744.1000 1023.1800 1745.7000 1023.6600 ;
        RECT 1744.1000 1028.6200 1745.7000 1029.1000 ;
        RECT 1744.1000 1034.0600 1745.7000 1034.5400 ;
        RECT 1736.3400 1023.1800 1737.9400 1023.6600 ;
        RECT 1736.3400 1028.6200 1737.9400 1029.1000 ;
        RECT 1736.3400 1034.0600 1737.9400 1034.5400 ;
        RECT 1744.1000 1012.3000 1745.7000 1012.7800 ;
        RECT 1744.1000 1017.7400 1745.7000 1018.2200 ;
        RECT 1736.3400 1012.3000 1737.9400 1012.7800 ;
        RECT 1736.3400 1017.7400 1737.9400 1018.2200 ;
        RECT 1744.1000 995.9800 1745.7000 996.4600 ;
        RECT 1744.1000 1001.4200 1745.7000 1001.9000 ;
        RECT 1744.1000 1006.8600 1745.7000 1007.3400 ;
        RECT 1736.3400 995.9800 1737.9400 996.4600 ;
        RECT 1736.3400 1001.4200 1737.9400 1001.9000 ;
        RECT 1736.3400 1006.8600 1737.9400 1007.3400 ;
        RECT 1744.1000 985.1000 1745.7000 985.5800 ;
        RECT 1744.1000 990.5400 1745.7000 991.0200 ;
        RECT 1736.3400 985.1000 1737.9400 985.5800 ;
        RECT 1736.3400 990.5400 1737.9400 991.0200 ;
        RECT 1933.8400 968.7800 1935.4400 969.2600 ;
        RECT 1933.8400 974.2200 1935.4400 974.7000 ;
        RECT 1933.8400 979.6600 1935.4400 980.1400 ;
        RECT 1924.1000 968.7800 1925.7000 969.2600 ;
        RECT 1924.1000 974.2200 1925.7000 974.7000 ;
        RECT 1924.1000 979.6600 1925.7000 980.1400 ;
        RECT 1933.8400 957.9000 1935.4400 958.3800 ;
        RECT 1933.8400 963.3400 1935.4400 963.8200 ;
        RECT 1924.1000 957.9000 1925.7000 958.3800 ;
        RECT 1924.1000 963.3400 1925.7000 963.8200 ;
        RECT 1933.8400 941.5800 1935.4400 942.0600 ;
        RECT 1933.8400 947.0200 1935.4400 947.5000 ;
        RECT 1933.8400 952.4600 1935.4400 952.9400 ;
        RECT 1924.1000 941.5800 1925.7000 942.0600 ;
        RECT 1924.1000 947.0200 1925.7000 947.5000 ;
        RECT 1924.1000 952.4600 1925.7000 952.9400 ;
        RECT 1933.8400 930.7000 1935.4400 931.1800 ;
        RECT 1933.8400 936.1400 1935.4400 936.6200 ;
        RECT 1924.1000 930.7000 1925.7000 931.1800 ;
        RECT 1924.1000 936.1400 1925.7000 936.6200 ;
        RECT 1879.1000 968.7800 1880.7000 969.2600 ;
        RECT 1879.1000 974.2200 1880.7000 974.7000 ;
        RECT 1879.1000 979.6600 1880.7000 980.1400 ;
        RECT 1879.1000 957.9000 1880.7000 958.3800 ;
        RECT 1879.1000 963.3400 1880.7000 963.8200 ;
        RECT 1879.1000 941.5800 1880.7000 942.0600 ;
        RECT 1879.1000 947.0200 1880.7000 947.5000 ;
        RECT 1879.1000 952.4600 1880.7000 952.9400 ;
        RECT 1879.1000 930.7000 1880.7000 931.1800 ;
        RECT 1879.1000 936.1400 1880.7000 936.6200 ;
        RECT 1933.8400 914.3800 1935.4400 914.8600 ;
        RECT 1933.8400 919.8200 1935.4400 920.3000 ;
        RECT 1933.8400 925.2600 1935.4400 925.7400 ;
        RECT 1924.1000 914.3800 1925.7000 914.8600 ;
        RECT 1924.1000 919.8200 1925.7000 920.3000 ;
        RECT 1924.1000 925.2600 1925.7000 925.7400 ;
        RECT 1933.8400 903.5000 1935.4400 903.9800 ;
        RECT 1933.8400 908.9400 1935.4400 909.4200 ;
        RECT 1924.1000 903.5000 1925.7000 903.9800 ;
        RECT 1924.1000 908.9400 1925.7000 909.4200 ;
        RECT 1933.8400 887.1800 1935.4400 887.6600 ;
        RECT 1933.8400 892.6200 1935.4400 893.1000 ;
        RECT 1933.8400 898.0600 1935.4400 898.5400 ;
        RECT 1924.1000 887.1800 1925.7000 887.6600 ;
        RECT 1924.1000 892.6200 1925.7000 893.1000 ;
        RECT 1924.1000 898.0600 1925.7000 898.5400 ;
        RECT 1924.1000 881.7400 1925.7000 882.2200 ;
        RECT 1933.8400 881.7400 1935.4400 882.2200 ;
        RECT 1879.1000 914.3800 1880.7000 914.8600 ;
        RECT 1879.1000 919.8200 1880.7000 920.3000 ;
        RECT 1879.1000 925.2600 1880.7000 925.7400 ;
        RECT 1879.1000 903.5000 1880.7000 903.9800 ;
        RECT 1879.1000 908.9400 1880.7000 909.4200 ;
        RECT 1879.1000 887.1800 1880.7000 887.6600 ;
        RECT 1879.1000 892.6200 1880.7000 893.1000 ;
        RECT 1879.1000 898.0600 1880.7000 898.5400 ;
        RECT 1879.1000 881.7400 1880.7000 882.2200 ;
        RECT 1834.1000 968.7800 1835.7000 969.2600 ;
        RECT 1834.1000 974.2200 1835.7000 974.7000 ;
        RECT 1834.1000 979.6600 1835.7000 980.1400 ;
        RECT 1834.1000 957.9000 1835.7000 958.3800 ;
        RECT 1834.1000 963.3400 1835.7000 963.8200 ;
        RECT 1789.1000 968.7800 1790.7000 969.2600 ;
        RECT 1789.1000 974.2200 1790.7000 974.7000 ;
        RECT 1789.1000 979.6600 1790.7000 980.1400 ;
        RECT 1789.1000 957.9000 1790.7000 958.3800 ;
        RECT 1789.1000 963.3400 1790.7000 963.8200 ;
        RECT 1834.1000 941.5800 1835.7000 942.0600 ;
        RECT 1834.1000 947.0200 1835.7000 947.5000 ;
        RECT 1834.1000 952.4600 1835.7000 952.9400 ;
        RECT 1834.1000 930.7000 1835.7000 931.1800 ;
        RECT 1834.1000 936.1400 1835.7000 936.6200 ;
        RECT 1789.1000 941.5800 1790.7000 942.0600 ;
        RECT 1789.1000 947.0200 1790.7000 947.5000 ;
        RECT 1789.1000 952.4600 1790.7000 952.9400 ;
        RECT 1789.1000 930.7000 1790.7000 931.1800 ;
        RECT 1789.1000 936.1400 1790.7000 936.6200 ;
        RECT 1744.1000 968.7800 1745.7000 969.2600 ;
        RECT 1744.1000 974.2200 1745.7000 974.7000 ;
        RECT 1744.1000 979.6600 1745.7000 980.1400 ;
        RECT 1736.3400 968.7800 1737.9400 969.2600 ;
        RECT 1736.3400 974.2200 1737.9400 974.7000 ;
        RECT 1736.3400 979.6600 1737.9400 980.1400 ;
        RECT 1744.1000 957.9000 1745.7000 958.3800 ;
        RECT 1744.1000 963.3400 1745.7000 963.8200 ;
        RECT 1736.3400 957.9000 1737.9400 958.3800 ;
        RECT 1736.3400 963.3400 1737.9400 963.8200 ;
        RECT 1744.1000 941.5800 1745.7000 942.0600 ;
        RECT 1744.1000 947.0200 1745.7000 947.5000 ;
        RECT 1744.1000 952.4600 1745.7000 952.9400 ;
        RECT 1736.3400 941.5800 1737.9400 942.0600 ;
        RECT 1736.3400 947.0200 1737.9400 947.5000 ;
        RECT 1736.3400 952.4600 1737.9400 952.9400 ;
        RECT 1744.1000 930.7000 1745.7000 931.1800 ;
        RECT 1744.1000 936.1400 1745.7000 936.6200 ;
        RECT 1736.3400 930.7000 1737.9400 931.1800 ;
        RECT 1736.3400 936.1400 1737.9400 936.6200 ;
        RECT 1834.1000 914.3800 1835.7000 914.8600 ;
        RECT 1834.1000 919.8200 1835.7000 920.3000 ;
        RECT 1834.1000 925.2600 1835.7000 925.7400 ;
        RECT 1834.1000 903.5000 1835.7000 903.9800 ;
        RECT 1834.1000 908.9400 1835.7000 909.4200 ;
        RECT 1789.1000 914.3800 1790.7000 914.8600 ;
        RECT 1789.1000 919.8200 1790.7000 920.3000 ;
        RECT 1789.1000 925.2600 1790.7000 925.7400 ;
        RECT 1789.1000 903.5000 1790.7000 903.9800 ;
        RECT 1789.1000 908.9400 1790.7000 909.4200 ;
        RECT 1834.1000 887.1800 1835.7000 887.6600 ;
        RECT 1834.1000 892.6200 1835.7000 893.1000 ;
        RECT 1834.1000 898.0600 1835.7000 898.5400 ;
        RECT 1834.1000 881.7400 1835.7000 882.2200 ;
        RECT 1789.1000 887.1800 1790.7000 887.6600 ;
        RECT 1789.1000 892.6200 1790.7000 893.1000 ;
        RECT 1789.1000 898.0600 1790.7000 898.5400 ;
        RECT 1789.1000 881.7400 1790.7000 882.2200 ;
        RECT 1744.1000 914.3800 1745.7000 914.8600 ;
        RECT 1744.1000 919.8200 1745.7000 920.3000 ;
        RECT 1744.1000 925.2600 1745.7000 925.7400 ;
        RECT 1736.3400 914.3800 1737.9400 914.8600 ;
        RECT 1736.3400 919.8200 1737.9400 920.3000 ;
        RECT 1736.3400 925.2600 1737.9400 925.7400 ;
        RECT 1744.1000 903.5000 1745.7000 903.9800 ;
        RECT 1744.1000 908.9400 1745.7000 909.4200 ;
        RECT 1736.3400 903.5000 1737.9400 903.9800 ;
        RECT 1736.3400 908.9400 1737.9400 909.4200 ;
        RECT 1744.1000 887.1800 1745.7000 887.6600 ;
        RECT 1744.1000 892.6200 1745.7000 893.1000 ;
        RECT 1744.1000 898.0600 1745.7000 898.5400 ;
        RECT 1736.3400 887.1800 1737.9400 887.6600 ;
        RECT 1736.3400 892.6200 1737.9400 893.1000 ;
        RECT 1736.3400 898.0600 1737.9400 898.5400 ;
        RECT 1736.3400 881.7400 1737.9400 882.2200 ;
        RECT 1744.1000 881.7400 1745.7000 882.2200 ;
        RECT 1730.7800 1084.0500 1941.0000 1085.6500 ;
        RECT 1730.7800 877.5500 1941.0000 879.1500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 872.1200 1737.9400 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 1090.1600 1737.9400 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 872.1200 1935.4400 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 1090.1600 1935.4400 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 877.5500 1732.3800 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 877.5500 1941.0000 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 1084.0500 1732.3800 1085.6500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 1084.0500 1941.0000 1085.6500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 647.9100 1925.7000 856.0100 ;
        RECT 1879.1000 647.9100 1880.7000 856.0100 ;
        RECT 1834.1000 647.9100 1835.7000 856.0100 ;
        RECT 1789.1000 647.9100 1790.7000 856.0100 ;
        RECT 1744.1000 647.9100 1745.7000 856.0100 ;
        RECT 1933.8400 642.4800 1935.4400 862.1200 ;
        RECT 1736.3400 642.4800 1737.9400 862.1200 ;
      LAYER met3 ;
        RECT 1933.8400 837.0600 1935.4400 837.5400 ;
        RECT 1933.8400 842.5000 1935.4400 842.9800 ;
        RECT 1924.1000 837.0600 1925.7000 837.5400 ;
        RECT 1924.1000 842.5000 1925.7000 842.9800 ;
        RECT 1924.1000 847.9400 1925.7000 848.4200 ;
        RECT 1933.8400 847.9400 1935.4400 848.4200 ;
        RECT 1933.8400 826.1800 1935.4400 826.6600 ;
        RECT 1933.8400 831.6200 1935.4400 832.1000 ;
        RECT 1924.1000 826.1800 1925.7000 826.6600 ;
        RECT 1924.1000 831.6200 1925.7000 832.1000 ;
        RECT 1933.8400 809.8600 1935.4400 810.3400 ;
        RECT 1933.8400 815.3000 1935.4400 815.7800 ;
        RECT 1924.1000 809.8600 1925.7000 810.3400 ;
        RECT 1924.1000 815.3000 1925.7000 815.7800 ;
        RECT 1924.1000 820.7400 1925.7000 821.2200 ;
        RECT 1933.8400 820.7400 1935.4400 821.2200 ;
        RECT 1879.1000 837.0600 1880.7000 837.5400 ;
        RECT 1879.1000 842.5000 1880.7000 842.9800 ;
        RECT 1879.1000 847.9400 1880.7000 848.4200 ;
        RECT 1879.1000 826.1800 1880.7000 826.6600 ;
        RECT 1879.1000 831.6200 1880.7000 832.1000 ;
        RECT 1879.1000 809.8600 1880.7000 810.3400 ;
        RECT 1879.1000 815.3000 1880.7000 815.7800 ;
        RECT 1879.1000 820.7400 1880.7000 821.2200 ;
        RECT 1933.8400 793.5400 1935.4400 794.0200 ;
        RECT 1933.8400 798.9800 1935.4400 799.4600 ;
        RECT 1933.8400 804.4200 1935.4400 804.9000 ;
        RECT 1924.1000 793.5400 1925.7000 794.0200 ;
        RECT 1924.1000 798.9800 1925.7000 799.4600 ;
        RECT 1924.1000 804.4200 1925.7000 804.9000 ;
        RECT 1933.8400 782.6600 1935.4400 783.1400 ;
        RECT 1933.8400 788.1000 1935.4400 788.5800 ;
        RECT 1924.1000 782.6600 1925.7000 783.1400 ;
        RECT 1924.1000 788.1000 1925.7000 788.5800 ;
        RECT 1933.8400 766.3400 1935.4400 766.8200 ;
        RECT 1933.8400 771.7800 1935.4400 772.2600 ;
        RECT 1933.8400 777.2200 1935.4400 777.7000 ;
        RECT 1924.1000 766.3400 1925.7000 766.8200 ;
        RECT 1924.1000 771.7800 1925.7000 772.2600 ;
        RECT 1924.1000 777.2200 1925.7000 777.7000 ;
        RECT 1933.8400 755.4600 1935.4400 755.9400 ;
        RECT 1933.8400 760.9000 1935.4400 761.3800 ;
        RECT 1924.1000 755.4600 1925.7000 755.9400 ;
        RECT 1924.1000 760.9000 1925.7000 761.3800 ;
        RECT 1879.1000 793.5400 1880.7000 794.0200 ;
        RECT 1879.1000 798.9800 1880.7000 799.4600 ;
        RECT 1879.1000 804.4200 1880.7000 804.9000 ;
        RECT 1879.1000 782.6600 1880.7000 783.1400 ;
        RECT 1879.1000 788.1000 1880.7000 788.5800 ;
        RECT 1879.1000 766.3400 1880.7000 766.8200 ;
        RECT 1879.1000 771.7800 1880.7000 772.2600 ;
        RECT 1879.1000 777.2200 1880.7000 777.7000 ;
        RECT 1879.1000 755.4600 1880.7000 755.9400 ;
        RECT 1879.1000 760.9000 1880.7000 761.3800 ;
        RECT 1834.1000 837.0600 1835.7000 837.5400 ;
        RECT 1834.1000 842.5000 1835.7000 842.9800 ;
        RECT 1834.1000 847.9400 1835.7000 848.4200 ;
        RECT 1789.1000 837.0600 1790.7000 837.5400 ;
        RECT 1789.1000 842.5000 1790.7000 842.9800 ;
        RECT 1789.1000 847.9400 1790.7000 848.4200 ;
        RECT 1834.1000 826.1800 1835.7000 826.6600 ;
        RECT 1834.1000 831.6200 1835.7000 832.1000 ;
        RECT 1834.1000 809.8600 1835.7000 810.3400 ;
        RECT 1834.1000 815.3000 1835.7000 815.7800 ;
        RECT 1834.1000 820.7400 1835.7000 821.2200 ;
        RECT 1789.1000 826.1800 1790.7000 826.6600 ;
        RECT 1789.1000 831.6200 1790.7000 832.1000 ;
        RECT 1789.1000 809.8600 1790.7000 810.3400 ;
        RECT 1789.1000 815.3000 1790.7000 815.7800 ;
        RECT 1789.1000 820.7400 1790.7000 821.2200 ;
        RECT 1744.1000 837.0600 1745.7000 837.5400 ;
        RECT 1744.1000 842.5000 1745.7000 842.9800 ;
        RECT 1736.3400 837.0600 1737.9400 837.5400 ;
        RECT 1736.3400 842.5000 1737.9400 842.9800 ;
        RECT 1736.3400 847.9400 1737.9400 848.4200 ;
        RECT 1744.1000 847.9400 1745.7000 848.4200 ;
        RECT 1744.1000 826.1800 1745.7000 826.6600 ;
        RECT 1744.1000 831.6200 1745.7000 832.1000 ;
        RECT 1736.3400 826.1800 1737.9400 826.6600 ;
        RECT 1736.3400 831.6200 1737.9400 832.1000 ;
        RECT 1744.1000 809.8600 1745.7000 810.3400 ;
        RECT 1744.1000 815.3000 1745.7000 815.7800 ;
        RECT 1736.3400 809.8600 1737.9400 810.3400 ;
        RECT 1736.3400 815.3000 1737.9400 815.7800 ;
        RECT 1736.3400 820.7400 1737.9400 821.2200 ;
        RECT 1744.1000 820.7400 1745.7000 821.2200 ;
        RECT 1834.1000 793.5400 1835.7000 794.0200 ;
        RECT 1834.1000 798.9800 1835.7000 799.4600 ;
        RECT 1834.1000 804.4200 1835.7000 804.9000 ;
        RECT 1834.1000 782.6600 1835.7000 783.1400 ;
        RECT 1834.1000 788.1000 1835.7000 788.5800 ;
        RECT 1789.1000 793.5400 1790.7000 794.0200 ;
        RECT 1789.1000 798.9800 1790.7000 799.4600 ;
        RECT 1789.1000 804.4200 1790.7000 804.9000 ;
        RECT 1789.1000 782.6600 1790.7000 783.1400 ;
        RECT 1789.1000 788.1000 1790.7000 788.5800 ;
        RECT 1834.1000 766.3400 1835.7000 766.8200 ;
        RECT 1834.1000 771.7800 1835.7000 772.2600 ;
        RECT 1834.1000 777.2200 1835.7000 777.7000 ;
        RECT 1834.1000 755.4600 1835.7000 755.9400 ;
        RECT 1834.1000 760.9000 1835.7000 761.3800 ;
        RECT 1789.1000 766.3400 1790.7000 766.8200 ;
        RECT 1789.1000 771.7800 1790.7000 772.2600 ;
        RECT 1789.1000 777.2200 1790.7000 777.7000 ;
        RECT 1789.1000 755.4600 1790.7000 755.9400 ;
        RECT 1789.1000 760.9000 1790.7000 761.3800 ;
        RECT 1744.1000 793.5400 1745.7000 794.0200 ;
        RECT 1744.1000 798.9800 1745.7000 799.4600 ;
        RECT 1744.1000 804.4200 1745.7000 804.9000 ;
        RECT 1736.3400 793.5400 1737.9400 794.0200 ;
        RECT 1736.3400 798.9800 1737.9400 799.4600 ;
        RECT 1736.3400 804.4200 1737.9400 804.9000 ;
        RECT 1744.1000 782.6600 1745.7000 783.1400 ;
        RECT 1744.1000 788.1000 1745.7000 788.5800 ;
        RECT 1736.3400 782.6600 1737.9400 783.1400 ;
        RECT 1736.3400 788.1000 1737.9400 788.5800 ;
        RECT 1744.1000 766.3400 1745.7000 766.8200 ;
        RECT 1744.1000 771.7800 1745.7000 772.2600 ;
        RECT 1744.1000 777.2200 1745.7000 777.7000 ;
        RECT 1736.3400 766.3400 1737.9400 766.8200 ;
        RECT 1736.3400 771.7800 1737.9400 772.2600 ;
        RECT 1736.3400 777.2200 1737.9400 777.7000 ;
        RECT 1744.1000 755.4600 1745.7000 755.9400 ;
        RECT 1744.1000 760.9000 1745.7000 761.3800 ;
        RECT 1736.3400 755.4600 1737.9400 755.9400 ;
        RECT 1736.3400 760.9000 1737.9400 761.3800 ;
        RECT 1933.8400 739.1400 1935.4400 739.6200 ;
        RECT 1933.8400 744.5800 1935.4400 745.0600 ;
        RECT 1933.8400 750.0200 1935.4400 750.5000 ;
        RECT 1924.1000 739.1400 1925.7000 739.6200 ;
        RECT 1924.1000 744.5800 1925.7000 745.0600 ;
        RECT 1924.1000 750.0200 1925.7000 750.5000 ;
        RECT 1933.8400 728.2600 1935.4400 728.7400 ;
        RECT 1933.8400 733.7000 1935.4400 734.1800 ;
        RECT 1924.1000 728.2600 1925.7000 728.7400 ;
        RECT 1924.1000 733.7000 1925.7000 734.1800 ;
        RECT 1933.8400 711.9400 1935.4400 712.4200 ;
        RECT 1933.8400 717.3800 1935.4400 717.8600 ;
        RECT 1933.8400 722.8200 1935.4400 723.3000 ;
        RECT 1924.1000 711.9400 1925.7000 712.4200 ;
        RECT 1924.1000 717.3800 1925.7000 717.8600 ;
        RECT 1924.1000 722.8200 1925.7000 723.3000 ;
        RECT 1933.8400 701.0600 1935.4400 701.5400 ;
        RECT 1933.8400 706.5000 1935.4400 706.9800 ;
        RECT 1924.1000 701.0600 1925.7000 701.5400 ;
        RECT 1924.1000 706.5000 1925.7000 706.9800 ;
        RECT 1879.1000 739.1400 1880.7000 739.6200 ;
        RECT 1879.1000 744.5800 1880.7000 745.0600 ;
        RECT 1879.1000 750.0200 1880.7000 750.5000 ;
        RECT 1879.1000 728.2600 1880.7000 728.7400 ;
        RECT 1879.1000 733.7000 1880.7000 734.1800 ;
        RECT 1879.1000 711.9400 1880.7000 712.4200 ;
        RECT 1879.1000 717.3800 1880.7000 717.8600 ;
        RECT 1879.1000 722.8200 1880.7000 723.3000 ;
        RECT 1879.1000 701.0600 1880.7000 701.5400 ;
        RECT 1879.1000 706.5000 1880.7000 706.9800 ;
        RECT 1933.8400 684.7400 1935.4400 685.2200 ;
        RECT 1933.8400 690.1800 1935.4400 690.6600 ;
        RECT 1933.8400 695.6200 1935.4400 696.1000 ;
        RECT 1924.1000 684.7400 1925.7000 685.2200 ;
        RECT 1924.1000 690.1800 1925.7000 690.6600 ;
        RECT 1924.1000 695.6200 1925.7000 696.1000 ;
        RECT 1933.8400 673.8600 1935.4400 674.3400 ;
        RECT 1933.8400 679.3000 1935.4400 679.7800 ;
        RECT 1924.1000 673.8600 1925.7000 674.3400 ;
        RECT 1924.1000 679.3000 1925.7000 679.7800 ;
        RECT 1933.8400 657.5400 1935.4400 658.0200 ;
        RECT 1933.8400 662.9800 1935.4400 663.4600 ;
        RECT 1933.8400 668.4200 1935.4400 668.9000 ;
        RECT 1924.1000 657.5400 1925.7000 658.0200 ;
        RECT 1924.1000 662.9800 1925.7000 663.4600 ;
        RECT 1924.1000 668.4200 1925.7000 668.9000 ;
        RECT 1924.1000 652.1000 1925.7000 652.5800 ;
        RECT 1933.8400 652.1000 1935.4400 652.5800 ;
        RECT 1879.1000 684.7400 1880.7000 685.2200 ;
        RECT 1879.1000 690.1800 1880.7000 690.6600 ;
        RECT 1879.1000 695.6200 1880.7000 696.1000 ;
        RECT 1879.1000 673.8600 1880.7000 674.3400 ;
        RECT 1879.1000 679.3000 1880.7000 679.7800 ;
        RECT 1879.1000 657.5400 1880.7000 658.0200 ;
        RECT 1879.1000 662.9800 1880.7000 663.4600 ;
        RECT 1879.1000 668.4200 1880.7000 668.9000 ;
        RECT 1879.1000 652.1000 1880.7000 652.5800 ;
        RECT 1834.1000 739.1400 1835.7000 739.6200 ;
        RECT 1834.1000 744.5800 1835.7000 745.0600 ;
        RECT 1834.1000 750.0200 1835.7000 750.5000 ;
        RECT 1834.1000 728.2600 1835.7000 728.7400 ;
        RECT 1834.1000 733.7000 1835.7000 734.1800 ;
        RECT 1789.1000 739.1400 1790.7000 739.6200 ;
        RECT 1789.1000 744.5800 1790.7000 745.0600 ;
        RECT 1789.1000 750.0200 1790.7000 750.5000 ;
        RECT 1789.1000 728.2600 1790.7000 728.7400 ;
        RECT 1789.1000 733.7000 1790.7000 734.1800 ;
        RECT 1834.1000 711.9400 1835.7000 712.4200 ;
        RECT 1834.1000 717.3800 1835.7000 717.8600 ;
        RECT 1834.1000 722.8200 1835.7000 723.3000 ;
        RECT 1834.1000 701.0600 1835.7000 701.5400 ;
        RECT 1834.1000 706.5000 1835.7000 706.9800 ;
        RECT 1789.1000 711.9400 1790.7000 712.4200 ;
        RECT 1789.1000 717.3800 1790.7000 717.8600 ;
        RECT 1789.1000 722.8200 1790.7000 723.3000 ;
        RECT 1789.1000 701.0600 1790.7000 701.5400 ;
        RECT 1789.1000 706.5000 1790.7000 706.9800 ;
        RECT 1744.1000 739.1400 1745.7000 739.6200 ;
        RECT 1744.1000 744.5800 1745.7000 745.0600 ;
        RECT 1744.1000 750.0200 1745.7000 750.5000 ;
        RECT 1736.3400 739.1400 1737.9400 739.6200 ;
        RECT 1736.3400 744.5800 1737.9400 745.0600 ;
        RECT 1736.3400 750.0200 1737.9400 750.5000 ;
        RECT 1744.1000 728.2600 1745.7000 728.7400 ;
        RECT 1744.1000 733.7000 1745.7000 734.1800 ;
        RECT 1736.3400 728.2600 1737.9400 728.7400 ;
        RECT 1736.3400 733.7000 1737.9400 734.1800 ;
        RECT 1744.1000 711.9400 1745.7000 712.4200 ;
        RECT 1744.1000 717.3800 1745.7000 717.8600 ;
        RECT 1744.1000 722.8200 1745.7000 723.3000 ;
        RECT 1736.3400 711.9400 1737.9400 712.4200 ;
        RECT 1736.3400 717.3800 1737.9400 717.8600 ;
        RECT 1736.3400 722.8200 1737.9400 723.3000 ;
        RECT 1744.1000 701.0600 1745.7000 701.5400 ;
        RECT 1744.1000 706.5000 1745.7000 706.9800 ;
        RECT 1736.3400 701.0600 1737.9400 701.5400 ;
        RECT 1736.3400 706.5000 1737.9400 706.9800 ;
        RECT 1834.1000 684.7400 1835.7000 685.2200 ;
        RECT 1834.1000 690.1800 1835.7000 690.6600 ;
        RECT 1834.1000 695.6200 1835.7000 696.1000 ;
        RECT 1834.1000 673.8600 1835.7000 674.3400 ;
        RECT 1834.1000 679.3000 1835.7000 679.7800 ;
        RECT 1789.1000 684.7400 1790.7000 685.2200 ;
        RECT 1789.1000 690.1800 1790.7000 690.6600 ;
        RECT 1789.1000 695.6200 1790.7000 696.1000 ;
        RECT 1789.1000 673.8600 1790.7000 674.3400 ;
        RECT 1789.1000 679.3000 1790.7000 679.7800 ;
        RECT 1834.1000 657.5400 1835.7000 658.0200 ;
        RECT 1834.1000 662.9800 1835.7000 663.4600 ;
        RECT 1834.1000 668.4200 1835.7000 668.9000 ;
        RECT 1834.1000 652.1000 1835.7000 652.5800 ;
        RECT 1789.1000 657.5400 1790.7000 658.0200 ;
        RECT 1789.1000 662.9800 1790.7000 663.4600 ;
        RECT 1789.1000 668.4200 1790.7000 668.9000 ;
        RECT 1789.1000 652.1000 1790.7000 652.5800 ;
        RECT 1744.1000 684.7400 1745.7000 685.2200 ;
        RECT 1744.1000 690.1800 1745.7000 690.6600 ;
        RECT 1744.1000 695.6200 1745.7000 696.1000 ;
        RECT 1736.3400 684.7400 1737.9400 685.2200 ;
        RECT 1736.3400 690.1800 1737.9400 690.6600 ;
        RECT 1736.3400 695.6200 1737.9400 696.1000 ;
        RECT 1744.1000 673.8600 1745.7000 674.3400 ;
        RECT 1744.1000 679.3000 1745.7000 679.7800 ;
        RECT 1736.3400 673.8600 1737.9400 674.3400 ;
        RECT 1736.3400 679.3000 1737.9400 679.7800 ;
        RECT 1744.1000 657.5400 1745.7000 658.0200 ;
        RECT 1744.1000 662.9800 1745.7000 663.4600 ;
        RECT 1744.1000 668.4200 1745.7000 668.9000 ;
        RECT 1736.3400 657.5400 1737.9400 658.0200 ;
        RECT 1736.3400 662.9800 1737.9400 663.4600 ;
        RECT 1736.3400 668.4200 1737.9400 668.9000 ;
        RECT 1736.3400 652.1000 1737.9400 652.5800 ;
        RECT 1744.1000 652.1000 1745.7000 652.5800 ;
        RECT 1730.7800 854.4100 1941.0000 856.0100 ;
        RECT 1730.7800 647.9100 1941.0000 649.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 642.4800 1737.9400 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 860.5200 1737.9400 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 642.4800 1935.4400 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 860.5200 1935.4400 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 647.9100 1732.3800 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 647.9100 1941.0000 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 854.4100 1732.3800 856.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 854.4100 1941.0000 856.0100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 1924.1000 418.2700 1925.7000 626.3700 ;
        RECT 1879.1000 418.2700 1880.7000 626.3700 ;
        RECT 1834.1000 418.2700 1835.7000 626.3700 ;
        RECT 1789.1000 418.2700 1790.7000 626.3700 ;
        RECT 1744.1000 418.2700 1745.7000 626.3700 ;
        RECT 1933.8400 412.8400 1935.4400 632.4800 ;
        RECT 1736.3400 412.8400 1737.9400 632.4800 ;
      LAYER met3 ;
        RECT 1933.8400 607.4200 1935.4400 607.9000 ;
        RECT 1933.8400 612.8600 1935.4400 613.3400 ;
        RECT 1924.1000 607.4200 1925.7000 607.9000 ;
        RECT 1924.1000 612.8600 1925.7000 613.3400 ;
        RECT 1924.1000 618.3000 1925.7000 618.7800 ;
        RECT 1933.8400 618.3000 1935.4400 618.7800 ;
        RECT 1933.8400 596.5400 1935.4400 597.0200 ;
        RECT 1933.8400 601.9800 1935.4400 602.4600 ;
        RECT 1924.1000 596.5400 1925.7000 597.0200 ;
        RECT 1924.1000 601.9800 1925.7000 602.4600 ;
        RECT 1933.8400 580.2200 1935.4400 580.7000 ;
        RECT 1933.8400 585.6600 1935.4400 586.1400 ;
        RECT 1924.1000 580.2200 1925.7000 580.7000 ;
        RECT 1924.1000 585.6600 1925.7000 586.1400 ;
        RECT 1924.1000 591.1000 1925.7000 591.5800 ;
        RECT 1933.8400 591.1000 1935.4400 591.5800 ;
        RECT 1879.1000 607.4200 1880.7000 607.9000 ;
        RECT 1879.1000 612.8600 1880.7000 613.3400 ;
        RECT 1879.1000 618.3000 1880.7000 618.7800 ;
        RECT 1879.1000 596.5400 1880.7000 597.0200 ;
        RECT 1879.1000 601.9800 1880.7000 602.4600 ;
        RECT 1879.1000 580.2200 1880.7000 580.7000 ;
        RECT 1879.1000 585.6600 1880.7000 586.1400 ;
        RECT 1879.1000 591.1000 1880.7000 591.5800 ;
        RECT 1933.8400 563.9000 1935.4400 564.3800 ;
        RECT 1933.8400 569.3400 1935.4400 569.8200 ;
        RECT 1933.8400 574.7800 1935.4400 575.2600 ;
        RECT 1924.1000 563.9000 1925.7000 564.3800 ;
        RECT 1924.1000 569.3400 1925.7000 569.8200 ;
        RECT 1924.1000 574.7800 1925.7000 575.2600 ;
        RECT 1933.8400 553.0200 1935.4400 553.5000 ;
        RECT 1933.8400 558.4600 1935.4400 558.9400 ;
        RECT 1924.1000 553.0200 1925.7000 553.5000 ;
        RECT 1924.1000 558.4600 1925.7000 558.9400 ;
        RECT 1933.8400 536.7000 1935.4400 537.1800 ;
        RECT 1933.8400 542.1400 1935.4400 542.6200 ;
        RECT 1933.8400 547.5800 1935.4400 548.0600 ;
        RECT 1924.1000 536.7000 1925.7000 537.1800 ;
        RECT 1924.1000 542.1400 1925.7000 542.6200 ;
        RECT 1924.1000 547.5800 1925.7000 548.0600 ;
        RECT 1933.8400 525.8200 1935.4400 526.3000 ;
        RECT 1933.8400 531.2600 1935.4400 531.7400 ;
        RECT 1924.1000 525.8200 1925.7000 526.3000 ;
        RECT 1924.1000 531.2600 1925.7000 531.7400 ;
        RECT 1879.1000 563.9000 1880.7000 564.3800 ;
        RECT 1879.1000 569.3400 1880.7000 569.8200 ;
        RECT 1879.1000 574.7800 1880.7000 575.2600 ;
        RECT 1879.1000 553.0200 1880.7000 553.5000 ;
        RECT 1879.1000 558.4600 1880.7000 558.9400 ;
        RECT 1879.1000 536.7000 1880.7000 537.1800 ;
        RECT 1879.1000 542.1400 1880.7000 542.6200 ;
        RECT 1879.1000 547.5800 1880.7000 548.0600 ;
        RECT 1879.1000 525.8200 1880.7000 526.3000 ;
        RECT 1879.1000 531.2600 1880.7000 531.7400 ;
        RECT 1834.1000 607.4200 1835.7000 607.9000 ;
        RECT 1834.1000 612.8600 1835.7000 613.3400 ;
        RECT 1834.1000 618.3000 1835.7000 618.7800 ;
        RECT 1789.1000 607.4200 1790.7000 607.9000 ;
        RECT 1789.1000 612.8600 1790.7000 613.3400 ;
        RECT 1789.1000 618.3000 1790.7000 618.7800 ;
        RECT 1834.1000 596.5400 1835.7000 597.0200 ;
        RECT 1834.1000 601.9800 1835.7000 602.4600 ;
        RECT 1834.1000 580.2200 1835.7000 580.7000 ;
        RECT 1834.1000 585.6600 1835.7000 586.1400 ;
        RECT 1834.1000 591.1000 1835.7000 591.5800 ;
        RECT 1789.1000 596.5400 1790.7000 597.0200 ;
        RECT 1789.1000 601.9800 1790.7000 602.4600 ;
        RECT 1789.1000 580.2200 1790.7000 580.7000 ;
        RECT 1789.1000 585.6600 1790.7000 586.1400 ;
        RECT 1789.1000 591.1000 1790.7000 591.5800 ;
        RECT 1744.1000 607.4200 1745.7000 607.9000 ;
        RECT 1744.1000 612.8600 1745.7000 613.3400 ;
        RECT 1736.3400 607.4200 1737.9400 607.9000 ;
        RECT 1736.3400 612.8600 1737.9400 613.3400 ;
        RECT 1736.3400 618.3000 1737.9400 618.7800 ;
        RECT 1744.1000 618.3000 1745.7000 618.7800 ;
        RECT 1744.1000 596.5400 1745.7000 597.0200 ;
        RECT 1744.1000 601.9800 1745.7000 602.4600 ;
        RECT 1736.3400 596.5400 1737.9400 597.0200 ;
        RECT 1736.3400 601.9800 1737.9400 602.4600 ;
        RECT 1744.1000 580.2200 1745.7000 580.7000 ;
        RECT 1744.1000 585.6600 1745.7000 586.1400 ;
        RECT 1736.3400 580.2200 1737.9400 580.7000 ;
        RECT 1736.3400 585.6600 1737.9400 586.1400 ;
        RECT 1736.3400 591.1000 1737.9400 591.5800 ;
        RECT 1744.1000 591.1000 1745.7000 591.5800 ;
        RECT 1834.1000 563.9000 1835.7000 564.3800 ;
        RECT 1834.1000 569.3400 1835.7000 569.8200 ;
        RECT 1834.1000 574.7800 1835.7000 575.2600 ;
        RECT 1834.1000 553.0200 1835.7000 553.5000 ;
        RECT 1834.1000 558.4600 1835.7000 558.9400 ;
        RECT 1789.1000 563.9000 1790.7000 564.3800 ;
        RECT 1789.1000 569.3400 1790.7000 569.8200 ;
        RECT 1789.1000 574.7800 1790.7000 575.2600 ;
        RECT 1789.1000 553.0200 1790.7000 553.5000 ;
        RECT 1789.1000 558.4600 1790.7000 558.9400 ;
        RECT 1834.1000 536.7000 1835.7000 537.1800 ;
        RECT 1834.1000 542.1400 1835.7000 542.6200 ;
        RECT 1834.1000 547.5800 1835.7000 548.0600 ;
        RECT 1834.1000 525.8200 1835.7000 526.3000 ;
        RECT 1834.1000 531.2600 1835.7000 531.7400 ;
        RECT 1789.1000 536.7000 1790.7000 537.1800 ;
        RECT 1789.1000 542.1400 1790.7000 542.6200 ;
        RECT 1789.1000 547.5800 1790.7000 548.0600 ;
        RECT 1789.1000 525.8200 1790.7000 526.3000 ;
        RECT 1789.1000 531.2600 1790.7000 531.7400 ;
        RECT 1744.1000 563.9000 1745.7000 564.3800 ;
        RECT 1744.1000 569.3400 1745.7000 569.8200 ;
        RECT 1744.1000 574.7800 1745.7000 575.2600 ;
        RECT 1736.3400 563.9000 1737.9400 564.3800 ;
        RECT 1736.3400 569.3400 1737.9400 569.8200 ;
        RECT 1736.3400 574.7800 1737.9400 575.2600 ;
        RECT 1744.1000 553.0200 1745.7000 553.5000 ;
        RECT 1744.1000 558.4600 1745.7000 558.9400 ;
        RECT 1736.3400 553.0200 1737.9400 553.5000 ;
        RECT 1736.3400 558.4600 1737.9400 558.9400 ;
        RECT 1744.1000 536.7000 1745.7000 537.1800 ;
        RECT 1744.1000 542.1400 1745.7000 542.6200 ;
        RECT 1744.1000 547.5800 1745.7000 548.0600 ;
        RECT 1736.3400 536.7000 1737.9400 537.1800 ;
        RECT 1736.3400 542.1400 1737.9400 542.6200 ;
        RECT 1736.3400 547.5800 1737.9400 548.0600 ;
        RECT 1744.1000 525.8200 1745.7000 526.3000 ;
        RECT 1744.1000 531.2600 1745.7000 531.7400 ;
        RECT 1736.3400 525.8200 1737.9400 526.3000 ;
        RECT 1736.3400 531.2600 1737.9400 531.7400 ;
        RECT 1933.8400 509.5000 1935.4400 509.9800 ;
        RECT 1933.8400 514.9400 1935.4400 515.4200 ;
        RECT 1933.8400 520.3800 1935.4400 520.8600 ;
        RECT 1924.1000 509.5000 1925.7000 509.9800 ;
        RECT 1924.1000 514.9400 1925.7000 515.4200 ;
        RECT 1924.1000 520.3800 1925.7000 520.8600 ;
        RECT 1933.8400 498.6200 1935.4400 499.1000 ;
        RECT 1933.8400 504.0600 1935.4400 504.5400 ;
        RECT 1924.1000 498.6200 1925.7000 499.1000 ;
        RECT 1924.1000 504.0600 1925.7000 504.5400 ;
        RECT 1933.8400 482.3000 1935.4400 482.7800 ;
        RECT 1933.8400 487.7400 1935.4400 488.2200 ;
        RECT 1933.8400 493.1800 1935.4400 493.6600 ;
        RECT 1924.1000 482.3000 1925.7000 482.7800 ;
        RECT 1924.1000 487.7400 1925.7000 488.2200 ;
        RECT 1924.1000 493.1800 1925.7000 493.6600 ;
        RECT 1933.8400 471.4200 1935.4400 471.9000 ;
        RECT 1933.8400 476.8600 1935.4400 477.3400 ;
        RECT 1924.1000 471.4200 1925.7000 471.9000 ;
        RECT 1924.1000 476.8600 1925.7000 477.3400 ;
        RECT 1879.1000 509.5000 1880.7000 509.9800 ;
        RECT 1879.1000 514.9400 1880.7000 515.4200 ;
        RECT 1879.1000 520.3800 1880.7000 520.8600 ;
        RECT 1879.1000 498.6200 1880.7000 499.1000 ;
        RECT 1879.1000 504.0600 1880.7000 504.5400 ;
        RECT 1879.1000 482.3000 1880.7000 482.7800 ;
        RECT 1879.1000 487.7400 1880.7000 488.2200 ;
        RECT 1879.1000 493.1800 1880.7000 493.6600 ;
        RECT 1879.1000 471.4200 1880.7000 471.9000 ;
        RECT 1879.1000 476.8600 1880.7000 477.3400 ;
        RECT 1933.8400 455.1000 1935.4400 455.5800 ;
        RECT 1933.8400 460.5400 1935.4400 461.0200 ;
        RECT 1933.8400 465.9800 1935.4400 466.4600 ;
        RECT 1924.1000 455.1000 1925.7000 455.5800 ;
        RECT 1924.1000 460.5400 1925.7000 461.0200 ;
        RECT 1924.1000 465.9800 1925.7000 466.4600 ;
        RECT 1933.8400 444.2200 1935.4400 444.7000 ;
        RECT 1933.8400 449.6600 1935.4400 450.1400 ;
        RECT 1924.1000 444.2200 1925.7000 444.7000 ;
        RECT 1924.1000 449.6600 1925.7000 450.1400 ;
        RECT 1933.8400 427.9000 1935.4400 428.3800 ;
        RECT 1933.8400 433.3400 1935.4400 433.8200 ;
        RECT 1933.8400 438.7800 1935.4400 439.2600 ;
        RECT 1924.1000 427.9000 1925.7000 428.3800 ;
        RECT 1924.1000 433.3400 1925.7000 433.8200 ;
        RECT 1924.1000 438.7800 1925.7000 439.2600 ;
        RECT 1924.1000 422.4600 1925.7000 422.9400 ;
        RECT 1933.8400 422.4600 1935.4400 422.9400 ;
        RECT 1879.1000 455.1000 1880.7000 455.5800 ;
        RECT 1879.1000 460.5400 1880.7000 461.0200 ;
        RECT 1879.1000 465.9800 1880.7000 466.4600 ;
        RECT 1879.1000 444.2200 1880.7000 444.7000 ;
        RECT 1879.1000 449.6600 1880.7000 450.1400 ;
        RECT 1879.1000 427.9000 1880.7000 428.3800 ;
        RECT 1879.1000 433.3400 1880.7000 433.8200 ;
        RECT 1879.1000 438.7800 1880.7000 439.2600 ;
        RECT 1879.1000 422.4600 1880.7000 422.9400 ;
        RECT 1834.1000 509.5000 1835.7000 509.9800 ;
        RECT 1834.1000 514.9400 1835.7000 515.4200 ;
        RECT 1834.1000 520.3800 1835.7000 520.8600 ;
        RECT 1834.1000 498.6200 1835.7000 499.1000 ;
        RECT 1834.1000 504.0600 1835.7000 504.5400 ;
        RECT 1789.1000 509.5000 1790.7000 509.9800 ;
        RECT 1789.1000 514.9400 1790.7000 515.4200 ;
        RECT 1789.1000 520.3800 1790.7000 520.8600 ;
        RECT 1789.1000 498.6200 1790.7000 499.1000 ;
        RECT 1789.1000 504.0600 1790.7000 504.5400 ;
        RECT 1834.1000 482.3000 1835.7000 482.7800 ;
        RECT 1834.1000 487.7400 1835.7000 488.2200 ;
        RECT 1834.1000 493.1800 1835.7000 493.6600 ;
        RECT 1834.1000 471.4200 1835.7000 471.9000 ;
        RECT 1834.1000 476.8600 1835.7000 477.3400 ;
        RECT 1789.1000 482.3000 1790.7000 482.7800 ;
        RECT 1789.1000 487.7400 1790.7000 488.2200 ;
        RECT 1789.1000 493.1800 1790.7000 493.6600 ;
        RECT 1789.1000 471.4200 1790.7000 471.9000 ;
        RECT 1789.1000 476.8600 1790.7000 477.3400 ;
        RECT 1744.1000 509.5000 1745.7000 509.9800 ;
        RECT 1744.1000 514.9400 1745.7000 515.4200 ;
        RECT 1744.1000 520.3800 1745.7000 520.8600 ;
        RECT 1736.3400 509.5000 1737.9400 509.9800 ;
        RECT 1736.3400 514.9400 1737.9400 515.4200 ;
        RECT 1736.3400 520.3800 1737.9400 520.8600 ;
        RECT 1744.1000 498.6200 1745.7000 499.1000 ;
        RECT 1744.1000 504.0600 1745.7000 504.5400 ;
        RECT 1736.3400 498.6200 1737.9400 499.1000 ;
        RECT 1736.3400 504.0600 1737.9400 504.5400 ;
        RECT 1744.1000 482.3000 1745.7000 482.7800 ;
        RECT 1744.1000 487.7400 1745.7000 488.2200 ;
        RECT 1744.1000 493.1800 1745.7000 493.6600 ;
        RECT 1736.3400 482.3000 1737.9400 482.7800 ;
        RECT 1736.3400 487.7400 1737.9400 488.2200 ;
        RECT 1736.3400 493.1800 1737.9400 493.6600 ;
        RECT 1744.1000 471.4200 1745.7000 471.9000 ;
        RECT 1744.1000 476.8600 1745.7000 477.3400 ;
        RECT 1736.3400 471.4200 1737.9400 471.9000 ;
        RECT 1736.3400 476.8600 1737.9400 477.3400 ;
        RECT 1834.1000 455.1000 1835.7000 455.5800 ;
        RECT 1834.1000 460.5400 1835.7000 461.0200 ;
        RECT 1834.1000 465.9800 1835.7000 466.4600 ;
        RECT 1834.1000 444.2200 1835.7000 444.7000 ;
        RECT 1834.1000 449.6600 1835.7000 450.1400 ;
        RECT 1789.1000 455.1000 1790.7000 455.5800 ;
        RECT 1789.1000 460.5400 1790.7000 461.0200 ;
        RECT 1789.1000 465.9800 1790.7000 466.4600 ;
        RECT 1789.1000 444.2200 1790.7000 444.7000 ;
        RECT 1789.1000 449.6600 1790.7000 450.1400 ;
        RECT 1834.1000 427.9000 1835.7000 428.3800 ;
        RECT 1834.1000 433.3400 1835.7000 433.8200 ;
        RECT 1834.1000 438.7800 1835.7000 439.2600 ;
        RECT 1834.1000 422.4600 1835.7000 422.9400 ;
        RECT 1789.1000 427.9000 1790.7000 428.3800 ;
        RECT 1789.1000 433.3400 1790.7000 433.8200 ;
        RECT 1789.1000 438.7800 1790.7000 439.2600 ;
        RECT 1789.1000 422.4600 1790.7000 422.9400 ;
        RECT 1744.1000 455.1000 1745.7000 455.5800 ;
        RECT 1744.1000 460.5400 1745.7000 461.0200 ;
        RECT 1744.1000 465.9800 1745.7000 466.4600 ;
        RECT 1736.3400 455.1000 1737.9400 455.5800 ;
        RECT 1736.3400 460.5400 1737.9400 461.0200 ;
        RECT 1736.3400 465.9800 1737.9400 466.4600 ;
        RECT 1744.1000 444.2200 1745.7000 444.7000 ;
        RECT 1744.1000 449.6600 1745.7000 450.1400 ;
        RECT 1736.3400 444.2200 1737.9400 444.7000 ;
        RECT 1736.3400 449.6600 1737.9400 450.1400 ;
        RECT 1744.1000 427.9000 1745.7000 428.3800 ;
        RECT 1744.1000 433.3400 1745.7000 433.8200 ;
        RECT 1744.1000 438.7800 1745.7000 439.2600 ;
        RECT 1736.3400 427.9000 1737.9400 428.3800 ;
        RECT 1736.3400 433.3400 1737.9400 433.8200 ;
        RECT 1736.3400 438.7800 1737.9400 439.2600 ;
        RECT 1736.3400 422.4600 1737.9400 422.9400 ;
        RECT 1744.1000 422.4600 1745.7000 422.9400 ;
        RECT 1730.7800 624.7700 1941.0000 626.3700 ;
        RECT 1730.7800 418.2700 1941.0000 419.8700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 412.8400 1737.9400 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1736.3400 630.8800 1737.9400 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 412.8400 1935.4400 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1933.8400 630.8800 1935.4400 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 418.2700 1732.3800 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 418.2700 1941.0000 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1730.7800 624.7700 1732.3800 626.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1939.4000 624.7700 1941.0000 626.3700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'N_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1956.4600 2479.6000 1958.0600 2509.8600 ;
        RECT 2154.1600 2479.6000 2155.7600 2509.8600 ;
      LAYER met3 ;
        RECT 2154.1600 2497.3800 2155.7600 2497.8600 ;
        RECT 1956.4600 2497.3800 1958.0600 2497.8600 ;
        RECT 2154.1600 2491.9400 2155.7600 2492.4200 ;
        RECT 2154.1600 2486.5000 2155.7600 2486.9800 ;
        RECT 1956.4600 2491.9400 1958.0600 2492.4200 ;
        RECT 1956.4600 2486.5000 1958.0600 2486.9800 ;
        RECT 1951.0000 2503.1000 2161.2200 2504.7000 ;
        RECT 1951.0000 2483.5700 2161.2200 2485.1700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.4600 2479.6000 1958.0600 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.4600 2508.2600 1958.0600 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.1600 2479.6000 2155.7600 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.1600 2508.2600 2155.7600 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2483.5700 1952.6000 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2483.5700 2161.2200 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2503.1000 1952.6000 2504.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2503.1000 2161.2200 2504.7000 ;
    END
# end of P/G pin shape extracted from block 'N_term_DSP'


# P/G pin shape extracted from block 'S_term_DSP'
    PORT
      LAYER met4 ;
        RECT 1956.4600 142.9400 1958.0600 173.2000 ;
        RECT 2154.1600 142.9400 2155.7600 173.2000 ;
      LAYER met3 ;
        RECT 2154.1600 160.7200 2155.7600 161.2000 ;
        RECT 1956.4600 160.7200 1958.0600 161.2000 ;
        RECT 2154.1600 155.2800 2155.7600 155.7600 ;
        RECT 2154.1600 149.8400 2155.7600 150.3200 ;
        RECT 1956.4600 155.2800 1958.0600 155.7600 ;
        RECT 1956.4600 149.8400 1958.0600 150.3200 ;
        RECT 1951.0000 166.4400 2161.2200 168.0400 ;
        RECT 1951.0000 146.9100 2161.2200 148.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.4600 142.9400 1958.0600 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.4600 171.6000 1958.0600 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.1600 142.9400 2155.7600 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.1600 171.6000 2155.7600 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 146.9100 1952.6000 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 146.9100 2161.2200 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 166.4400 1952.6000 168.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 166.4400 2161.2200 168.0400 ;
    END
# end of P/G pin shape extracted from block 'S_term_DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1956.5600 2020.3200 1958.1600 2470.1400 ;
        RECT 2154.0600 2020.3200 2155.6600 2470.1400 ;
        RECT 1964.3200 2025.7500 1965.9200 2464.5400 ;
        RECT 2009.3200 2025.7500 2010.9200 2464.5400 ;
        RECT 2054.3200 2025.7500 2055.9200 2464.5400 ;
        RECT 2099.3200 2025.7500 2100.9200 2464.5400 ;
        RECT 2144.3200 2025.7500 2145.9200 2464.5400 ;
      LAYER met3 ;
        RECT 2154.0600 2459.7000 2155.6600 2460.1800 ;
        RECT 2154.0600 2454.2600 2155.6600 2454.7400 ;
        RECT 2154.0600 2448.8200 2155.6600 2449.3000 ;
        RECT 2154.0600 2443.3800 2155.6600 2443.8600 ;
        RECT 2154.0600 2437.9400 2155.6600 2438.4200 ;
        RECT 2154.0600 2432.5000 2155.6600 2432.9800 ;
        RECT 2154.0600 2427.0600 2155.6600 2427.5400 ;
        RECT 2154.0600 2421.6200 2155.6600 2422.1000 ;
        RECT 2154.0600 2416.1800 2155.6600 2416.6600 ;
        RECT 2154.0600 2410.7400 2155.6600 2411.2200 ;
        RECT 2154.0600 2405.3000 2155.6600 2405.7800 ;
        RECT 2154.0600 2399.8600 2155.6600 2400.3400 ;
        RECT 2154.0600 2394.4200 2155.6600 2394.9000 ;
        RECT 2154.0600 2388.9800 2155.6600 2389.4600 ;
        RECT 2154.0600 2383.5400 2155.6600 2384.0200 ;
        RECT 2154.0600 2378.1000 2155.6600 2378.5800 ;
        RECT 2154.0600 2372.6600 2155.6600 2373.1400 ;
        RECT 2154.0600 2367.2200 2155.6600 2367.7000 ;
        RECT 2154.0600 2361.7800 2155.6600 2362.2600 ;
        RECT 2154.0600 2356.3400 2155.6600 2356.8200 ;
        RECT 2154.0600 2350.9000 2155.6600 2351.3800 ;
        RECT 2154.0600 2345.4600 2155.6600 2345.9400 ;
        RECT 2154.0600 2340.0200 2155.6600 2340.5000 ;
        RECT 2154.0600 2334.5800 2155.6600 2335.0600 ;
        RECT 2154.0600 2323.7000 2155.6600 2324.1800 ;
        RECT 2154.0600 2318.2600 2155.6600 2318.7400 ;
        RECT 2154.0600 2312.8200 2155.6600 2313.3000 ;
        RECT 2154.0600 2307.3800 2155.6600 2307.8600 ;
        RECT 2154.0600 2301.9400 2155.6600 2302.4200 ;
        RECT 2154.0600 2329.1400 2155.6600 2329.6200 ;
        RECT 2154.0600 2296.5000 2155.6600 2296.9800 ;
        RECT 2154.0600 2291.0600 2155.6600 2291.5400 ;
        RECT 2154.0600 2285.6200 2155.6600 2286.1000 ;
        RECT 2154.0600 2280.1800 2155.6600 2280.6600 ;
        RECT 2154.0600 2274.7400 2155.6600 2275.2200 ;
        RECT 2154.0600 2269.3000 2155.6600 2269.7800 ;
        RECT 2154.0600 2263.8600 2155.6600 2264.3400 ;
        RECT 2154.0600 2258.4200 2155.6600 2258.9000 ;
        RECT 2154.0600 2252.9800 2155.6600 2253.4600 ;
        RECT 2154.0600 2247.5400 2155.6600 2248.0200 ;
        RECT 1956.5600 2459.7000 1958.1600 2460.1800 ;
        RECT 1956.5600 2454.2600 1958.1600 2454.7400 ;
        RECT 1956.5600 2448.8200 1958.1600 2449.3000 ;
        RECT 1956.5600 2443.3800 1958.1600 2443.8600 ;
        RECT 1956.5600 2437.9400 1958.1600 2438.4200 ;
        RECT 1956.5600 2432.5000 1958.1600 2432.9800 ;
        RECT 1956.5600 2427.0600 1958.1600 2427.5400 ;
        RECT 1956.5600 2421.6200 1958.1600 2422.1000 ;
        RECT 1956.5600 2416.1800 1958.1600 2416.6600 ;
        RECT 1956.5600 2410.7400 1958.1600 2411.2200 ;
        RECT 1956.5600 2405.3000 1958.1600 2405.7800 ;
        RECT 1956.5600 2399.8600 1958.1600 2400.3400 ;
        RECT 1956.5600 2394.4200 1958.1600 2394.9000 ;
        RECT 1956.5600 2388.9800 1958.1600 2389.4600 ;
        RECT 1956.5600 2383.5400 1958.1600 2384.0200 ;
        RECT 1956.5600 2378.1000 1958.1600 2378.5800 ;
        RECT 1956.5600 2372.6600 1958.1600 2373.1400 ;
        RECT 1956.5600 2367.2200 1958.1600 2367.7000 ;
        RECT 1956.5600 2361.7800 1958.1600 2362.2600 ;
        RECT 1956.5600 2356.3400 1958.1600 2356.8200 ;
        RECT 1956.5600 2350.9000 1958.1600 2351.3800 ;
        RECT 1956.5600 2345.4600 1958.1600 2345.9400 ;
        RECT 1956.5600 2340.0200 1958.1600 2340.5000 ;
        RECT 1956.5600 2334.5800 1958.1600 2335.0600 ;
        RECT 1956.5600 2323.7000 1958.1600 2324.1800 ;
        RECT 1956.5600 2318.2600 1958.1600 2318.7400 ;
        RECT 1956.5600 2312.8200 1958.1600 2313.3000 ;
        RECT 1956.5600 2307.3800 1958.1600 2307.8600 ;
        RECT 1956.5600 2301.9400 1958.1600 2302.4200 ;
        RECT 1956.5600 2329.1400 1958.1600 2329.6200 ;
        RECT 1956.5600 2296.5000 1958.1600 2296.9800 ;
        RECT 1956.5600 2291.0600 1958.1600 2291.5400 ;
        RECT 1956.5600 2285.6200 1958.1600 2286.1000 ;
        RECT 1956.5600 2280.1800 1958.1600 2280.6600 ;
        RECT 1956.5600 2274.7400 1958.1600 2275.2200 ;
        RECT 1956.5600 2269.3000 1958.1600 2269.7800 ;
        RECT 1956.5600 2263.8600 1958.1600 2264.3400 ;
        RECT 1956.5600 2258.4200 1958.1600 2258.9000 ;
        RECT 1956.5600 2252.9800 1958.1600 2253.4600 ;
        RECT 1956.5600 2247.5400 1958.1600 2248.0200 ;
        RECT 2154.0600 2242.1000 2155.6600 2242.5800 ;
        RECT 2154.0600 2236.6600 2155.6600 2237.1400 ;
        RECT 2154.0600 2231.2200 2155.6600 2231.7000 ;
        RECT 2154.0600 2225.7800 2155.6600 2226.2600 ;
        RECT 2154.0600 2220.3400 2155.6600 2220.8200 ;
        RECT 2154.0600 2214.9000 2155.6600 2215.3800 ;
        RECT 2154.0600 2209.4600 2155.6600 2209.9400 ;
        RECT 2154.0600 2204.0200 2155.6600 2204.5000 ;
        RECT 2154.0600 2198.5800 2155.6600 2199.0600 ;
        RECT 2154.0600 2193.1400 2155.6600 2193.6200 ;
        RECT 2154.0600 2187.7000 2155.6600 2188.1800 ;
        RECT 2154.0600 2182.2600 2155.6600 2182.7400 ;
        RECT 2154.0600 2176.8200 2155.6600 2177.3000 ;
        RECT 2154.0600 2171.3800 2155.6600 2171.8600 ;
        RECT 2154.0600 2165.9400 2155.6600 2166.4200 ;
        RECT 2154.0600 2155.0600 2155.6600 2155.5400 ;
        RECT 2154.0600 2149.6200 2155.6600 2150.1000 ;
        RECT 2154.0600 2144.1800 2155.6600 2144.6600 ;
        RECT 2154.0600 2138.7400 2155.6600 2139.2200 ;
        RECT 2154.0600 2133.3000 2155.6600 2133.7800 ;
        RECT 2154.0600 2160.5000 2155.6600 2160.9800 ;
        RECT 2154.0600 2127.8600 2155.6600 2128.3400 ;
        RECT 2154.0600 2122.4200 2155.6600 2122.9000 ;
        RECT 2154.0600 2116.9800 2155.6600 2117.4600 ;
        RECT 2154.0600 2111.5400 2155.6600 2112.0200 ;
        RECT 2154.0600 2106.1000 2155.6600 2106.5800 ;
        RECT 2154.0600 2100.6600 2155.6600 2101.1400 ;
        RECT 2154.0600 2095.2200 2155.6600 2095.7000 ;
        RECT 2154.0600 2089.7800 2155.6600 2090.2600 ;
        RECT 2154.0600 2084.3400 2155.6600 2084.8200 ;
        RECT 2154.0600 2078.9000 2155.6600 2079.3800 ;
        RECT 2154.0600 2073.4600 2155.6600 2073.9400 ;
        RECT 2154.0600 2068.0200 2155.6600 2068.5000 ;
        RECT 2154.0600 2062.5800 2155.6600 2063.0600 ;
        RECT 2154.0600 2057.1400 2155.6600 2057.6200 ;
        RECT 2154.0600 2051.7000 2155.6600 2052.1800 ;
        RECT 2154.0600 2046.2600 2155.6600 2046.7400 ;
        RECT 2154.0600 2040.8200 2155.6600 2041.3000 ;
        RECT 2154.0600 2035.3800 2155.6600 2035.8600 ;
        RECT 2154.0600 2029.9400 2155.6600 2030.4200 ;
        RECT 1956.5600 2242.1000 1958.1600 2242.5800 ;
        RECT 1956.5600 2236.6600 1958.1600 2237.1400 ;
        RECT 1956.5600 2231.2200 1958.1600 2231.7000 ;
        RECT 1956.5600 2225.7800 1958.1600 2226.2600 ;
        RECT 1956.5600 2220.3400 1958.1600 2220.8200 ;
        RECT 1956.5600 2214.9000 1958.1600 2215.3800 ;
        RECT 1956.5600 2209.4600 1958.1600 2209.9400 ;
        RECT 1956.5600 2204.0200 1958.1600 2204.5000 ;
        RECT 1956.5600 2198.5800 1958.1600 2199.0600 ;
        RECT 1956.5600 2193.1400 1958.1600 2193.6200 ;
        RECT 1956.5600 2187.7000 1958.1600 2188.1800 ;
        RECT 1956.5600 2182.2600 1958.1600 2182.7400 ;
        RECT 1956.5600 2176.8200 1958.1600 2177.3000 ;
        RECT 1956.5600 2171.3800 1958.1600 2171.8600 ;
        RECT 1956.5600 2165.9400 1958.1600 2166.4200 ;
        RECT 1956.5600 2155.0600 1958.1600 2155.5400 ;
        RECT 1956.5600 2149.6200 1958.1600 2150.1000 ;
        RECT 1956.5600 2144.1800 1958.1600 2144.6600 ;
        RECT 1956.5600 2138.7400 1958.1600 2139.2200 ;
        RECT 1956.5600 2133.3000 1958.1600 2133.7800 ;
        RECT 1956.5600 2160.5000 1958.1600 2160.9800 ;
        RECT 1956.5600 2127.8600 1958.1600 2128.3400 ;
        RECT 1956.5600 2122.4200 1958.1600 2122.9000 ;
        RECT 1956.5600 2116.9800 1958.1600 2117.4600 ;
        RECT 1956.5600 2111.5400 1958.1600 2112.0200 ;
        RECT 1956.5600 2106.1000 1958.1600 2106.5800 ;
        RECT 1956.5600 2100.6600 1958.1600 2101.1400 ;
        RECT 1956.5600 2095.2200 1958.1600 2095.7000 ;
        RECT 1956.5600 2089.7800 1958.1600 2090.2600 ;
        RECT 1956.5600 2084.3400 1958.1600 2084.8200 ;
        RECT 1956.5600 2078.9000 1958.1600 2079.3800 ;
        RECT 1956.5600 2073.4600 1958.1600 2073.9400 ;
        RECT 1956.5600 2068.0200 1958.1600 2068.5000 ;
        RECT 1956.5600 2062.5800 1958.1600 2063.0600 ;
        RECT 1956.5600 2057.1400 1958.1600 2057.6200 ;
        RECT 1956.5600 2051.7000 1958.1600 2052.1800 ;
        RECT 1956.5600 2046.2600 1958.1600 2046.7400 ;
        RECT 1956.5600 2040.8200 1958.1600 2041.3000 ;
        RECT 1956.5600 2035.3800 1958.1600 2035.8600 ;
        RECT 1956.5600 2029.9400 1958.1600 2030.4200 ;
        RECT 1951.0000 2462.9400 2161.2200 2464.5400 ;
        RECT 1951.0000 2025.7500 2161.2200 2027.3500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 2020.3200 1958.1600 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 2468.5400 1958.1600 2470.1400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 2020.3200 2155.6600 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 2468.5400 2155.6600 2470.1400 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2025.7500 1952.6000 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2025.7500 2161.2200 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2462.9400 1952.6000 2464.5400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2462.9400 2161.2200 2464.5400 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1956.5600 1561.0400 1958.1600 2010.8600 ;
        RECT 2154.0600 1561.0400 2155.6600 2010.8600 ;
        RECT 1964.3200 1566.4700 1965.9200 2005.2600 ;
        RECT 2009.3200 1566.4700 2010.9200 2005.2600 ;
        RECT 2054.3200 1566.4700 2055.9200 2005.2600 ;
        RECT 2099.3200 1566.4700 2100.9200 2005.2600 ;
        RECT 2144.3200 1566.4700 2145.9200 2005.2600 ;
      LAYER met3 ;
        RECT 2154.0600 2000.4200 2155.6600 2000.9000 ;
        RECT 2154.0600 1994.9800 2155.6600 1995.4600 ;
        RECT 2154.0600 1989.5400 2155.6600 1990.0200 ;
        RECT 2154.0600 1984.1000 2155.6600 1984.5800 ;
        RECT 2154.0600 1978.6600 2155.6600 1979.1400 ;
        RECT 2154.0600 1973.2200 2155.6600 1973.7000 ;
        RECT 2154.0600 1967.7800 2155.6600 1968.2600 ;
        RECT 2154.0600 1962.3400 2155.6600 1962.8200 ;
        RECT 2154.0600 1956.9000 2155.6600 1957.3800 ;
        RECT 2154.0600 1951.4600 2155.6600 1951.9400 ;
        RECT 2154.0600 1946.0200 2155.6600 1946.5000 ;
        RECT 2154.0600 1940.5800 2155.6600 1941.0600 ;
        RECT 2154.0600 1935.1400 2155.6600 1935.6200 ;
        RECT 2154.0600 1929.7000 2155.6600 1930.1800 ;
        RECT 2154.0600 1924.2600 2155.6600 1924.7400 ;
        RECT 2154.0600 1918.8200 2155.6600 1919.3000 ;
        RECT 2154.0600 1913.3800 2155.6600 1913.8600 ;
        RECT 2154.0600 1907.9400 2155.6600 1908.4200 ;
        RECT 2154.0600 1902.5000 2155.6600 1902.9800 ;
        RECT 2154.0600 1897.0600 2155.6600 1897.5400 ;
        RECT 2154.0600 1891.6200 2155.6600 1892.1000 ;
        RECT 2154.0600 1886.1800 2155.6600 1886.6600 ;
        RECT 2154.0600 1880.7400 2155.6600 1881.2200 ;
        RECT 2154.0600 1875.3000 2155.6600 1875.7800 ;
        RECT 2154.0600 1864.4200 2155.6600 1864.9000 ;
        RECT 2154.0600 1858.9800 2155.6600 1859.4600 ;
        RECT 2154.0600 1853.5400 2155.6600 1854.0200 ;
        RECT 2154.0600 1848.1000 2155.6600 1848.5800 ;
        RECT 2154.0600 1842.6600 2155.6600 1843.1400 ;
        RECT 2154.0600 1869.8600 2155.6600 1870.3400 ;
        RECT 2154.0600 1837.2200 2155.6600 1837.7000 ;
        RECT 2154.0600 1831.7800 2155.6600 1832.2600 ;
        RECT 2154.0600 1826.3400 2155.6600 1826.8200 ;
        RECT 2154.0600 1820.9000 2155.6600 1821.3800 ;
        RECT 2154.0600 1815.4600 2155.6600 1815.9400 ;
        RECT 2154.0600 1810.0200 2155.6600 1810.5000 ;
        RECT 2154.0600 1804.5800 2155.6600 1805.0600 ;
        RECT 2154.0600 1799.1400 2155.6600 1799.6200 ;
        RECT 2154.0600 1793.7000 2155.6600 1794.1800 ;
        RECT 2154.0600 1788.2600 2155.6600 1788.7400 ;
        RECT 1956.5600 2000.4200 1958.1600 2000.9000 ;
        RECT 1956.5600 1994.9800 1958.1600 1995.4600 ;
        RECT 1956.5600 1989.5400 1958.1600 1990.0200 ;
        RECT 1956.5600 1984.1000 1958.1600 1984.5800 ;
        RECT 1956.5600 1978.6600 1958.1600 1979.1400 ;
        RECT 1956.5600 1973.2200 1958.1600 1973.7000 ;
        RECT 1956.5600 1967.7800 1958.1600 1968.2600 ;
        RECT 1956.5600 1962.3400 1958.1600 1962.8200 ;
        RECT 1956.5600 1956.9000 1958.1600 1957.3800 ;
        RECT 1956.5600 1951.4600 1958.1600 1951.9400 ;
        RECT 1956.5600 1946.0200 1958.1600 1946.5000 ;
        RECT 1956.5600 1940.5800 1958.1600 1941.0600 ;
        RECT 1956.5600 1935.1400 1958.1600 1935.6200 ;
        RECT 1956.5600 1929.7000 1958.1600 1930.1800 ;
        RECT 1956.5600 1924.2600 1958.1600 1924.7400 ;
        RECT 1956.5600 1918.8200 1958.1600 1919.3000 ;
        RECT 1956.5600 1913.3800 1958.1600 1913.8600 ;
        RECT 1956.5600 1907.9400 1958.1600 1908.4200 ;
        RECT 1956.5600 1902.5000 1958.1600 1902.9800 ;
        RECT 1956.5600 1897.0600 1958.1600 1897.5400 ;
        RECT 1956.5600 1891.6200 1958.1600 1892.1000 ;
        RECT 1956.5600 1886.1800 1958.1600 1886.6600 ;
        RECT 1956.5600 1880.7400 1958.1600 1881.2200 ;
        RECT 1956.5600 1875.3000 1958.1600 1875.7800 ;
        RECT 1956.5600 1864.4200 1958.1600 1864.9000 ;
        RECT 1956.5600 1858.9800 1958.1600 1859.4600 ;
        RECT 1956.5600 1853.5400 1958.1600 1854.0200 ;
        RECT 1956.5600 1848.1000 1958.1600 1848.5800 ;
        RECT 1956.5600 1842.6600 1958.1600 1843.1400 ;
        RECT 1956.5600 1869.8600 1958.1600 1870.3400 ;
        RECT 1956.5600 1837.2200 1958.1600 1837.7000 ;
        RECT 1956.5600 1831.7800 1958.1600 1832.2600 ;
        RECT 1956.5600 1826.3400 1958.1600 1826.8200 ;
        RECT 1956.5600 1820.9000 1958.1600 1821.3800 ;
        RECT 1956.5600 1815.4600 1958.1600 1815.9400 ;
        RECT 1956.5600 1810.0200 1958.1600 1810.5000 ;
        RECT 1956.5600 1804.5800 1958.1600 1805.0600 ;
        RECT 1956.5600 1799.1400 1958.1600 1799.6200 ;
        RECT 1956.5600 1793.7000 1958.1600 1794.1800 ;
        RECT 1956.5600 1788.2600 1958.1600 1788.7400 ;
        RECT 2154.0600 1782.8200 2155.6600 1783.3000 ;
        RECT 2154.0600 1777.3800 2155.6600 1777.8600 ;
        RECT 2154.0600 1771.9400 2155.6600 1772.4200 ;
        RECT 2154.0600 1766.5000 2155.6600 1766.9800 ;
        RECT 2154.0600 1761.0600 2155.6600 1761.5400 ;
        RECT 2154.0600 1755.6200 2155.6600 1756.1000 ;
        RECT 2154.0600 1750.1800 2155.6600 1750.6600 ;
        RECT 2154.0600 1744.7400 2155.6600 1745.2200 ;
        RECT 2154.0600 1739.3000 2155.6600 1739.7800 ;
        RECT 2154.0600 1733.8600 2155.6600 1734.3400 ;
        RECT 2154.0600 1728.4200 2155.6600 1728.9000 ;
        RECT 2154.0600 1722.9800 2155.6600 1723.4600 ;
        RECT 2154.0600 1717.5400 2155.6600 1718.0200 ;
        RECT 2154.0600 1712.1000 2155.6600 1712.5800 ;
        RECT 2154.0600 1706.6600 2155.6600 1707.1400 ;
        RECT 2154.0600 1695.7800 2155.6600 1696.2600 ;
        RECT 2154.0600 1690.3400 2155.6600 1690.8200 ;
        RECT 2154.0600 1684.9000 2155.6600 1685.3800 ;
        RECT 2154.0600 1679.4600 2155.6600 1679.9400 ;
        RECT 2154.0600 1674.0200 2155.6600 1674.5000 ;
        RECT 2154.0600 1701.2200 2155.6600 1701.7000 ;
        RECT 2154.0600 1668.5800 2155.6600 1669.0600 ;
        RECT 2154.0600 1663.1400 2155.6600 1663.6200 ;
        RECT 2154.0600 1657.7000 2155.6600 1658.1800 ;
        RECT 2154.0600 1652.2600 2155.6600 1652.7400 ;
        RECT 2154.0600 1646.8200 2155.6600 1647.3000 ;
        RECT 2154.0600 1641.3800 2155.6600 1641.8600 ;
        RECT 2154.0600 1635.9400 2155.6600 1636.4200 ;
        RECT 2154.0600 1630.5000 2155.6600 1630.9800 ;
        RECT 2154.0600 1625.0600 2155.6600 1625.5400 ;
        RECT 2154.0600 1619.6200 2155.6600 1620.1000 ;
        RECT 2154.0600 1614.1800 2155.6600 1614.6600 ;
        RECT 2154.0600 1608.7400 2155.6600 1609.2200 ;
        RECT 2154.0600 1603.3000 2155.6600 1603.7800 ;
        RECT 2154.0600 1597.8600 2155.6600 1598.3400 ;
        RECT 2154.0600 1592.4200 2155.6600 1592.9000 ;
        RECT 2154.0600 1586.9800 2155.6600 1587.4600 ;
        RECT 2154.0600 1581.5400 2155.6600 1582.0200 ;
        RECT 2154.0600 1576.1000 2155.6600 1576.5800 ;
        RECT 2154.0600 1570.6600 2155.6600 1571.1400 ;
        RECT 1956.5600 1782.8200 1958.1600 1783.3000 ;
        RECT 1956.5600 1777.3800 1958.1600 1777.8600 ;
        RECT 1956.5600 1771.9400 1958.1600 1772.4200 ;
        RECT 1956.5600 1766.5000 1958.1600 1766.9800 ;
        RECT 1956.5600 1761.0600 1958.1600 1761.5400 ;
        RECT 1956.5600 1755.6200 1958.1600 1756.1000 ;
        RECT 1956.5600 1750.1800 1958.1600 1750.6600 ;
        RECT 1956.5600 1744.7400 1958.1600 1745.2200 ;
        RECT 1956.5600 1739.3000 1958.1600 1739.7800 ;
        RECT 1956.5600 1733.8600 1958.1600 1734.3400 ;
        RECT 1956.5600 1728.4200 1958.1600 1728.9000 ;
        RECT 1956.5600 1722.9800 1958.1600 1723.4600 ;
        RECT 1956.5600 1717.5400 1958.1600 1718.0200 ;
        RECT 1956.5600 1712.1000 1958.1600 1712.5800 ;
        RECT 1956.5600 1706.6600 1958.1600 1707.1400 ;
        RECT 1956.5600 1695.7800 1958.1600 1696.2600 ;
        RECT 1956.5600 1690.3400 1958.1600 1690.8200 ;
        RECT 1956.5600 1684.9000 1958.1600 1685.3800 ;
        RECT 1956.5600 1679.4600 1958.1600 1679.9400 ;
        RECT 1956.5600 1674.0200 1958.1600 1674.5000 ;
        RECT 1956.5600 1701.2200 1958.1600 1701.7000 ;
        RECT 1956.5600 1668.5800 1958.1600 1669.0600 ;
        RECT 1956.5600 1663.1400 1958.1600 1663.6200 ;
        RECT 1956.5600 1657.7000 1958.1600 1658.1800 ;
        RECT 1956.5600 1652.2600 1958.1600 1652.7400 ;
        RECT 1956.5600 1646.8200 1958.1600 1647.3000 ;
        RECT 1956.5600 1641.3800 1958.1600 1641.8600 ;
        RECT 1956.5600 1635.9400 1958.1600 1636.4200 ;
        RECT 1956.5600 1630.5000 1958.1600 1630.9800 ;
        RECT 1956.5600 1625.0600 1958.1600 1625.5400 ;
        RECT 1956.5600 1619.6200 1958.1600 1620.1000 ;
        RECT 1956.5600 1614.1800 1958.1600 1614.6600 ;
        RECT 1956.5600 1608.7400 1958.1600 1609.2200 ;
        RECT 1956.5600 1603.3000 1958.1600 1603.7800 ;
        RECT 1956.5600 1597.8600 1958.1600 1598.3400 ;
        RECT 1956.5600 1592.4200 1958.1600 1592.9000 ;
        RECT 1956.5600 1586.9800 1958.1600 1587.4600 ;
        RECT 1956.5600 1581.5400 1958.1600 1582.0200 ;
        RECT 1956.5600 1576.1000 1958.1600 1576.5800 ;
        RECT 1956.5600 1570.6600 1958.1600 1571.1400 ;
        RECT 1951.0000 2003.6600 2161.2200 2005.2600 ;
        RECT 1951.0000 1566.4700 2161.2200 1568.0700 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 1561.0400 1958.1600 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 2009.2600 1958.1600 2010.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 1561.0400 2155.6600 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 2009.2600 2155.6600 2010.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1566.4700 1952.6000 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1566.4700 2161.2200 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 2003.6600 1952.6000 2005.2600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 2003.6600 2161.2200 2005.2600 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1956.5600 1101.7600 1958.1600 1551.5800 ;
        RECT 2154.0600 1101.7600 2155.6600 1551.5800 ;
        RECT 1964.3200 1107.1900 1965.9200 1545.9800 ;
        RECT 2009.3200 1107.1900 2010.9200 1545.9800 ;
        RECT 2054.3200 1107.1900 2055.9200 1545.9800 ;
        RECT 2099.3200 1107.1900 2100.9200 1545.9800 ;
        RECT 2144.3200 1107.1900 2145.9200 1545.9800 ;
      LAYER met3 ;
        RECT 2154.0600 1541.1400 2155.6600 1541.6200 ;
        RECT 2154.0600 1535.7000 2155.6600 1536.1800 ;
        RECT 2154.0600 1530.2600 2155.6600 1530.7400 ;
        RECT 2154.0600 1524.8200 2155.6600 1525.3000 ;
        RECT 2154.0600 1519.3800 2155.6600 1519.8600 ;
        RECT 2154.0600 1513.9400 2155.6600 1514.4200 ;
        RECT 2154.0600 1508.5000 2155.6600 1508.9800 ;
        RECT 2154.0600 1503.0600 2155.6600 1503.5400 ;
        RECT 2154.0600 1497.6200 2155.6600 1498.1000 ;
        RECT 2154.0600 1492.1800 2155.6600 1492.6600 ;
        RECT 2154.0600 1486.7400 2155.6600 1487.2200 ;
        RECT 2154.0600 1481.3000 2155.6600 1481.7800 ;
        RECT 2154.0600 1475.8600 2155.6600 1476.3400 ;
        RECT 2154.0600 1470.4200 2155.6600 1470.9000 ;
        RECT 2154.0600 1464.9800 2155.6600 1465.4600 ;
        RECT 2154.0600 1459.5400 2155.6600 1460.0200 ;
        RECT 2154.0600 1454.1000 2155.6600 1454.5800 ;
        RECT 2154.0600 1448.6600 2155.6600 1449.1400 ;
        RECT 2154.0600 1443.2200 2155.6600 1443.7000 ;
        RECT 2154.0600 1437.7800 2155.6600 1438.2600 ;
        RECT 2154.0600 1432.3400 2155.6600 1432.8200 ;
        RECT 2154.0600 1426.9000 2155.6600 1427.3800 ;
        RECT 2154.0600 1421.4600 2155.6600 1421.9400 ;
        RECT 2154.0600 1416.0200 2155.6600 1416.5000 ;
        RECT 2154.0600 1405.1400 2155.6600 1405.6200 ;
        RECT 2154.0600 1399.7000 2155.6600 1400.1800 ;
        RECT 2154.0600 1394.2600 2155.6600 1394.7400 ;
        RECT 2154.0600 1388.8200 2155.6600 1389.3000 ;
        RECT 2154.0600 1383.3800 2155.6600 1383.8600 ;
        RECT 2154.0600 1410.5800 2155.6600 1411.0600 ;
        RECT 2154.0600 1377.9400 2155.6600 1378.4200 ;
        RECT 2154.0600 1372.5000 2155.6600 1372.9800 ;
        RECT 2154.0600 1367.0600 2155.6600 1367.5400 ;
        RECT 2154.0600 1361.6200 2155.6600 1362.1000 ;
        RECT 2154.0600 1356.1800 2155.6600 1356.6600 ;
        RECT 2154.0600 1350.7400 2155.6600 1351.2200 ;
        RECT 2154.0600 1345.3000 2155.6600 1345.7800 ;
        RECT 2154.0600 1339.8600 2155.6600 1340.3400 ;
        RECT 2154.0600 1334.4200 2155.6600 1334.9000 ;
        RECT 2154.0600 1328.9800 2155.6600 1329.4600 ;
        RECT 1956.5600 1541.1400 1958.1600 1541.6200 ;
        RECT 1956.5600 1535.7000 1958.1600 1536.1800 ;
        RECT 1956.5600 1530.2600 1958.1600 1530.7400 ;
        RECT 1956.5600 1524.8200 1958.1600 1525.3000 ;
        RECT 1956.5600 1519.3800 1958.1600 1519.8600 ;
        RECT 1956.5600 1513.9400 1958.1600 1514.4200 ;
        RECT 1956.5600 1508.5000 1958.1600 1508.9800 ;
        RECT 1956.5600 1503.0600 1958.1600 1503.5400 ;
        RECT 1956.5600 1497.6200 1958.1600 1498.1000 ;
        RECT 1956.5600 1492.1800 1958.1600 1492.6600 ;
        RECT 1956.5600 1486.7400 1958.1600 1487.2200 ;
        RECT 1956.5600 1481.3000 1958.1600 1481.7800 ;
        RECT 1956.5600 1475.8600 1958.1600 1476.3400 ;
        RECT 1956.5600 1470.4200 1958.1600 1470.9000 ;
        RECT 1956.5600 1464.9800 1958.1600 1465.4600 ;
        RECT 1956.5600 1459.5400 1958.1600 1460.0200 ;
        RECT 1956.5600 1454.1000 1958.1600 1454.5800 ;
        RECT 1956.5600 1448.6600 1958.1600 1449.1400 ;
        RECT 1956.5600 1443.2200 1958.1600 1443.7000 ;
        RECT 1956.5600 1437.7800 1958.1600 1438.2600 ;
        RECT 1956.5600 1432.3400 1958.1600 1432.8200 ;
        RECT 1956.5600 1426.9000 1958.1600 1427.3800 ;
        RECT 1956.5600 1421.4600 1958.1600 1421.9400 ;
        RECT 1956.5600 1416.0200 1958.1600 1416.5000 ;
        RECT 1956.5600 1405.1400 1958.1600 1405.6200 ;
        RECT 1956.5600 1399.7000 1958.1600 1400.1800 ;
        RECT 1956.5600 1394.2600 1958.1600 1394.7400 ;
        RECT 1956.5600 1388.8200 1958.1600 1389.3000 ;
        RECT 1956.5600 1383.3800 1958.1600 1383.8600 ;
        RECT 1956.5600 1410.5800 1958.1600 1411.0600 ;
        RECT 1956.5600 1377.9400 1958.1600 1378.4200 ;
        RECT 1956.5600 1372.5000 1958.1600 1372.9800 ;
        RECT 1956.5600 1367.0600 1958.1600 1367.5400 ;
        RECT 1956.5600 1361.6200 1958.1600 1362.1000 ;
        RECT 1956.5600 1356.1800 1958.1600 1356.6600 ;
        RECT 1956.5600 1350.7400 1958.1600 1351.2200 ;
        RECT 1956.5600 1345.3000 1958.1600 1345.7800 ;
        RECT 1956.5600 1339.8600 1958.1600 1340.3400 ;
        RECT 1956.5600 1334.4200 1958.1600 1334.9000 ;
        RECT 1956.5600 1328.9800 1958.1600 1329.4600 ;
        RECT 2154.0600 1323.5400 2155.6600 1324.0200 ;
        RECT 2154.0600 1318.1000 2155.6600 1318.5800 ;
        RECT 2154.0600 1312.6600 2155.6600 1313.1400 ;
        RECT 2154.0600 1307.2200 2155.6600 1307.7000 ;
        RECT 2154.0600 1301.7800 2155.6600 1302.2600 ;
        RECT 2154.0600 1296.3400 2155.6600 1296.8200 ;
        RECT 2154.0600 1290.9000 2155.6600 1291.3800 ;
        RECT 2154.0600 1285.4600 2155.6600 1285.9400 ;
        RECT 2154.0600 1280.0200 2155.6600 1280.5000 ;
        RECT 2154.0600 1274.5800 2155.6600 1275.0600 ;
        RECT 2154.0600 1269.1400 2155.6600 1269.6200 ;
        RECT 2154.0600 1263.7000 2155.6600 1264.1800 ;
        RECT 2154.0600 1258.2600 2155.6600 1258.7400 ;
        RECT 2154.0600 1252.8200 2155.6600 1253.3000 ;
        RECT 2154.0600 1247.3800 2155.6600 1247.8600 ;
        RECT 2154.0600 1236.5000 2155.6600 1236.9800 ;
        RECT 2154.0600 1231.0600 2155.6600 1231.5400 ;
        RECT 2154.0600 1225.6200 2155.6600 1226.1000 ;
        RECT 2154.0600 1220.1800 2155.6600 1220.6600 ;
        RECT 2154.0600 1214.7400 2155.6600 1215.2200 ;
        RECT 2154.0600 1241.9400 2155.6600 1242.4200 ;
        RECT 2154.0600 1209.3000 2155.6600 1209.7800 ;
        RECT 2154.0600 1203.8600 2155.6600 1204.3400 ;
        RECT 2154.0600 1198.4200 2155.6600 1198.9000 ;
        RECT 2154.0600 1192.9800 2155.6600 1193.4600 ;
        RECT 2154.0600 1187.5400 2155.6600 1188.0200 ;
        RECT 2154.0600 1182.1000 2155.6600 1182.5800 ;
        RECT 2154.0600 1176.6600 2155.6600 1177.1400 ;
        RECT 2154.0600 1171.2200 2155.6600 1171.7000 ;
        RECT 2154.0600 1165.7800 2155.6600 1166.2600 ;
        RECT 2154.0600 1160.3400 2155.6600 1160.8200 ;
        RECT 2154.0600 1154.9000 2155.6600 1155.3800 ;
        RECT 2154.0600 1149.4600 2155.6600 1149.9400 ;
        RECT 2154.0600 1144.0200 2155.6600 1144.5000 ;
        RECT 2154.0600 1138.5800 2155.6600 1139.0600 ;
        RECT 2154.0600 1133.1400 2155.6600 1133.6200 ;
        RECT 2154.0600 1127.7000 2155.6600 1128.1800 ;
        RECT 2154.0600 1122.2600 2155.6600 1122.7400 ;
        RECT 2154.0600 1116.8200 2155.6600 1117.3000 ;
        RECT 2154.0600 1111.3800 2155.6600 1111.8600 ;
        RECT 1956.5600 1323.5400 1958.1600 1324.0200 ;
        RECT 1956.5600 1318.1000 1958.1600 1318.5800 ;
        RECT 1956.5600 1312.6600 1958.1600 1313.1400 ;
        RECT 1956.5600 1307.2200 1958.1600 1307.7000 ;
        RECT 1956.5600 1301.7800 1958.1600 1302.2600 ;
        RECT 1956.5600 1296.3400 1958.1600 1296.8200 ;
        RECT 1956.5600 1290.9000 1958.1600 1291.3800 ;
        RECT 1956.5600 1285.4600 1958.1600 1285.9400 ;
        RECT 1956.5600 1280.0200 1958.1600 1280.5000 ;
        RECT 1956.5600 1274.5800 1958.1600 1275.0600 ;
        RECT 1956.5600 1269.1400 1958.1600 1269.6200 ;
        RECT 1956.5600 1263.7000 1958.1600 1264.1800 ;
        RECT 1956.5600 1258.2600 1958.1600 1258.7400 ;
        RECT 1956.5600 1252.8200 1958.1600 1253.3000 ;
        RECT 1956.5600 1247.3800 1958.1600 1247.8600 ;
        RECT 1956.5600 1236.5000 1958.1600 1236.9800 ;
        RECT 1956.5600 1231.0600 1958.1600 1231.5400 ;
        RECT 1956.5600 1225.6200 1958.1600 1226.1000 ;
        RECT 1956.5600 1220.1800 1958.1600 1220.6600 ;
        RECT 1956.5600 1214.7400 1958.1600 1215.2200 ;
        RECT 1956.5600 1241.9400 1958.1600 1242.4200 ;
        RECT 1956.5600 1209.3000 1958.1600 1209.7800 ;
        RECT 1956.5600 1203.8600 1958.1600 1204.3400 ;
        RECT 1956.5600 1198.4200 1958.1600 1198.9000 ;
        RECT 1956.5600 1192.9800 1958.1600 1193.4600 ;
        RECT 1956.5600 1187.5400 1958.1600 1188.0200 ;
        RECT 1956.5600 1182.1000 1958.1600 1182.5800 ;
        RECT 1956.5600 1176.6600 1958.1600 1177.1400 ;
        RECT 1956.5600 1171.2200 1958.1600 1171.7000 ;
        RECT 1956.5600 1165.7800 1958.1600 1166.2600 ;
        RECT 1956.5600 1160.3400 1958.1600 1160.8200 ;
        RECT 1956.5600 1154.9000 1958.1600 1155.3800 ;
        RECT 1956.5600 1149.4600 1958.1600 1149.9400 ;
        RECT 1956.5600 1144.0200 1958.1600 1144.5000 ;
        RECT 1956.5600 1138.5800 1958.1600 1139.0600 ;
        RECT 1956.5600 1133.1400 1958.1600 1133.6200 ;
        RECT 1956.5600 1127.7000 1958.1600 1128.1800 ;
        RECT 1956.5600 1122.2600 1958.1600 1122.7400 ;
        RECT 1956.5600 1116.8200 1958.1600 1117.3000 ;
        RECT 1956.5600 1111.3800 1958.1600 1111.8600 ;
        RECT 1951.0000 1544.3800 2161.2200 1545.9800 ;
        RECT 1951.0000 1107.1900 2161.2200 1108.7900 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 1101.7600 1958.1600 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 1549.9800 1958.1600 1551.5800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 1101.7600 2155.6600 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 1549.9800 2155.6600 1551.5800 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1107.1900 1952.6000 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1107.1900 2161.2200 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1544.3800 1952.6000 1545.9800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1544.3800 2161.2200 1545.9800 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1956.5600 642.4800 1958.1600 1092.3000 ;
        RECT 2154.0600 642.4800 2155.6600 1092.3000 ;
        RECT 1964.3200 647.9100 1965.9200 1086.7000 ;
        RECT 2009.3200 647.9100 2010.9200 1086.7000 ;
        RECT 2054.3200 647.9100 2055.9200 1086.7000 ;
        RECT 2099.3200 647.9100 2100.9200 1086.7000 ;
        RECT 2144.3200 647.9100 2145.9200 1086.7000 ;
      LAYER met3 ;
        RECT 2154.0600 1081.8600 2155.6600 1082.3400 ;
        RECT 2154.0600 1076.4200 2155.6600 1076.9000 ;
        RECT 2154.0600 1070.9800 2155.6600 1071.4600 ;
        RECT 2154.0600 1065.5400 2155.6600 1066.0200 ;
        RECT 2154.0600 1060.1000 2155.6600 1060.5800 ;
        RECT 2154.0600 1054.6600 2155.6600 1055.1400 ;
        RECT 2154.0600 1049.2200 2155.6600 1049.7000 ;
        RECT 2154.0600 1043.7800 2155.6600 1044.2600 ;
        RECT 2154.0600 1038.3400 2155.6600 1038.8200 ;
        RECT 2154.0600 1032.9000 2155.6600 1033.3800 ;
        RECT 2154.0600 1027.4600 2155.6600 1027.9400 ;
        RECT 2154.0600 1022.0200 2155.6600 1022.5000 ;
        RECT 2154.0600 1016.5800 2155.6600 1017.0600 ;
        RECT 2154.0600 1011.1400 2155.6600 1011.6200 ;
        RECT 2154.0600 1005.7000 2155.6600 1006.1800 ;
        RECT 2154.0600 1000.2600 2155.6600 1000.7400 ;
        RECT 2154.0600 994.8200 2155.6600 995.3000 ;
        RECT 2154.0600 989.3800 2155.6600 989.8600 ;
        RECT 2154.0600 983.9400 2155.6600 984.4200 ;
        RECT 2154.0600 978.5000 2155.6600 978.9800 ;
        RECT 2154.0600 973.0600 2155.6600 973.5400 ;
        RECT 2154.0600 967.6200 2155.6600 968.1000 ;
        RECT 2154.0600 962.1800 2155.6600 962.6600 ;
        RECT 2154.0600 956.7400 2155.6600 957.2200 ;
        RECT 2154.0600 945.8600 2155.6600 946.3400 ;
        RECT 2154.0600 940.4200 2155.6600 940.9000 ;
        RECT 2154.0600 934.9800 2155.6600 935.4600 ;
        RECT 2154.0600 929.5400 2155.6600 930.0200 ;
        RECT 2154.0600 924.1000 2155.6600 924.5800 ;
        RECT 2154.0600 951.3000 2155.6600 951.7800 ;
        RECT 2154.0600 918.6600 2155.6600 919.1400 ;
        RECT 2154.0600 913.2200 2155.6600 913.7000 ;
        RECT 2154.0600 907.7800 2155.6600 908.2600 ;
        RECT 2154.0600 902.3400 2155.6600 902.8200 ;
        RECT 2154.0600 896.9000 2155.6600 897.3800 ;
        RECT 2154.0600 891.4600 2155.6600 891.9400 ;
        RECT 2154.0600 886.0200 2155.6600 886.5000 ;
        RECT 2154.0600 880.5800 2155.6600 881.0600 ;
        RECT 2154.0600 875.1400 2155.6600 875.6200 ;
        RECT 2154.0600 869.7000 2155.6600 870.1800 ;
        RECT 1956.5600 1081.8600 1958.1600 1082.3400 ;
        RECT 1956.5600 1076.4200 1958.1600 1076.9000 ;
        RECT 1956.5600 1070.9800 1958.1600 1071.4600 ;
        RECT 1956.5600 1065.5400 1958.1600 1066.0200 ;
        RECT 1956.5600 1060.1000 1958.1600 1060.5800 ;
        RECT 1956.5600 1054.6600 1958.1600 1055.1400 ;
        RECT 1956.5600 1049.2200 1958.1600 1049.7000 ;
        RECT 1956.5600 1043.7800 1958.1600 1044.2600 ;
        RECT 1956.5600 1038.3400 1958.1600 1038.8200 ;
        RECT 1956.5600 1032.9000 1958.1600 1033.3800 ;
        RECT 1956.5600 1027.4600 1958.1600 1027.9400 ;
        RECT 1956.5600 1022.0200 1958.1600 1022.5000 ;
        RECT 1956.5600 1016.5800 1958.1600 1017.0600 ;
        RECT 1956.5600 1011.1400 1958.1600 1011.6200 ;
        RECT 1956.5600 1005.7000 1958.1600 1006.1800 ;
        RECT 1956.5600 1000.2600 1958.1600 1000.7400 ;
        RECT 1956.5600 994.8200 1958.1600 995.3000 ;
        RECT 1956.5600 989.3800 1958.1600 989.8600 ;
        RECT 1956.5600 983.9400 1958.1600 984.4200 ;
        RECT 1956.5600 978.5000 1958.1600 978.9800 ;
        RECT 1956.5600 973.0600 1958.1600 973.5400 ;
        RECT 1956.5600 967.6200 1958.1600 968.1000 ;
        RECT 1956.5600 962.1800 1958.1600 962.6600 ;
        RECT 1956.5600 956.7400 1958.1600 957.2200 ;
        RECT 1956.5600 945.8600 1958.1600 946.3400 ;
        RECT 1956.5600 940.4200 1958.1600 940.9000 ;
        RECT 1956.5600 934.9800 1958.1600 935.4600 ;
        RECT 1956.5600 929.5400 1958.1600 930.0200 ;
        RECT 1956.5600 924.1000 1958.1600 924.5800 ;
        RECT 1956.5600 951.3000 1958.1600 951.7800 ;
        RECT 1956.5600 918.6600 1958.1600 919.1400 ;
        RECT 1956.5600 913.2200 1958.1600 913.7000 ;
        RECT 1956.5600 907.7800 1958.1600 908.2600 ;
        RECT 1956.5600 902.3400 1958.1600 902.8200 ;
        RECT 1956.5600 896.9000 1958.1600 897.3800 ;
        RECT 1956.5600 891.4600 1958.1600 891.9400 ;
        RECT 1956.5600 886.0200 1958.1600 886.5000 ;
        RECT 1956.5600 880.5800 1958.1600 881.0600 ;
        RECT 1956.5600 875.1400 1958.1600 875.6200 ;
        RECT 1956.5600 869.7000 1958.1600 870.1800 ;
        RECT 2154.0600 864.2600 2155.6600 864.7400 ;
        RECT 2154.0600 858.8200 2155.6600 859.3000 ;
        RECT 2154.0600 853.3800 2155.6600 853.8600 ;
        RECT 2154.0600 847.9400 2155.6600 848.4200 ;
        RECT 2154.0600 842.5000 2155.6600 842.9800 ;
        RECT 2154.0600 837.0600 2155.6600 837.5400 ;
        RECT 2154.0600 831.6200 2155.6600 832.1000 ;
        RECT 2154.0600 826.1800 2155.6600 826.6600 ;
        RECT 2154.0600 820.7400 2155.6600 821.2200 ;
        RECT 2154.0600 815.3000 2155.6600 815.7800 ;
        RECT 2154.0600 809.8600 2155.6600 810.3400 ;
        RECT 2154.0600 804.4200 2155.6600 804.9000 ;
        RECT 2154.0600 798.9800 2155.6600 799.4600 ;
        RECT 2154.0600 793.5400 2155.6600 794.0200 ;
        RECT 2154.0600 788.1000 2155.6600 788.5800 ;
        RECT 2154.0600 777.2200 2155.6600 777.7000 ;
        RECT 2154.0600 771.7800 2155.6600 772.2600 ;
        RECT 2154.0600 766.3400 2155.6600 766.8200 ;
        RECT 2154.0600 760.9000 2155.6600 761.3800 ;
        RECT 2154.0600 755.4600 2155.6600 755.9400 ;
        RECT 2154.0600 782.6600 2155.6600 783.1400 ;
        RECT 2154.0600 750.0200 2155.6600 750.5000 ;
        RECT 2154.0600 744.5800 2155.6600 745.0600 ;
        RECT 2154.0600 739.1400 2155.6600 739.6200 ;
        RECT 2154.0600 733.7000 2155.6600 734.1800 ;
        RECT 2154.0600 728.2600 2155.6600 728.7400 ;
        RECT 2154.0600 722.8200 2155.6600 723.3000 ;
        RECT 2154.0600 717.3800 2155.6600 717.8600 ;
        RECT 2154.0600 711.9400 2155.6600 712.4200 ;
        RECT 2154.0600 706.5000 2155.6600 706.9800 ;
        RECT 2154.0600 701.0600 2155.6600 701.5400 ;
        RECT 2154.0600 695.6200 2155.6600 696.1000 ;
        RECT 2154.0600 690.1800 2155.6600 690.6600 ;
        RECT 2154.0600 684.7400 2155.6600 685.2200 ;
        RECT 2154.0600 679.3000 2155.6600 679.7800 ;
        RECT 2154.0600 673.8600 2155.6600 674.3400 ;
        RECT 2154.0600 668.4200 2155.6600 668.9000 ;
        RECT 2154.0600 662.9800 2155.6600 663.4600 ;
        RECT 2154.0600 657.5400 2155.6600 658.0200 ;
        RECT 2154.0600 652.1000 2155.6600 652.5800 ;
        RECT 1956.5600 864.2600 1958.1600 864.7400 ;
        RECT 1956.5600 858.8200 1958.1600 859.3000 ;
        RECT 1956.5600 853.3800 1958.1600 853.8600 ;
        RECT 1956.5600 847.9400 1958.1600 848.4200 ;
        RECT 1956.5600 842.5000 1958.1600 842.9800 ;
        RECT 1956.5600 837.0600 1958.1600 837.5400 ;
        RECT 1956.5600 831.6200 1958.1600 832.1000 ;
        RECT 1956.5600 826.1800 1958.1600 826.6600 ;
        RECT 1956.5600 820.7400 1958.1600 821.2200 ;
        RECT 1956.5600 815.3000 1958.1600 815.7800 ;
        RECT 1956.5600 809.8600 1958.1600 810.3400 ;
        RECT 1956.5600 804.4200 1958.1600 804.9000 ;
        RECT 1956.5600 798.9800 1958.1600 799.4600 ;
        RECT 1956.5600 793.5400 1958.1600 794.0200 ;
        RECT 1956.5600 788.1000 1958.1600 788.5800 ;
        RECT 1956.5600 777.2200 1958.1600 777.7000 ;
        RECT 1956.5600 771.7800 1958.1600 772.2600 ;
        RECT 1956.5600 766.3400 1958.1600 766.8200 ;
        RECT 1956.5600 760.9000 1958.1600 761.3800 ;
        RECT 1956.5600 755.4600 1958.1600 755.9400 ;
        RECT 1956.5600 782.6600 1958.1600 783.1400 ;
        RECT 1956.5600 750.0200 1958.1600 750.5000 ;
        RECT 1956.5600 744.5800 1958.1600 745.0600 ;
        RECT 1956.5600 739.1400 1958.1600 739.6200 ;
        RECT 1956.5600 733.7000 1958.1600 734.1800 ;
        RECT 1956.5600 728.2600 1958.1600 728.7400 ;
        RECT 1956.5600 722.8200 1958.1600 723.3000 ;
        RECT 1956.5600 717.3800 1958.1600 717.8600 ;
        RECT 1956.5600 711.9400 1958.1600 712.4200 ;
        RECT 1956.5600 706.5000 1958.1600 706.9800 ;
        RECT 1956.5600 701.0600 1958.1600 701.5400 ;
        RECT 1956.5600 695.6200 1958.1600 696.1000 ;
        RECT 1956.5600 690.1800 1958.1600 690.6600 ;
        RECT 1956.5600 684.7400 1958.1600 685.2200 ;
        RECT 1956.5600 679.3000 1958.1600 679.7800 ;
        RECT 1956.5600 673.8600 1958.1600 674.3400 ;
        RECT 1956.5600 668.4200 1958.1600 668.9000 ;
        RECT 1956.5600 662.9800 1958.1600 663.4600 ;
        RECT 1956.5600 657.5400 1958.1600 658.0200 ;
        RECT 1956.5600 652.1000 1958.1600 652.5800 ;
        RECT 1951.0000 1085.1000 2161.2200 1086.7000 ;
        RECT 1951.0000 647.9100 2161.2200 649.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 642.4800 1958.1600 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 1090.7000 1958.1600 1092.3000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 642.4800 2155.6600 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 1090.7000 2155.6600 1092.3000 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 647.9100 1952.6000 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 647.9100 2161.2200 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 1085.1000 1952.6000 1086.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 1085.1000 2161.2200 1086.7000 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'DSP'
    PORT
      LAYER met4 ;
        RECT 1956.5600 183.2000 1958.1600 633.0200 ;
        RECT 2154.0600 183.2000 2155.6600 633.0200 ;
        RECT 1964.3200 188.6300 1965.9200 627.4200 ;
        RECT 2009.3200 188.6300 2010.9200 627.4200 ;
        RECT 2054.3200 188.6300 2055.9200 627.4200 ;
        RECT 2099.3200 188.6300 2100.9200 627.4200 ;
        RECT 2144.3200 188.6300 2145.9200 627.4200 ;
      LAYER met3 ;
        RECT 2154.0600 622.5800 2155.6600 623.0600 ;
        RECT 2154.0600 617.1400 2155.6600 617.6200 ;
        RECT 2154.0600 611.7000 2155.6600 612.1800 ;
        RECT 2154.0600 606.2600 2155.6600 606.7400 ;
        RECT 2154.0600 600.8200 2155.6600 601.3000 ;
        RECT 2154.0600 595.3800 2155.6600 595.8600 ;
        RECT 2154.0600 589.9400 2155.6600 590.4200 ;
        RECT 2154.0600 584.5000 2155.6600 584.9800 ;
        RECT 2154.0600 579.0600 2155.6600 579.5400 ;
        RECT 2154.0600 573.6200 2155.6600 574.1000 ;
        RECT 2154.0600 568.1800 2155.6600 568.6600 ;
        RECT 2154.0600 562.7400 2155.6600 563.2200 ;
        RECT 2154.0600 557.3000 2155.6600 557.7800 ;
        RECT 2154.0600 551.8600 2155.6600 552.3400 ;
        RECT 2154.0600 546.4200 2155.6600 546.9000 ;
        RECT 2154.0600 540.9800 2155.6600 541.4600 ;
        RECT 2154.0600 535.5400 2155.6600 536.0200 ;
        RECT 2154.0600 530.1000 2155.6600 530.5800 ;
        RECT 2154.0600 524.6600 2155.6600 525.1400 ;
        RECT 2154.0600 519.2200 2155.6600 519.7000 ;
        RECT 2154.0600 513.7800 2155.6600 514.2600 ;
        RECT 2154.0600 508.3400 2155.6600 508.8200 ;
        RECT 2154.0600 502.9000 2155.6600 503.3800 ;
        RECT 2154.0600 497.4600 2155.6600 497.9400 ;
        RECT 2154.0600 486.5800 2155.6600 487.0600 ;
        RECT 2154.0600 481.1400 2155.6600 481.6200 ;
        RECT 2154.0600 475.7000 2155.6600 476.1800 ;
        RECT 2154.0600 470.2600 2155.6600 470.7400 ;
        RECT 2154.0600 464.8200 2155.6600 465.3000 ;
        RECT 2154.0600 492.0200 2155.6600 492.5000 ;
        RECT 2154.0600 459.3800 2155.6600 459.8600 ;
        RECT 2154.0600 453.9400 2155.6600 454.4200 ;
        RECT 2154.0600 448.5000 2155.6600 448.9800 ;
        RECT 2154.0600 443.0600 2155.6600 443.5400 ;
        RECT 2154.0600 437.6200 2155.6600 438.1000 ;
        RECT 2154.0600 432.1800 2155.6600 432.6600 ;
        RECT 2154.0600 426.7400 2155.6600 427.2200 ;
        RECT 2154.0600 421.3000 2155.6600 421.7800 ;
        RECT 2154.0600 415.8600 2155.6600 416.3400 ;
        RECT 2154.0600 410.4200 2155.6600 410.9000 ;
        RECT 1956.5600 622.5800 1958.1600 623.0600 ;
        RECT 1956.5600 617.1400 1958.1600 617.6200 ;
        RECT 1956.5600 611.7000 1958.1600 612.1800 ;
        RECT 1956.5600 606.2600 1958.1600 606.7400 ;
        RECT 1956.5600 600.8200 1958.1600 601.3000 ;
        RECT 1956.5600 595.3800 1958.1600 595.8600 ;
        RECT 1956.5600 589.9400 1958.1600 590.4200 ;
        RECT 1956.5600 584.5000 1958.1600 584.9800 ;
        RECT 1956.5600 579.0600 1958.1600 579.5400 ;
        RECT 1956.5600 573.6200 1958.1600 574.1000 ;
        RECT 1956.5600 568.1800 1958.1600 568.6600 ;
        RECT 1956.5600 562.7400 1958.1600 563.2200 ;
        RECT 1956.5600 557.3000 1958.1600 557.7800 ;
        RECT 1956.5600 551.8600 1958.1600 552.3400 ;
        RECT 1956.5600 546.4200 1958.1600 546.9000 ;
        RECT 1956.5600 540.9800 1958.1600 541.4600 ;
        RECT 1956.5600 535.5400 1958.1600 536.0200 ;
        RECT 1956.5600 530.1000 1958.1600 530.5800 ;
        RECT 1956.5600 524.6600 1958.1600 525.1400 ;
        RECT 1956.5600 519.2200 1958.1600 519.7000 ;
        RECT 1956.5600 513.7800 1958.1600 514.2600 ;
        RECT 1956.5600 508.3400 1958.1600 508.8200 ;
        RECT 1956.5600 502.9000 1958.1600 503.3800 ;
        RECT 1956.5600 497.4600 1958.1600 497.9400 ;
        RECT 1956.5600 486.5800 1958.1600 487.0600 ;
        RECT 1956.5600 481.1400 1958.1600 481.6200 ;
        RECT 1956.5600 475.7000 1958.1600 476.1800 ;
        RECT 1956.5600 470.2600 1958.1600 470.7400 ;
        RECT 1956.5600 464.8200 1958.1600 465.3000 ;
        RECT 1956.5600 492.0200 1958.1600 492.5000 ;
        RECT 1956.5600 459.3800 1958.1600 459.8600 ;
        RECT 1956.5600 453.9400 1958.1600 454.4200 ;
        RECT 1956.5600 448.5000 1958.1600 448.9800 ;
        RECT 1956.5600 443.0600 1958.1600 443.5400 ;
        RECT 1956.5600 437.6200 1958.1600 438.1000 ;
        RECT 1956.5600 432.1800 1958.1600 432.6600 ;
        RECT 1956.5600 426.7400 1958.1600 427.2200 ;
        RECT 1956.5600 421.3000 1958.1600 421.7800 ;
        RECT 1956.5600 415.8600 1958.1600 416.3400 ;
        RECT 1956.5600 410.4200 1958.1600 410.9000 ;
        RECT 2154.0600 404.9800 2155.6600 405.4600 ;
        RECT 2154.0600 399.5400 2155.6600 400.0200 ;
        RECT 2154.0600 394.1000 2155.6600 394.5800 ;
        RECT 2154.0600 388.6600 2155.6600 389.1400 ;
        RECT 2154.0600 383.2200 2155.6600 383.7000 ;
        RECT 2154.0600 377.7800 2155.6600 378.2600 ;
        RECT 2154.0600 372.3400 2155.6600 372.8200 ;
        RECT 2154.0600 366.9000 2155.6600 367.3800 ;
        RECT 2154.0600 361.4600 2155.6600 361.9400 ;
        RECT 2154.0600 356.0200 2155.6600 356.5000 ;
        RECT 2154.0600 350.5800 2155.6600 351.0600 ;
        RECT 2154.0600 345.1400 2155.6600 345.6200 ;
        RECT 2154.0600 339.7000 2155.6600 340.1800 ;
        RECT 2154.0600 334.2600 2155.6600 334.7400 ;
        RECT 2154.0600 328.8200 2155.6600 329.3000 ;
        RECT 2154.0600 317.9400 2155.6600 318.4200 ;
        RECT 2154.0600 312.5000 2155.6600 312.9800 ;
        RECT 2154.0600 307.0600 2155.6600 307.5400 ;
        RECT 2154.0600 301.6200 2155.6600 302.1000 ;
        RECT 2154.0600 296.1800 2155.6600 296.6600 ;
        RECT 2154.0600 323.3800 2155.6600 323.8600 ;
        RECT 2154.0600 290.7400 2155.6600 291.2200 ;
        RECT 2154.0600 285.3000 2155.6600 285.7800 ;
        RECT 2154.0600 279.8600 2155.6600 280.3400 ;
        RECT 2154.0600 274.4200 2155.6600 274.9000 ;
        RECT 2154.0600 268.9800 2155.6600 269.4600 ;
        RECT 2154.0600 263.5400 2155.6600 264.0200 ;
        RECT 2154.0600 258.1000 2155.6600 258.5800 ;
        RECT 2154.0600 252.6600 2155.6600 253.1400 ;
        RECT 2154.0600 247.2200 2155.6600 247.7000 ;
        RECT 2154.0600 241.7800 2155.6600 242.2600 ;
        RECT 2154.0600 236.3400 2155.6600 236.8200 ;
        RECT 2154.0600 230.9000 2155.6600 231.3800 ;
        RECT 2154.0600 225.4600 2155.6600 225.9400 ;
        RECT 2154.0600 220.0200 2155.6600 220.5000 ;
        RECT 2154.0600 214.5800 2155.6600 215.0600 ;
        RECT 2154.0600 209.1400 2155.6600 209.6200 ;
        RECT 2154.0600 203.7000 2155.6600 204.1800 ;
        RECT 2154.0600 198.2600 2155.6600 198.7400 ;
        RECT 2154.0600 192.8200 2155.6600 193.3000 ;
        RECT 1956.5600 404.9800 1958.1600 405.4600 ;
        RECT 1956.5600 399.5400 1958.1600 400.0200 ;
        RECT 1956.5600 394.1000 1958.1600 394.5800 ;
        RECT 1956.5600 388.6600 1958.1600 389.1400 ;
        RECT 1956.5600 383.2200 1958.1600 383.7000 ;
        RECT 1956.5600 377.7800 1958.1600 378.2600 ;
        RECT 1956.5600 372.3400 1958.1600 372.8200 ;
        RECT 1956.5600 366.9000 1958.1600 367.3800 ;
        RECT 1956.5600 361.4600 1958.1600 361.9400 ;
        RECT 1956.5600 356.0200 1958.1600 356.5000 ;
        RECT 1956.5600 350.5800 1958.1600 351.0600 ;
        RECT 1956.5600 345.1400 1958.1600 345.6200 ;
        RECT 1956.5600 339.7000 1958.1600 340.1800 ;
        RECT 1956.5600 334.2600 1958.1600 334.7400 ;
        RECT 1956.5600 328.8200 1958.1600 329.3000 ;
        RECT 1956.5600 317.9400 1958.1600 318.4200 ;
        RECT 1956.5600 312.5000 1958.1600 312.9800 ;
        RECT 1956.5600 307.0600 1958.1600 307.5400 ;
        RECT 1956.5600 301.6200 1958.1600 302.1000 ;
        RECT 1956.5600 296.1800 1958.1600 296.6600 ;
        RECT 1956.5600 323.3800 1958.1600 323.8600 ;
        RECT 1956.5600 290.7400 1958.1600 291.2200 ;
        RECT 1956.5600 285.3000 1958.1600 285.7800 ;
        RECT 1956.5600 279.8600 1958.1600 280.3400 ;
        RECT 1956.5600 274.4200 1958.1600 274.9000 ;
        RECT 1956.5600 268.9800 1958.1600 269.4600 ;
        RECT 1956.5600 263.5400 1958.1600 264.0200 ;
        RECT 1956.5600 258.1000 1958.1600 258.5800 ;
        RECT 1956.5600 252.6600 1958.1600 253.1400 ;
        RECT 1956.5600 247.2200 1958.1600 247.7000 ;
        RECT 1956.5600 241.7800 1958.1600 242.2600 ;
        RECT 1956.5600 236.3400 1958.1600 236.8200 ;
        RECT 1956.5600 230.9000 1958.1600 231.3800 ;
        RECT 1956.5600 225.4600 1958.1600 225.9400 ;
        RECT 1956.5600 220.0200 1958.1600 220.5000 ;
        RECT 1956.5600 214.5800 1958.1600 215.0600 ;
        RECT 1956.5600 209.1400 1958.1600 209.6200 ;
        RECT 1956.5600 203.7000 1958.1600 204.1800 ;
        RECT 1956.5600 198.2600 1958.1600 198.7400 ;
        RECT 1956.5600 192.8200 1958.1600 193.3000 ;
        RECT 1951.0000 625.8200 2161.2200 627.4200 ;
        RECT 1951.0000 188.6300 2161.2200 190.2300 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 183.2000 1958.1600 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.5600 631.4200 1958.1600 633.0200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 183.2000 2155.6600 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2154.0600 631.4200 2155.6600 633.0200 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 188.6300 1952.6000 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 188.6300 2161.2200 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 1951.0000 625.8200 1952.6000 627.4200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2159.6200 625.8200 2161.2200 627.4200 ;
    END
# end of P/G pin shape extracted from block 'DSP'


# P/G pin shape extracted from block 'N_term_single'
    PORT
      LAYER met4 ;
        RECT 2176.6800 2479.6000 2178.2800 2509.8600 ;
        RECT 2374.3800 2479.6000 2375.9800 2509.8600 ;
      LAYER met3 ;
        RECT 2374.3800 2497.3800 2375.9800 2497.8600 ;
        RECT 2176.6800 2497.3800 2178.2800 2497.8600 ;
        RECT 2374.3800 2491.9400 2375.9800 2492.4200 ;
        RECT 2374.3800 2486.5000 2375.9800 2486.9800 ;
        RECT 2176.6800 2491.9400 2178.2800 2492.4200 ;
        RECT 2176.6800 2486.5000 2178.2800 2486.9800 ;
        RECT 2171.2200 2503.1000 2381.4400 2504.7000 ;
        RECT 2171.2200 2483.5700 2381.4400 2485.1700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.6800 2479.6000 2178.2800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.6800 2508.2600 2178.2800 2509.8600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.3800 2479.6000 2375.9800 2481.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.3800 2508.2600 2375.9800 2509.8600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2483.5700 2172.8200 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2483.5700 2381.4400 2485.1700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2503.1000 2172.8200 2504.7000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2503.1000 2381.4400 2504.7000 ;
    END
# end of P/G pin shape extracted from block 'N_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 188.6300 2366.1400 396.7300 ;
        RECT 2319.5400 188.6300 2321.1400 396.7300 ;
        RECT 2274.5400 188.6300 2276.1400 396.7300 ;
        RECT 2229.5400 188.6300 2231.1400 396.7300 ;
        RECT 2184.5400 188.6300 2186.1400 396.7300 ;
        RECT 2374.2800 183.2000 2375.8800 402.8400 ;
        RECT 2176.7800 183.2000 2178.3800 402.8400 ;
      LAYER met3 ;
        RECT 2374.2800 377.7800 2375.8800 378.2600 ;
        RECT 2374.2800 383.2200 2375.8800 383.7000 ;
        RECT 2364.5400 377.7800 2366.1400 378.2600 ;
        RECT 2364.5400 383.2200 2366.1400 383.7000 ;
        RECT 2364.5400 388.6600 2366.1400 389.1400 ;
        RECT 2374.2800 388.6600 2375.8800 389.1400 ;
        RECT 2374.2800 366.9000 2375.8800 367.3800 ;
        RECT 2374.2800 372.3400 2375.8800 372.8200 ;
        RECT 2364.5400 366.9000 2366.1400 367.3800 ;
        RECT 2364.5400 372.3400 2366.1400 372.8200 ;
        RECT 2374.2800 350.5800 2375.8800 351.0600 ;
        RECT 2374.2800 356.0200 2375.8800 356.5000 ;
        RECT 2364.5400 350.5800 2366.1400 351.0600 ;
        RECT 2364.5400 356.0200 2366.1400 356.5000 ;
        RECT 2364.5400 361.4600 2366.1400 361.9400 ;
        RECT 2374.2800 361.4600 2375.8800 361.9400 ;
        RECT 2319.5400 377.7800 2321.1400 378.2600 ;
        RECT 2319.5400 383.2200 2321.1400 383.7000 ;
        RECT 2319.5400 388.6600 2321.1400 389.1400 ;
        RECT 2319.5400 366.9000 2321.1400 367.3800 ;
        RECT 2319.5400 372.3400 2321.1400 372.8200 ;
        RECT 2319.5400 350.5800 2321.1400 351.0600 ;
        RECT 2319.5400 356.0200 2321.1400 356.5000 ;
        RECT 2319.5400 361.4600 2321.1400 361.9400 ;
        RECT 2374.2800 334.2600 2375.8800 334.7400 ;
        RECT 2374.2800 339.7000 2375.8800 340.1800 ;
        RECT 2374.2800 345.1400 2375.8800 345.6200 ;
        RECT 2364.5400 334.2600 2366.1400 334.7400 ;
        RECT 2364.5400 339.7000 2366.1400 340.1800 ;
        RECT 2364.5400 345.1400 2366.1400 345.6200 ;
        RECT 2374.2800 323.3800 2375.8800 323.8600 ;
        RECT 2374.2800 328.8200 2375.8800 329.3000 ;
        RECT 2364.5400 323.3800 2366.1400 323.8600 ;
        RECT 2364.5400 328.8200 2366.1400 329.3000 ;
        RECT 2374.2800 307.0600 2375.8800 307.5400 ;
        RECT 2374.2800 312.5000 2375.8800 312.9800 ;
        RECT 2374.2800 317.9400 2375.8800 318.4200 ;
        RECT 2364.5400 307.0600 2366.1400 307.5400 ;
        RECT 2364.5400 312.5000 2366.1400 312.9800 ;
        RECT 2364.5400 317.9400 2366.1400 318.4200 ;
        RECT 2374.2800 296.1800 2375.8800 296.6600 ;
        RECT 2374.2800 301.6200 2375.8800 302.1000 ;
        RECT 2364.5400 296.1800 2366.1400 296.6600 ;
        RECT 2364.5400 301.6200 2366.1400 302.1000 ;
        RECT 2319.5400 334.2600 2321.1400 334.7400 ;
        RECT 2319.5400 339.7000 2321.1400 340.1800 ;
        RECT 2319.5400 345.1400 2321.1400 345.6200 ;
        RECT 2319.5400 323.3800 2321.1400 323.8600 ;
        RECT 2319.5400 328.8200 2321.1400 329.3000 ;
        RECT 2319.5400 307.0600 2321.1400 307.5400 ;
        RECT 2319.5400 312.5000 2321.1400 312.9800 ;
        RECT 2319.5400 317.9400 2321.1400 318.4200 ;
        RECT 2319.5400 296.1800 2321.1400 296.6600 ;
        RECT 2319.5400 301.6200 2321.1400 302.1000 ;
        RECT 2274.5400 377.7800 2276.1400 378.2600 ;
        RECT 2274.5400 383.2200 2276.1400 383.7000 ;
        RECT 2274.5400 388.6600 2276.1400 389.1400 ;
        RECT 2229.5400 377.7800 2231.1400 378.2600 ;
        RECT 2229.5400 383.2200 2231.1400 383.7000 ;
        RECT 2229.5400 388.6600 2231.1400 389.1400 ;
        RECT 2274.5400 366.9000 2276.1400 367.3800 ;
        RECT 2274.5400 372.3400 2276.1400 372.8200 ;
        RECT 2274.5400 350.5800 2276.1400 351.0600 ;
        RECT 2274.5400 356.0200 2276.1400 356.5000 ;
        RECT 2274.5400 361.4600 2276.1400 361.9400 ;
        RECT 2229.5400 366.9000 2231.1400 367.3800 ;
        RECT 2229.5400 372.3400 2231.1400 372.8200 ;
        RECT 2229.5400 350.5800 2231.1400 351.0600 ;
        RECT 2229.5400 356.0200 2231.1400 356.5000 ;
        RECT 2229.5400 361.4600 2231.1400 361.9400 ;
        RECT 2184.5400 377.7800 2186.1400 378.2600 ;
        RECT 2184.5400 383.2200 2186.1400 383.7000 ;
        RECT 2176.7800 377.7800 2178.3800 378.2600 ;
        RECT 2176.7800 383.2200 2178.3800 383.7000 ;
        RECT 2176.7800 388.6600 2178.3800 389.1400 ;
        RECT 2184.5400 388.6600 2186.1400 389.1400 ;
        RECT 2184.5400 366.9000 2186.1400 367.3800 ;
        RECT 2184.5400 372.3400 2186.1400 372.8200 ;
        RECT 2176.7800 366.9000 2178.3800 367.3800 ;
        RECT 2176.7800 372.3400 2178.3800 372.8200 ;
        RECT 2184.5400 350.5800 2186.1400 351.0600 ;
        RECT 2184.5400 356.0200 2186.1400 356.5000 ;
        RECT 2176.7800 350.5800 2178.3800 351.0600 ;
        RECT 2176.7800 356.0200 2178.3800 356.5000 ;
        RECT 2176.7800 361.4600 2178.3800 361.9400 ;
        RECT 2184.5400 361.4600 2186.1400 361.9400 ;
        RECT 2274.5400 334.2600 2276.1400 334.7400 ;
        RECT 2274.5400 339.7000 2276.1400 340.1800 ;
        RECT 2274.5400 345.1400 2276.1400 345.6200 ;
        RECT 2274.5400 323.3800 2276.1400 323.8600 ;
        RECT 2274.5400 328.8200 2276.1400 329.3000 ;
        RECT 2229.5400 334.2600 2231.1400 334.7400 ;
        RECT 2229.5400 339.7000 2231.1400 340.1800 ;
        RECT 2229.5400 345.1400 2231.1400 345.6200 ;
        RECT 2229.5400 323.3800 2231.1400 323.8600 ;
        RECT 2229.5400 328.8200 2231.1400 329.3000 ;
        RECT 2274.5400 307.0600 2276.1400 307.5400 ;
        RECT 2274.5400 312.5000 2276.1400 312.9800 ;
        RECT 2274.5400 317.9400 2276.1400 318.4200 ;
        RECT 2274.5400 296.1800 2276.1400 296.6600 ;
        RECT 2274.5400 301.6200 2276.1400 302.1000 ;
        RECT 2229.5400 307.0600 2231.1400 307.5400 ;
        RECT 2229.5400 312.5000 2231.1400 312.9800 ;
        RECT 2229.5400 317.9400 2231.1400 318.4200 ;
        RECT 2229.5400 296.1800 2231.1400 296.6600 ;
        RECT 2229.5400 301.6200 2231.1400 302.1000 ;
        RECT 2184.5400 334.2600 2186.1400 334.7400 ;
        RECT 2184.5400 339.7000 2186.1400 340.1800 ;
        RECT 2184.5400 345.1400 2186.1400 345.6200 ;
        RECT 2176.7800 334.2600 2178.3800 334.7400 ;
        RECT 2176.7800 339.7000 2178.3800 340.1800 ;
        RECT 2176.7800 345.1400 2178.3800 345.6200 ;
        RECT 2184.5400 323.3800 2186.1400 323.8600 ;
        RECT 2184.5400 328.8200 2186.1400 329.3000 ;
        RECT 2176.7800 323.3800 2178.3800 323.8600 ;
        RECT 2176.7800 328.8200 2178.3800 329.3000 ;
        RECT 2184.5400 307.0600 2186.1400 307.5400 ;
        RECT 2184.5400 312.5000 2186.1400 312.9800 ;
        RECT 2184.5400 317.9400 2186.1400 318.4200 ;
        RECT 2176.7800 307.0600 2178.3800 307.5400 ;
        RECT 2176.7800 312.5000 2178.3800 312.9800 ;
        RECT 2176.7800 317.9400 2178.3800 318.4200 ;
        RECT 2184.5400 296.1800 2186.1400 296.6600 ;
        RECT 2184.5400 301.6200 2186.1400 302.1000 ;
        RECT 2176.7800 296.1800 2178.3800 296.6600 ;
        RECT 2176.7800 301.6200 2178.3800 302.1000 ;
        RECT 2374.2800 279.8600 2375.8800 280.3400 ;
        RECT 2374.2800 285.3000 2375.8800 285.7800 ;
        RECT 2374.2800 290.7400 2375.8800 291.2200 ;
        RECT 2364.5400 279.8600 2366.1400 280.3400 ;
        RECT 2364.5400 285.3000 2366.1400 285.7800 ;
        RECT 2364.5400 290.7400 2366.1400 291.2200 ;
        RECT 2374.2800 268.9800 2375.8800 269.4600 ;
        RECT 2374.2800 274.4200 2375.8800 274.9000 ;
        RECT 2364.5400 268.9800 2366.1400 269.4600 ;
        RECT 2364.5400 274.4200 2366.1400 274.9000 ;
        RECT 2374.2800 252.6600 2375.8800 253.1400 ;
        RECT 2374.2800 258.1000 2375.8800 258.5800 ;
        RECT 2374.2800 263.5400 2375.8800 264.0200 ;
        RECT 2364.5400 252.6600 2366.1400 253.1400 ;
        RECT 2364.5400 258.1000 2366.1400 258.5800 ;
        RECT 2364.5400 263.5400 2366.1400 264.0200 ;
        RECT 2374.2800 241.7800 2375.8800 242.2600 ;
        RECT 2374.2800 247.2200 2375.8800 247.7000 ;
        RECT 2364.5400 241.7800 2366.1400 242.2600 ;
        RECT 2364.5400 247.2200 2366.1400 247.7000 ;
        RECT 2319.5400 279.8600 2321.1400 280.3400 ;
        RECT 2319.5400 285.3000 2321.1400 285.7800 ;
        RECT 2319.5400 290.7400 2321.1400 291.2200 ;
        RECT 2319.5400 268.9800 2321.1400 269.4600 ;
        RECT 2319.5400 274.4200 2321.1400 274.9000 ;
        RECT 2319.5400 252.6600 2321.1400 253.1400 ;
        RECT 2319.5400 258.1000 2321.1400 258.5800 ;
        RECT 2319.5400 263.5400 2321.1400 264.0200 ;
        RECT 2319.5400 241.7800 2321.1400 242.2600 ;
        RECT 2319.5400 247.2200 2321.1400 247.7000 ;
        RECT 2374.2800 225.4600 2375.8800 225.9400 ;
        RECT 2374.2800 230.9000 2375.8800 231.3800 ;
        RECT 2374.2800 236.3400 2375.8800 236.8200 ;
        RECT 2364.5400 225.4600 2366.1400 225.9400 ;
        RECT 2364.5400 230.9000 2366.1400 231.3800 ;
        RECT 2364.5400 236.3400 2366.1400 236.8200 ;
        RECT 2374.2800 214.5800 2375.8800 215.0600 ;
        RECT 2374.2800 220.0200 2375.8800 220.5000 ;
        RECT 2364.5400 214.5800 2366.1400 215.0600 ;
        RECT 2364.5400 220.0200 2366.1400 220.5000 ;
        RECT 2374.2800 198.2600 2375.8800 198.7400 ;
        RECT 2374.2800 203.7000 2375.8800 204.1800 ;
        RECT 2374.2800 209.1400 2375.8800 209.6200 ;
        RECT 2364.5400 198.2600 2366.1400 198.7400 ;
        RECT 2364.5400 203.7000 2366.1400 204.1800 ;
        RECT 2364.5400 209.1400 2366.1400 209.6200 ;
        RECT 2364.5400 192.8200 2366.1400 193.3000 ;
        RECT 2374.2800 192.8200 2375.8800 193.3000 ;
        RECT 2319.5400 225.4600 2321.1400 225.9400 ;
        RECT 2319.5400 230.9000 2321.1400 231.3800 ;
        RECT 2319.5400 236.3400 2321.1400 236.8200 ;
        RECT 2319.5400 214.5800 2321.1400 215.0600 ;
        RECT 2319.5400 220.0200 2321.1400 220.5000 ;
        RECT 2319.5400 198.2600 2321.1400 198.7400 ;
        RECT 2319.5400 203.7000 2321.1400 204.1800 ;
        RECT 2319.5400 209.1400 2321.1400 209.6200 ;
        RECT 2319.5400 192.8200 2321.1400 193.3000 ;
        RECT 2274.5400 279.8600 2276.1400 280.3400 ;
        RECT 2274.5400 285.3000 2276.1400 285.7800 ;
        RECT 2274.5400 290.7400 2276.1400 291.2200 ;
        RECT 2274.5400 268.9800 2276.1400 269.4600 ;
        RECT 2274.5400 274.4200 2276.1400 274.9000 ;
        RECT 2229.5400 279.8600 2231.1400 280.3400 ;
        RECT 2229.5400 285.3000 2231.1400 285.7800 ;
        RECT 2229.5400 290.7400 2231.1400 291.2200 ;
        RECT 2229.5400 268.9800 2231.1400 269.4600 ;
        RECT 2229.5400 274.4200 2231.1400 274.9000 ;
        RECT 2274.5400 252.6600 2276.1400 253.1400 ;
        RECT 2274.5400 258.1000 2276.1400 258.5800 ;
        RECT 2274.5400 263.5400 2276.1400 264.0200 ;
        RECT 2274.5400 241.7800 2276.1400 242.2600 ;
        RECT 2274.5400 247.2200 2276.1400 247.7000 ;
        RECT 2229.5400 252.6600 2231.1400 253.1400 ;
        RECT 2229.5400 258.1000 2231.1400 258.5800 ;
        RECT 2229.5400 263.5400 2231.1400 264.0200 ;
        RECT 2229.5400 241.7800 2231.1400 242.2600 ;
        RECT 2229.5400 247.2200 2231.1400 247.7000 ;
        RECT 2184.5400 279.8600 2186.1400 280.3400 ;
        RECT 2184.5400 285.3000 2186.1400 285.7800 ;
        RECT 2184.5400 290.7400 2186.1400 291.2200 ;
        RECT 2176.7800 279.8600 2178.3800 280.3400 ;
        RECT 2176.7800 285.3000 2178.3800 285.7800 ;
        RECT 2176.7800 290.7400 2178.3800 291.2200 ;
        RECT 2184.5400 268.9800 2186.1400 269.4600 ;
        RECT 2184.5400 274.4200 2186.1400 274.9000 ;
        RECT 2176.7800 268.9800 2178.3800 269.4600 ;
        RECT 2176.7800 274.4200 2178.3800 274.9000 ;
        RECT 2184.5400 252.6600 2186.1400 253.1400 ;
        RECT 2184.5400 258.1000 2186.1400 258.5800 ;
        RECT 2184.5400 263.5400 2186.1400 264.0200 ;
        RECT 2176.7800 252.6600 2178.3800 253.1400 ;
        RECT 2176.7800 258.1000 2178.3800 258.5800 ;
        RECT 2176.7800 263.5400 2178.3800 264.0200 ;
        RECT 2184.5400 241.7800 2186.1400 242.2600 ;
        RECT 2184.5400 247.2200 2186.1400 247.7000 ;
        RECT 2176.7800 241.7800 2178.3800 242.2600 ;
        RECT 2176.7800 247.2200 2178.3800 247.7000 ;
        RECT 2274.5400 225.4600 2276.1400 225.9400 ;
        RECT 2274.5400 230.9000 2276.1400 231.3800 ;
        RECT 2274.5400 236.3400 2276.1400 236.8200 ;
        RECT 2274.5400 214.5800 2276.1400 215.0600 ;
        RECT 2274.5400 220.0200 2276.1400 220.5000 ;
        RECT 2229.5400 225.4600 2231.1400 225.9400 ;
        RECT 2229.5400 230.9000 2231.1400 231.3800 ;
        RECT 2229.5400 236.3400 2231.1400 236.8200 ;
        RECT 2229.5400 214.5800 2231.1400 215.0600 ;
        RECT 2229.5400 220.0200 2231.1400 220.5000 ;
        RECT 2274.5400 198.2600 2276.1400 198.7400 ;
        RECT 2274.5400 203.7000 2276.1400 204.1800 ;
        RECT 2274.5400 209.1400 2276.1400 209.6200 ;
        RECT 2274.5400 192.8200 2276.1400 193.3000 ;
        RECT 2229.5400 198.2600 2231.1400 198.7400 ;
        RECT 2229.5400 203.7000 2231.1400 204.1800 ;
        RECT 2229.5400 209.1400 2231.1400 209.6200 ;
        RECT 2229.5400 192.8200 2231.1400 193.3000 ;
        RECT 2184.5400 225.4600 2186.1400 225.9400 ;
        RECT 2184.5400 230.9000 2186.1400 231.3800 ;
        RECT 2184.5400 236.3400 2186.1400 236.8200 ;
        RECT 2176.7800 225.4600 2178.3800 225.9400 ;
        RECT 2176.7800 230.9000 2178.3800 231.3800 ;
        RECT 2176.7800 236.3400 2178.3800 236.8200 ;
        RECT 2184.5400 214.5800 2186.1400 215.0600 ;
        RECT 2184.5400 220.0200 2186.1400 220.5000 ;
        RECT 2176.7800 214.5800 2178.3800 215.0600 ;
        RECT 2176.7800 220.0200 2178.3800 220.5000 ;
        RECT 2184.5400 198.2600 2186.1400 198.7400 ;
        RECT 2184.5400 203.7000 2186.1400 204.1800 ;
        RECT 2184.5400 209.1400 2186.1400 209.6200 ;
        RECT 2176.7800 198.2600 2178.3800 198.7400 ;
        RECT 2176.7800 203.7000 2178.3800 204.1800 ;
        RECT 2176.7800 209.1400 2178.3800 209.6200 ;
        RECT 2176.7800 192.8200 2178.3800 193.3000 ;
        RECT 2184.5400 192.8200 2186.1400 193.3000 ;
        RECT 2171.2200 395.1300 2381.4400 396.7300 ;
        RECT 2171.2200 188.6300 2381.4400 190.2300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 183.2000 2178.3800 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 401.2400 2178.3800 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 183.2000 2375.8800 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 401.2400 2375.8800 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 188.6300 2172.8200 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 188.6300 2381.4400 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 395.1300 2172.8200 396.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 395.1300 2381.4400 396.7300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'S_term_single'
    PORT
      LAYER met4 ;
        RECT 2176.6800 142.9400 2178.2800 173.2000 ;
        RECT 2374.3800 142.9400 2375.9800 173.2000 ;
      LAYER met3 ;
        RECT 2374.3800 160.7200 2375.9800 161.2000 ;
        RECT 2176.6800 160.7200 2178.2800 161.2000 ;
        RECT 2374.3800 155.2800 2375.9800 155.7600 ;
        RECT 2374.3800 149.8400 2375.9800 150.3200 ;
        RECT 2176.6800 155.2800 2178.2800 155.7600 ;
        RECT 2176.6800 149.8400 2178.2800 150.3200 ;
        RECT 2171.2200 166.4400 2381.4400 168.0400 ;
        RECT 2171.2200 146.9100 2381.4400 148.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.6800 142.9400 2178.2800 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.6800 171.6000 2178.2800 173.2000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.3800 142.9400 2375.9800 144.5400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.3800 171.6000 2375.9800 173.2000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 146.9100 2172.8200 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 146.9100 2381.4400 148.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 166.4400 2172.8200 168.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 166.4400 2381.4400 168.0400 ;
    END
# end of P/G pin shape extracted from block 'S_term_single'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 2255.3900 2366.1400 2463.4900 ;
        RECT 2319.5400 2255.3900 2321.1400 2463.4900 ;
        RECT 2274.5400 2255.3900 2276.1400 2463.4900 ;
        RECT 2229.5400 2255.3900 2231.1400 2463.4900 ;
        RECT 2184.5400 2255.3900 2186.1400 2463.4900 ;
        RECT 2374.2800 2249.9600 2375.8800 2469.6000 ;
        RECT 2176.7800 2249.9600 2178.3800 2469.6000 ;
      LAYER met3 ;
        RECT 2374.2800 2444.5400 2375.8800 2445.0200 ;
        RECT 2374.2800 2449.9800 2375.8800 2450.4600 ;
        RECT 2364.5400 2444.5400 2366.1400 2445.0200 ;
        RECT 2364.5400 2449.9800 2366.1400 2450.4600 ;
        RECT 2364.5400 2455.4200 2366.1400 2455.9000 ;
        RECT 2374.2800 2455.4200 2375.8800 2455.9000 ;
        RECT 2374.2800 2433.6600 2375.8800 2434.1400 ;
        RECT 2374.2800 2439.1000 2375.8800 2439.5800 ;
        RECT 2364.5400 2433.6600 2366.1400 2434.1400 ;
        RECT 2364.5400 2439.1000 2366.1400 2439.5800 ;
        RECT 2374.2800 2417.3400 2375.8800 2417.8200 ;
        RECT 2374.2800 2422.7800 2375.8800 2423.2600 ;
        RECT 2364.5400 2417.3400 2366.1400 2417.8200 ;
        RECT 2364.5400 2422.7800 2366.1400 2423.2600 ;
        RECT 2364.5400 2428.2200 2366.1400 2428.7000 ;
        RECT 2374.2800 2428.2200 2375.8800 2428.7000 ;
        RECT 2319.5400 2444.5400 2321.1400 2445.0200 ;
        RECT 2319.5400 2449.9800 2321.1400 2450.4600 ;
        RECT 2319.5400 2455.4200 2321.1400 2455.9000 ;
        RECT 2319.5400 2433.6600 2321.1400 2434.1400 ;
        RECT 2319.5400 2439.1000 2321.1400 2439.5800 ;
        RECT 2319.5400 2417.3400 2321.1400 2417.8200 ;
        RECT 2319.5400 2422.7800 2321.1400 2423.2600 ;
        RECT 2319.5400 2428.2200 2321.1400 2428.7000 ;
        RECT 2374.2800 2401.0200 2375.8800 2401.5000 ;
        RECT 2374.2800 2406.4600 2375.8800 2406.9400 ;
        RECT 2374.2800 2411.9000 2375.8800 2412.3800 ;
        RECT 2364.5400 2401.0200 2366.1400 2401.5000 ;
        RECT 2364.5400 2406.4600 2366.1400 2406.9400 ;
        RECT 2364.5400 2411.9000 2366.1400 2412.3800 ;
        RECT 2374.2800 2390.1400 2375.8800 2390.6200 ;
        RECT 2374.2800 2395.5800 2375.8800 2396.0600 ;
        RECT 2364.5400 2390.1400 2366.1400 2390.6200 ;
        RECT 2364.5400 2395.5800 2366.1400 2396.0600 ;
        RECT 2374.2800 2373.8200 2375.8800 2374.3000 ;
        RECT 2374.2800 2379.2600 2375.8800 2379.7400 ;
        RECT 2374.2800 2384.7000 2375.8800 2385.1800 ;
        RECT 2364.5400 2373.8200 2366.1400 2374.3000 ;
        RECT 2364.5400 2379.2600 2366.1400 2379.7400 ;
        RECT 2364.5400 2384.7000 2366.1400 2385.1800 ;
        RECT 2374.2800 2362.9400 2375.8800 2363.4200 ;
        RECT 2374.2800 2368.3800 2375.8800 2368.8600 ;
        RECT 2364.5400 2362.9400 2366.1400 2363.4200 ;
        RECT 2364.5400 2368.3800 2366.1400 2368.8600 ;
        RECT 2319.5400 2401.0200 2321.1400 2401.5000 ;
        RECT 2319.5400 2406.4600 2321.1400 2406.9400 ;
        RECT 2319.5400 2411.9000 2321.1400 2412.3800 ;
        RECT 2319.5400 2390.1400 2321.1400 2390.6200 ;
        RECT 2319.5400 2395.5800 2321.1400 2396.0600 ;
        RECT 2319.5400 2373.8200 2321.1400 2374.3000 ;
        RECT 2319.5400 2379.2600 2321.1400 2379.7400 ;
        RECT 2319.5400 2384.7000 2321.1400 2385.1800 ;
        RECT 2319.5400 2362.9400 2321.1400 2363.4200 ;
        RECT 2319.5400 2368.3800 2321.1400 2368.8600 ;
        RECT 2274.5400 2444.5400 2276.1400 2445.0200 ;
        RECT 2274.5400 2449.9800 2276.1400 2450.4600 ;
        RECT 2274.5400 2455.4200 2276.1400 2455.9000 ;
        RECT 2229.5400 2444.5400 2231.1400 2445.0200 ;
        RECT 2229.5400 2449.9800 2231.1400 2450.4600 ;
        RECT 2229.5400 2455.4200 2231.1400 2455.9000 ;
        RECT 2274.5400 2433.6600 2276.1400 2434.1400 ;
        RECT 2274.5400 2439.1000 2276.1400 2439.5800 ;
        RECT 2274.5400 2417.3400 2276.1400 2417.8200 ;
        RECT 2274.5400 2422.7800 2276.1400 2423.2600 ;
        RECT 2274.5400 2428.2200 2276.1400 2428.7000 ;
        RECT 2229.5400 2433.6600 2231.1400 2434.1400 ;
        RECT 2229.5400 2439.1000 2231.1400 2439.5800 ;
        RECT 2229.5400 2417.3400 2231.1400 2417.8200 ;
        RECT 2229.5400 2422.7800 2231.1400 2423.2600 ;
        RECT 2229.5400 2428.2200 2231.1400 2428.7000 ;
        RECT 2184.5400 2444.5400 2186.1400 2445.0200 ;
        RECT 2184.5400 2449.9800 2186.1400 2450.4600 ;
        RECT 2176.7800 2444.5400 2178.3800 2445.0200 ;
        RECT 2176.7800 2449.9800 2178.3800 2450.4600 ;
        RECT 2176.7800 2455.4200 2178.3800 2455.9000 ;
        RECT 2184.5400 2455.4200 2186.1400 2455.9000 ;
        RECT 2184.5400 2433.6600 2186.1400 2434.1400 ;
        RECT 2184.5400 2439.1000 2186.1400 2439.5800 ;
        RECT 2176.7800 2433.6600 2178.3800 2434.1400 ;
        RECT 2176.7800 2439.1000 2178.3800 2439.5800 ;
        RECT 2184.5400 2417.3400 2186.1400 2417.8200 ;
        RECT 2184.5400 2422.7800 2186.1400 2423.2600 ;
        RECT 2176.7800 2417.3400 2178.3800 2417.8200 ;
        RECT 2176.7800 2422.7800 2178.3800 2423.2600 ;
        RECT 2176.7800 2428.2200 2178.3800 2428.7000 ;
        RECT 2184.5400 2428.2200 2186.1400 2428.7000 ;
        RECT 2274.5400 2401.0200 2276.1400 2401.5000 ;
        RECT 2274.5400 2406.4600 2276.1400 2406.9400 ;
        RECT 2274.5400 2411.9000 2276.1400 2412.3800 ;
        RECT 2274.5400 2390.1400 2276.1400 2390.6200 ;
        RECT 2274.5400 2395.5800 2276.1400 2396.0600 ;
        RECT 2229.5400 2401.0200 2231.1400 2401.5000 ;
        RECT 2229.5400 2406.4600 2231.1400 2406.9400 ;
        RECT 2229.5400 2411.9000 2231.1400 2412.3800 ;
        RECT 2229.5400 2390.1400 2231.1400 2390.6200 ;
        RECT 2229.5400 2395.5800 2231.1400 2396.0600 ;
        RECT 2274.5400 2373.8200 2276.1400 2374.3000 ;
        RECT 2274.5400 2379.2600 2276.1400 2379.7400 ;
        RECT 2274.5400 2384.7000 2276.1400 2385.1800 ;
        RECT 2274.5400 2362.9400 2276.1400 2363.4200 ;
        RECT 2274.5400 2368.3800 2276.1400 2368.8600 ;
        RECT 2229.5400 2373.8200 2231.1400 2374.3000 ;
        RECT 2229.5400 2379.2600 2231.1400 2379.7400 ;
        RECT 2229.5400 2384.7000 2231.1400 2385.1800 ;
        RECT 2229.5400 2362.9400 2231.1400 2363.4200 ;
        RECT 2229.5400 2368.3800 2231.1400 2368.8600 ;
        RECT 2184.5400 2401.0200 2186.1400 2401.5000 ;
        RECT 2184.5400 2406.4600 2186.1400 2406.9400 ;
        RECT 2184.5400 2411.9000 2186.1400 2412.3800 ;
        RECT 2176.7800 2401.0200 2178.3800 2401.5000 ;
        RECT 2176.7800 2406.4600 2178.3800 2406.9400 ;
        RECT 2176.7800 2411.9000 2178.3800 2412.3800 ;
        RECT 2184.5400 2390.1400 2186.1400 2390.6200 ;
        RECT 2184.5400 2395.5800 2186.1400 2396.0600 ;
        RECT 2176.7800 2390.1400 2178.3800 2390.6200 ;
        RECT 2176.7800 2395.5800 2178.3800 2396.0600 ;
        RECT 2184.5400 2373.8200 2186.1400 2374.3000 ;
        RECT 2184.5400 2379.2600 2186.1400 2379.7400 ;
        RECT 2184.5400 2384.7000 2186.1400 2385.1800 ;
        RECT 2176.7800 2373.8200 2178.3800 2374.3000 ;
        RECT 2176.7800 2379.2600 2178.3800 2379.7400 ;
        RECT 2176.7800 2384.7000 2178.3800 2385.1800 ;
        RECT 2184.5400 2362.9400 2186.1400 2363.4200 ;
        RECT 2184.5400 2368.3800 2186.1400 2368.8600 ;
        RECT 2176.7800 2362.9400 2178.3800 2363.4200 ;
        RECT 2176.7800 2368.3800 2178.3800 2368.8600 ;
        RECT 2374.2800 2346.6200 2375.8800 2347.1000 ;
        RECT 2374.2800 2352.0600 2375.8800 2352.5400 ;
        RECT 2374.2800 2357.5000 2375.8800 2357.9800 ;
        RECT 2364.5400 2346.6200 2366.1400 2347.1000 ;
        RECT 2364.5400 2352.0600 2366.1400 2352.5400 ;
        RECT 2364.5400 2357.5000 2366.1400 2357.9800 ;
        RECT 2374.2800 2335.7400 2375.8800 2336.2200 ;
        RECT 2374.2800 2341.1800 2375.8800 2341.6600 ;
        RECT 2364.5400 2335.7400 2366.1400 2336.2200 ;
        RECT 2364.5400 2341.1800 2366.1400 2341.6600 ;
        RECT 2374.2800 2319.4200 2375.8800 2319.9000 ;
        RECT 2374.2800 2324.8600 2375.8800 2325.3400 ;
        RECT 2374.2800 2330.3000 2375.8800 2330.7800 ;
        RECT 2364.5400 2319.4200 2366.1400 2319.9000 ;
        RECT 2364.5400 2324.8600 2366.1400 2325.3400 ;
        RECT 2364.5400 2330.3000 2366.1400 2330.7800 ;
        RECT 2374.2800 2308.5400 2375.8800 2309.0200 ;
        RECT 2374.2800 2313.9800 2375.8800 2314.4600 ;
        RECT 2364.5400 2308.5400 2366.1400 2309.0200 ;
        RECT 2364.5400 2313.9800 2366.1400 2314.4600 ;
        RECT 2319.5400 2346.6200 2321.1400 2347.1000 ;
        RECT 2319.5400 2352.0600 2321.1400 2352.5400 ;
        RECT 2319.5400 2357.5000 2321.1400 2357.9800 ;
        RECT 2319.5400 2335.7400 2321.1400 2336.2200 ;
        RECT 2319.5400 2341.1800 2321.1400 2341.6600 ;
        RECT 2319.5400 2319.4200 2321.1400 2319.9000 ;
        RECT 2319.5400 2324.8600 2321.1400 2325.3400 ;
        RECT 2319.5400 2330.3000 2321.1400 2330.7800 ;
        RECT 2319.5400 2308.5400 2321.1400 2309.0200 ;
        RECT 2319.5400 2313.9800 2321.1400 2314.4600 ;
        RECT 2374.2800 2292.2200 2375.8800 2292.7000 ;
        RECT 2374.2800 2297.6600 2375.8800 2298.1400 ;
        RECT 2374.2800 2303.1000 2375.8800 2303.5800 ;
        RECT 2364.5400 2292.2200 2366.1400 2292.7000 ;
        RECT 2364.5400 2297.6600 2366.1400 2298.1400 ;
        RECT 2364.5400 2303.1000 2366.1400 2303.5800 ;
        RECT 2374.2800 2281.3400 2375.8800 2281.8200 ;
        RECT 2374.2800 2286.7800 2375.8800 2287.2600 ;
        RECT 2364.5400 2281.3400 2366.1400 2281.8200 ;
        RECT 2364.5400 2286.7800 2366.1400 2287.2600 ;
        RECT 2374.2800 2265.0200 2375.8800 2265.5000 ;
        RECT 2374.2800 2270.4600 2375.8800 2270.9400 ;
        RECT 2374.2800 2275.9000 2375.8800 2276.3800 ;
        RECT 2364.5400 2265.0200 2366.1400 2265.5000 ;
        RECT 2364.5400 2270.4600 2366.1400 2270.9400 ;
        RECT 2364.5400 2275.9000 2366.1400 2276.3800 ;
        RECT 2364.5400 2259.5800 2366.1400 2260.0600 ;
        RECT 2374.2800 2259.5800 2375.8800 2260.0600 ;
        RECT 2319.5400 2292.2200 2321.1400 2292.7000 ;
        RECT 2319.5400 2297.6600 2321.1400 2298.1400 ;
        RECT 2319.5400 2303.1000 2321.1400 2303.5800 ;
        RECT 2319.5400 2281.3400 2321.1400 2281.8200 ;
        RECT 2319.5400 2286.7800 2321.1400 2287.2600 ;
        RECT 2319.5400 2265.0200 2321.1400 2265.5000 ;
        RECT 2319.5400 2270.4600 2321.1400 2270.9400 ;
        RECT 2319.5400 2275.9000 2321.1400 2276.3800 ;
        RECT 2319.5400 2259.5800 2321.1400 2260.0600 ;
        RECT 2274.5400 2346.6200 2276.1400 2347.1000 ;
        RECT 2274.5400 2352.0600 2276.1400 2352.5400 ;
        RECT 2274.5400 2357.5000 2276.1400 2357.9800 ;
        RECT 2274.5400 2335.7400 2276.1400 2336.2200 ;
        RECT 2274.5400 2341.1800 2276.1400 2341.6600 ;
        RECT 2229.5400 2346.6200 2231.1400 2347.1000 ;
        RECT 2229.5400 2352.0600 2231.1400 2352.5400 ;
        RECT 2229.5400 2357.5000 2231.1400 2357.9800 ;
        RECT 2229.5400 2335.7400 2231.1400 2336.2200 ;
        RECT 2229.5400 2341.1800 2231.1400 2341.6600 ;
        RECT 2274.5400 2319.4200 2276.1400 2319.9000 ;
        RECT 2274.5400 2324.8600 2276.1400 2325.3400 ;
        RECT 2274.5400 2330.3000 2276.1400 2330.7800 ;
        RECT 2274.5400 2308.5400 2276.1400 2309.0200 ;
        RECT 2274.5400 2313.9800 2276.1400 2314.4600 ;
        RECT 2229.5400 2319.4200 2231.1400 2319.9000 ;
        RECT 2229.5400 2324.8600 2231.1400 2325.3400 ;
        RECT 2229.5400 2330.3000 2231.1400 2330.7800 ;
        RECT 2229.5400 2308.5400 2231.1400 2309.0200 ;
        RECT 2229.5400 2313.9800 2231.1400 2314.4600 ;
        RECT 2184.5400 2346.6200 2186.1400 2347.1000 ;
        RECT 2184.5400 2352.0600 2186.1400 2352.5400 ;
        RECT 2184.5400 2357.5000 2186.1400 2357.9800 ;
        RECT 2176.7800 2346.6200 2178.3800 2347.1000 ;
        RECT 2176.7800 2352.0600 2178.3800 2352.5400 ;
        RECT 2176.7800 2357.5000 2178.3800 2357.9800 ;
        RECT 2184.5400 2335.7400 2186.1400 2336.2200 ;
        RECT 2184.5400 2341.1800 2186.1400 2341.6600 ;
        RECT 2176.7800 2335.7400 2178.3800 2336.2200 ;
        RECT 2176.7800 2341.1800 2178.3800 2341.6600 ;
        RECT 2184.5400 2319.4200 2186.1400 2319.9000 ;
        RECT 2184.5400 2324.8600 2186.1400 2325.3400 ;
        RECT 2184.5400 2330.3000 2186.1400 2330.7800 ;
        RECT 2176.7800 2319.4200 2178.3800 2319.9000 ;
        RECT 2176.7800 2324.8600 2178.3800 2325.3400 ;
        RECT 2176.7800 2330.3000 2178.3800 2330.7800 ;
        RECT 2184.5400 2308.5400 2186.1400 2309.0200 ;
        RECT 2184.5400 2313.9800 2186.1400 2314.4600 ;
        RECT 2176.7800 2308.5400 2178.3800 2309.0200 ;
        RECT 2176.7800 2313.9800 2178.3800 2314.4600 ;
        RECT 2274.5400 2292.2200 2276.1400 2292.7000 ;
        RECT 2274.5400 2297.6600 2276.1400 2298.1400 ;
        RECT 2274.5400 2303.1000 2276.1400 2303.5800 ;
        RECT 2274.5400 2281.3400 2276.1400 2281.8200 ;
        RECT 2274.5400 2286.7800 2276.1400 2287.2600 ;
        RECT 2229.5400 2292.2200 2231.1400 2292.7000 ;
        RECT 2229.5400 2297.6600 2231.1400 2298.1400 ;
        RECT 2229.5400 2303.1000 2231.1400 2303.5800 ;
        RECT 2229.5400 2281.3400 2231.1400 2281.8200 ;
        RECT 2229.5400 2286.7800 2231.1400 2287.2600 ;
        RECT 2274.5400 2265.0200 2276.1400 2265.5000 ;
        RECT 2274.5400 2270.4600 2276.1400 2270.9400 ;
        RECT 2274.5400 2275.9000 2276.1400 2276.3800 ;
        RECT 2274.5400 2259.5800 2276.1400 2260.0600 ;
        RECT 2229.5400 2265.0200 2231.1400 2265.5000 ;
        RECT 2229.5400 2270.4600 2231.1400 2270.9400 ;
        RECT 2229.5400 2275.9000 2231.1400 2276.3800 ;
        RECT 2229.5400 2259.5800 2231.1400 2260.0600 ;
        RECT 2184.5400 2292.2200 2186.1400 2292.7000 ;
        RECT 2184.5400 2297.6600 2186.1400 2298.1400 ;
        RECT 2184.5400 2303.1000 2186.1400 2303.5800 ;
        RECT 2176.7800 2292.2200 2178.3800 2292.7000 ;
        RECT 2176.7800 2297.6600 2178.3800 2298.1400 ;
        RECT 2176.7800 2303.1000 2178.3800 2303.5800 ;
        RECT 2184.5400 2281.3400 2186.1400 2281.8200 ;
        RECT 2184.5400 2286.7800 2186.1400 2287.2600 ;
        RECT 2176.7800 2281.3400 2178.3800 2281.8200 ;
        RECT 2176.7800 2286.7800 2178.3800 2287.2600 ;
        RECT 2184.5400 2265.0200 2186.1400 2265.5000 ;
        RECT 2184.5400 2270.4600 2186.1400 2270.9400 ;
        RECT 2184.5400 2275.9000 2186.1400 2276.3800 ;
        RECT 2176.7800 2265.0200 2178.3800 2265.5000 ;
        RECT 2176.7800 2270.4600 2178.3800 2270.9400 ;
        RECT 2176.7800 2275.9000 2178.3800 2276.3800 ;
        RECT 2176.7800 2259.5800 2178.3800 2260.0600 ;
        RECT 2184.5400 2259.5800 2186.1400 2260.0600 ;
        RECT 2171.2200 2461.8900 2381.4400 2463.4900 ;
        RECT 2171.2200 2255.3900 2381.4400 2256.9900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 2249.9600 2178.3800 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 2468.0000 2178.3800 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 2249.9600 2375.8800 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 2468.0000 2375.8800 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2255.3900 2172.8200 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2255.3900 2381.4400 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2461.8900 2172.8200 2463.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2461.8900 2381.4400 2463.4900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 2025.7500 2366.1400 2233.8500 ;
        RECT 2319.5400 2025.7500 2321.1400 2233.8500 ;
        RECT 2274.5400 2025.7500 2276.1400 2233.8500 ;
        RECT 2229.5400 2025.7500 2231.1400 2233.8500 ;
        RECT 2184.5400 2025.7500 2186.1400 2233.8500 ;
        RECT 2374.2800 2020.3200 2375.8800 2239.9600 ;
        RECT 2176.7800 2020.3200 2178.3800 2239.9600 ;
      LAYER met3 ;
        RECT 2374.2800 2214.9000 2375.8800 2215.3800 ;
        RECT 2374.2800 2220.3400 2375.8800 2220.8200 ;
        RECT 2364.5400 2214.9000 2366.1400 2215.3800 ;
        RECT 2364.5400 2220.3400 2366.1400 2220.8200 ;
        RECT 2364.5400 2225.7800 2366.1400 2226.2600 ;
        RECT 2374.2800 2225.7800 2375.8800 2226.2600 ;
        RECT 2374.2800 2204.0200 2375.8800 2204.5000 ;
        RECT 2374.2800 2209.4600 2375.8800 2209.9400 ;
        RECT 2364.5400 2204.0200 2366.1400 2204.5000 ;
        RECT 2364.5400 2209.4600 2366.1400 2209.9400 ;
        RECT 2374.2800 2187.7000 2375.8800 2188.1800 ;
        RECT 2374.2800 2193.1400 2375.8800 2193.6200 ;
        RECT 2364.5400 2187.7000 2366.1400 2188.1800 ;
        RECT 2364.5400 2193.1400 2366.1400 2193.6200 ;
        RECT 2364.5400 2198.5800 2366.1400 2199.0600 ;
        RECT 2374.2800 2198.5800 2375.8800 2199.0600 ;
        RECT 2319.5400 2214.9000 2321.1400 2215.3800 ;
        RECT 2319.5400 2220.3400 2321.1400 2220.8200 ;
        RECT 2319.5400 2225.7800 2321.1400 2226.2600 ;
        RECT 2319.5400 2204.0200 2321.1400 2204.5000 ;
        RECT 2319.5400 2209.4600 2321.1400 2209.9400 ;
        RECT 2319.5400 2187.7000 2321.1400 2188.1800 ;
        RECT 2319.5400 2193.1400 2321.1400 2193.6200 ;
        RECT 2319.5400 2198.5800 2321.1400 2199.0600 ;
        RECT 2374.2800 2171.3800 2375.8800 2171.8600 ;
        RECT 2374.2800 2176.8200 2375.8800 2177.3000 ;
        RECT 2374.2800 2182.2600 2375.8800 2182.7400 ;
        RECT 2364.5400 2171.3800 2366.1400 2171.8600 ;
        RECT 2364.5400 2176.8200 2366.1400 2177.3000 ;
        RECT 2364.5400 2182.2600 2366.1400 2182.7400 ;
        RECT 2374.2800 2160.5000 2375.8800 2160.9800 ;
        RECT 2374.2800 2165.9400 2375.8800 2166.4200 ;
        RECT 2364.5400 2160.5000 2366.1400 2160.9800 ;
        RECT 2364.5400 2165.9400 2366.1400 2166.4200 ;
        RECT 2374.2800 2144.1800 2375.8800 2144.6600 ;
        RECT 2374.2800 2149.6200 2375.8800 2150.1000 ;
        RECT 2374.2800 2155.0600 2375.8800 2155.5400 ;
        RECT 2364.5400 2144.1800 2366.1400 2144.6600 ;
        RECT 2364.5400 2149.6200 2366.1400 2150.1000 ;
        RECT 2364.5400 2155.0600 2366.1400 2155.5400 ;
        RECT 2374.2800 2133.3000 2375.8800 2133.7800 ;
        RECT 2374.2800 2138.7400 2375.8800 2139.2200 ;
        RECT 2364.5400 2133.3000 2366.1400 2133.7800 ;
        RECT 2364.5400 2138.7400 2366.1400 2139.2200 ;
        RECT 2319.5400 2171.3800 2321.1400 2171.8600 ;
        RECT 2319.5400 2176.8200 2321.1400 2177.3000 ;
        RECT 2319.5400 2182.2600 2321.1400 2182.7400 ;
        RECT 2319.5400 2160.5000 2321.1400 2160.9800 ;
        RECT 2319.5400 2165.9400 2321.1400 2166.4200 ;
        RECT 2319.5400 2144.1800 2321.1400 2144.6600 ;
        RECT 2319.5400 2149.6200 2321.1400 2150.1000 ;
        RECT 2319.5400 2155.0600 2321.1400 2155.5400 ;
        RECT 2319.5400 2133.3000 2321.1400 2133.7800 ;
        RECT 2319.5400 2138.7400 2321.1400 2139.2200 ;
        RECT 2274.5400 2214.9000 2276.1400 2215.3800 ;
        RECT 2274.5400 2220.3400 2276.1400 2220.8200 ;
        RECT 2274.5400 2225.7800 2276.1400 2226.2600 ;
        RECT 2229.5400 2214.9000 2231.1400 2215.3800 ;
        RECT 2229.5400 2220.3400 2231.1400 2220.8200 ;
        RECT 2229.5400 2225.7800 2231.1400 2226.2600 ;
        RECT 2274.5400 2204.0200 2276.1400 2204.5000 ;
        RECT 2274.5400 2209.4600 2276.1400 2209.9400 ;
        RECT 2274.5400 2187.7000 2276.1400 2188.1800 ;
        RECT 2274.5400 2193.1400 2276.1400 2193.6200 ;
        RECT 2274.5400 2198.5800 2276.1400 2199.0600 ;
        RECT 2229.5400 2204.0200 2231.1400 2204.5000 ;
        RECT 2229.5400 2209.4600 2231.1400 2209.9400 ;
        RECT 2229.5400 2187.7000 2231.1400 2188.1800 ;
        RECT 2229.5400 2193.1400 2231.1400 2193.6200 ;
        RECT 2229.5400 2198.5800 2231.1400 2199.0600 ;
        RECT 2184.5400 2214.9000 2186.1400 2215.3800 ;
        RECT 2184.5400 2220.3400 2186.1400 2220.8200 ;
        RECT 2176.7800 2214.9000 2178.3800 2215.3800 ;
        RECT 2176.7800 2220.3400 2178.3800 2220.8200 ;
        RECT 2176.7800 2225.7800 2178.3800 2226.2600 ;
        RECT 2184.5400 2225.7800 2186.1400 2226.2600 ;
        RECT 2184.5400 2204.0200 2186.1400 2204.5000 ;
        RECT 2184.5400 2209.4600 2186.1400 2209.9400 ;
        RECT 2176.7800 2204.0200 2178.3800 2204.5000 ;
        RECT 2176.7800 2209.4600 2178.3800 2209.9400 ;
        RECT 2184.5400 2187.7000 2186.1400 2188.1800 ;
        RECT 2184.5400 2193.1400 2186.1400 2193.6200 ;
        RECT 2176.7800 2187.7000 2178.3800 2188.1800 ;
        RECT 2176.7800 2193.1400 2178.3800 2193.6200 ;
        RECT 2176.7800 2198.5800 2178.3800 2199.0600 ;
        RECT 2184.5400 2198.5800 2186.1400 2199.0600 ;
        RECT 2274.5400 2171.3800 2276.1400 2171.8600 ;
        RECT 2274.5400 2176.8200 2276.1400 2177.3000 ;
        RECT 2274.5400 2182.2600 2276.1400 2182.7400 ;
        RECT 2274.5400 2160.5000 2276.1400 2160.9800 ;
        RECT 2274.5400 2165.9400 2276.1400 2166.4200 ;
        RECT 2229.5400 2171.3800 2231.1400 2171.8600 ;
        RECT 2229.5400 2176.8200 2231.1400 2177.3000 ;
        RECT 2229.5400 2182.2600 2231.1400 2182.7400 ;
        RECT 2229.5400 2160.5000 2231.1400 2160.9800 ;
        RECT 2229.5400 2165.9400 2231.1400 2166.4200 ;
        RECT 2274.5400 2144.1800 2276.1400 2144.6600 ;
        RECT 2274.5400 2149.6200 2276.1400 2150.1000 ;
        RECT 2274.5400 2155.0600 2276.1400 2155.5400 ;
        RECT 2274.5400 2133.3000 2276.1400 2133.7800 ;
        RECT 2274.5400 2138.7400 2276.1400 2139.2200 ;
        RECT 2229.5400 2144.1800 2231.1400 2144.6600 ;
        RECT 2229.5400 2149.6200 2231.1400 2150.1000 ;
        RECT 2229.5400 2155.0600 2231.1400 2155.5400 ;
        RECT 2229.5400 2133.3000 2231.1400 2133.7800 ;
        RECT 2229.5400 2138.7400 2231.1400 2139.2200 ;
        RECT 2184.5400 2171.3800 2186.1400 2171.8600 ;
        RECT 2184.5400 2176.8200 2186.1400 2177.3000 ;
        RECT 2184.5400 2182.2600 2186.1400 2182.7400 ;
        RECT 2176.7800 2171.3800 2178.3800 2171.8600 ;
        RECT 2176.7800 2176.8200 2178.3800 2177.3000 ;
        RECT 2176.7800 2182.2600 2178.3800 2182.7400 ;
        RECT 2184.5400 2160.5000 2186.1400 2160.9800 ;
        RECT 2184.5400 2165.9400 2186.1400 2166.4200 ;
        RECT 2176.7800 2160.5000 2178.3800 2160.9800 ;
        RECT 2176.7800 2165.9400 2178.3800 2166.4200 ;
        RECT 2184.5400 2144.1800 2186.1400 2144.6600 ;
        RECT 2184.5400 2149.6200 2186.1400 2150.1000 ;
        RECT 2184.5400 2155.0600 2186.1400 2155.5400 ;
        RECT 2176.7800 2144.1800 2178.3800 2144.6600 ;
        RECT 2176.7800 2149.6200 2178.3800 2150.1000 ;
        RECT 2176.7800 2155.0600 2178.3800 2155.5400 ;
        RECT 2184.5400 2133.3000 2186.1400 2133.7800 ;
        RECT 2184.5400 2138.7400 2186.1400 2139.2200 ;
        RECT 2176.7800 2133.3000 2178.3800 2133.7800 ;
        RECT 2176.7800 2138.7400 2178.3800 2139.2200 ;
        RECT 2374.2800 2116.9800 2375.8800 2117.4600 ;
        RECT 2374.2800 2122.4200 2375.8800 2122.9000 ;
        RECT 2374.2800 2127.8600 2375.8800 2128.3400 ;
        RECT 2364.5400 2116.9800 2366.1400 2117.4600 ;
        RECT 2364.5400 2122.4200 2366.1400 2122.9000 ;
        RECT 2364.5400 2127.8600 2366.1400 2128.3400 ;
        RECT 2374.2800 2106.1000 2375.8800 2106.5800 ;
        RECT 2374.2800 2111.5400 2375.8800 2112.0200 ;
        RECT 2364.5400 2106.1000 2366.1400 2106.5800 ;
        RECT 2364.5400 2111.5400 2366.1400 2112.0200 ;
        RECT 2374.2800 2089.7800 2375.8800 2090.2600 ;
        RECT 2374.2800 2095.2200 2375.8800 2095.7000 ;
        RECT 2374.2800 2100.6600 2375.8800 2101.1400 ;
        RECT 2364.5400 2089.7800 2366.1400 2090.2600 ;
        RECT 2364.5400 2095.2200 2366.1400 2095.7000 ;
        RECT 2364.5400 2100.6600 2366.1400 2101.1400 ;
        RECT 2374.2800 2078.9000 2375.8800 2079.3800 ;
        RECT 2374.2800 2084.3400 2375.8800 2084.8200 ;
        RECT 2364.5400 2078.9000 2366.1400 2079.3800 ;
        RECT 2364.5400 2084.3400 2366.1400 2084.8200 ;
        RECT 2319.5400 2116.9800 2321.1400 2117.4600 ;
        RECT 2319.5400 2122.4200 2321.1400 2122.9000 ;
        RECT 2319.5400 2127.8600 2321.1400 2128.3400 ;
        RECT 2319.5400 2106.1000 2321.1400 2106.5800 ;
        RECT 2319.5400 2111.5400 2321.1400 2112.0200 ;
        RECT 2319.5400 2089.7800 2321.1400 2090.2600 ;
        RECT 2319.5400 2095.2200 2321.1400 2095.7000 ;
        RECT 2319.5400 2100.6600 2321.1400 2101.1400 ;
        RECT 2319.5400 2078.9000 2321.1400 2079.3800 ;
        RECT 2319.5400 2084.3400 2321.1400 2084.8200 ;
        RECT 2374.2800 2062.5800 2375.8800 2063.0600 ;
        RECT 2374.2800 2068.0200 2375.8800 2068.5000 ;
        RECT 2374.2800 2073.4600 2375.8800 2073.9400 ;
        RECT 2364.5400 2062.5800 2366.1400 2063.0600 ;
        RECT 2364.5400 2068.0200 2366.1400 2068.5000 ;
        RECT 2364.5400 2073.4600 2366.1400 2073.9400 ;
        RECT 2374.2800 2051.7000 2375.8800 2052.1800 ;
        RECT 2374.2800 2057.1400 2375.8800 2057.6200 ;
        RECT 2364.5400 2051.7000 2366.1400 2052.1800 ;
        RECT 2364.5400 2057.1400 2366.1400 2057.6200 ;
        RECT 2374.2800 2035.3800 2375.8800 2035.8600 ;
        RECT 2374.2800 2040.8200 2375.8800 2041.3000 ;
        RECT 2374.2800 2046.2600 2375.8800 2046.7400 ;
        RECT 2364.5400 2035.3800 2366.1400 2035.8600 ;
        RECT 2364.5400 2040.8200 2366.1400 2041.3000 ;
        RECT 2364.5400 2046.2600 2366.1400 2046.7400 ;
        RECT 2364.5400 2029.9400 2366.1400 2030.4200 ;
        RECT 2374.2800 2029.9400 2375.8800 2030.4200 ;
        RECT 2319.5400 2062.5800 2321.1400 2063.0600 ;
        RECT 2319.5400 2068.0200 2321.1400 2068.5000 ;
        RECT 2319.5400 2073.4600 2321.1400 2073.9400 ;
        RECT 2319.5400 2051.7000 2321.1400 2052.1800 ;
        RECT 2319.5400 2057.1400 2321.1400 2057.6200 ;
        RECT 2319.5400 2035.3800 2321.1400 2035.8600 ;
        RECT 2319.5400 2040.8200 2321.1400 2041.3000 ;
        RECT 2319.5400 2046.2600 2321.1400 2046.7400 ;
        RECT 2319.5400 2029.9400 2321.1400 2030.4200 ;
        RECT 2274.5400 2116.9800 2276.1400 2117.4600 ;
        RECT 2274.5400 2122.4200 2276.1400 2122.9000 ;
        RECT 2274.5400 2127.8600 2276.1400 2128.3400 ;
        RECT 2274.5400 2106.1000 2276.1400 2106.5800 ;
        RECT 2274.5400 2111.5400 2276.1400 2112.0200 ;
        RECT 2229.5400 2116.9800 2231.1400 2117.4600 ;
        RECT 2229.5400 2122.4200 2231.1400 2122.9000 ;
        RECT 2229.5400 2127.8600 2231.1400 2128.3400 ;
        RECT 2229.5400 2106.1000 2231.1400 2106.5800 ;
        RECT 2229.5400 2111.5400 2231.1400 2112.0200 ;
        RECT 2274.5400 2089.7800 2276.1400 2090.2600 ;
        RECT 2274.5400 2095.2200 2276.1400 2095.7000 ;
        RECT 2274.5400 2100.6600 2276.1400 2101.1400 ;
        RECT 2274.5400 2078.9000 2276.1400 2079.3800 ;
        RECT 2274.5400 2084.3400 2276.1400 2084.8200 ;
        RECT 2229.5400 2089.7800 2231.1400 2090.2600 ;
        RECT 2229.5400 2095.2200 2231.1400 2095.7000 ;
        RECT 2229.5400 2100.6600 2231.1400 2101.1400 ;
        RECT 2229.5400 2078.9000 2231.1400 2079.3800 ;
        RECT 2229.5400 2084.3400 2231.1400 2084.8200 ;
        RECT 2184.5400 2116.9800 2186.1400 2117.4600 ;
        RECT 2184.5400 2122.4200 2186.1400 2122.9000 ;
        RECT 2184.5400 2127.8600 2186.1400 2128.3400 ;
        RECT 2176.7800 2116.9800 2178.3800 2117.4600 ;
        RECT 2176.7800 2122.4200 2178.3800 2122.9000 ;
        RECT 2176.7800 2127.8600 2178.3800 2128.3400 ;
        RECT 2184.5400 2106.1000 2186.1400 2106.5800 ;
        RECT 2184.5400 2111.5400 2186.1400 2112.0200 ;
        RECT 2176.7800 2106.1000 2178.3800 2106.5800 ;
        RECT 2176.7800 2111.5400 2178.3800 2112.0200 ;
        RECT 2184.5400 2089.7800 2186.1400 2090.2600 ;
        RECT 2184.5400 2095.2200 2186.1400 2095.7000 ;
        RECT 2184.5400 2100.6600 2186.1400 2101.1400 ;
        RECT 2176.7800 2089.7800 2178.3800 2090.2600 ;
        RECT 2176.7800 2095.2200 2178.3800 2095.7000 ;
        RECT 2176.7800 2100.6600 2178.3800 2101.1400 ;
        RECT 2184.5400 2078.9000 2186.1400 2079.3800 ;
        RECT 2184.5400 2084.3400 2186.1400 2084.8200 ;
        RECT 2176.7800 2078.9000 2178.3800 2079.3800 ;
        RECT 2176.7800 2084.3400 2178.3800 2084.8200 ;
        RECT 2274.5400 2062.5800 2276.1400 2063.0600 ;
        RECT 2274.5400 2068.0200 2276.1400 2068.5000 ;
        RECT 2274.5400 2073.4600 2276.1400 2073.9400 ;
        RECT 2274.5400 2051.7000 2276.1400 2052.1800 ;
        RECT 2274.5400 2057.1400 2276.1400 2057.6200 ;
        RECT 2229.5400 2062.5800 2231.1400 2063.0600 ;
        RECT 2229.5400 2068.0200 2231.1400 2068.5000 ;
        RECT 2229.5400 2073.4600 2231.1400 2073.9400 ;
        RECT 2229.5400 2051.7000 2231.1400 2052.1800 ;
        RECT 2229.5400 2057.1400 2231.1400 2057.6200 ;
        RECT 2274.5400 2035.3800 2276.1400 2035.8600 ;
        RECT 2274.5400 2040.8200 2276.1400 2041.3000 ;
        RECT 2274.5400 2046.2600 2276.1400 2046.7400 ;
        RECT 2274.5400 2029.9400 2276.1400 2030.4200 ;
        RECT 2229.5400 2035.3800 2231.1400 2035.8600 ;
        RECT 2229.5400 2040.8200 2231.1400 2041.3000 ;
        RECT 2229.5400 2046.2600 2231.1400 2046.7400 ;
        RECT 2229.5400 2029.9400 2231.1400 2030.4200 ;
        RECT 2184.5400 2062.5800 2186.1400 2063.0600 ;
        RECT 2184.5400 2068.0200 2186.1400 2068.5000 ;
        RECT 2184.5400 2073.4600 2186.1400 2073.9400 ;
        RECT 2176.7800 2062.5800 2178.3800 2063.0600 ;
        RECT 2176.7800 2068.0200 2178.3800 2068.5000 ;
        RECT 2176.7800 2073.4600 2178.3800 2073.9400 ;
        RECT 2184.5400 2051.7000 2186.1400 2052.1800 ;
        RECT 2184.5400 2057.1400 2186.1400 2057.6200 ;
        RECT 2176.7800 2051.7000 2178.3800 2052.1800 ;
        RECT 2176.7800 2057.1400 2178.3800 2057.6200 ;
        RECT 2184.5400 2035.3800 2186.1400 2035.8600 ;
        RECT 2184.5400 2040.8200 2186.1400 2041.3000 ;
        RECT 2184.5400 2046.2600 2186.1400 2046.7400 ;
        RECT 2176.7800 2035.3800 2178.3800 2035.8600 ;
        RECT 2176.7800 2040.8200 2178.3800 2041.3000 ;
        RECT 2176.7800 2046.2600 2178.3800 2046.7400 ;
        RECT 2176.7800 2029.9400 2178.3800 2030.4200 ;
        RECT 2184.5400 2029.9400 2186.1400 2030.4200 ;
        RECT 2171.2200 2232.2500 2381.4400 2233.8500 ;
        RECT 2171.2200 2025.7500 2381.4400 2027.3500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 2020.3200 2178.3800 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 2238.3600 2178.3800 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 2020.3200 2375.8800 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 2238.3600 2375.8800 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2025.7500 2172.8200 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2025.7500 2381.4400 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2232.2500 2172.8200 2233.8500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2232.2500 2381.4400 2233.8500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 1796.1100 2366.1400 2004.2100 ;
        RECT 2319.5400 1796.1100 2321.1400 2004.2100 ;
        RECT 2274.5400 1796.1100 2276.1400 2004.2100 ;
        RECT 2229.5400 1796.1100 2231.1400 2004.2100 ;
        RECT 2184.5400 1796.1100 2186.1400 2004.2100 ;
        RECT 2374.2800 1790.6800 2375.8800 2010.3200 ;
        RECT 2176.7800 1790.6800 2178.3800 2010.3200 ;
      LAYER met3 ;
        RECT 2374.2800 1985.2600 2375.8800 1985.7400 ;
        RECT 2374.2800 1990.7000 2375.8800 1991.1800 ;
        RECT 2364.5400 1985.2600 2366.1400 1985.7400 ;
        RECT 2364.5400 1990.7000 2366.1400 1991.1800 ;
        RECT 2364.5400 1996.1400 2366.1400 1996.6200 ;
        RECT 2374.2800 1996.1400 2375.8800 1996.6200 ;
        RECT 2374.2800 1974.3800 2375.8800 1974.8600 ;
        RECT 2374.2800 1979.8200 2375.8800 1980.3000 ;
        RECT 2364.5400 1974.3800 2366.1400 1974.8600 ;
        RECT 2364.5400 1979.8200 2366.1400 1980.3000 ;
        RECT 2374.2800 1958.0600 2375.8800 1958.5400 ;
        RECT 2374.2800 1963.5000 2375.8800 1963.9800 ;
        RECT 2364.5400 1958.0600 2366.1400 1958.5400 ;
        RECT 2364.5400 1963.5000 2366.1400 1963.9800 ;
        RECT 2364.5400 1968.9400 2366.1400 1969.4200 ;
        RECT 2374.2800 1968.9400 2375.8800 1969.4200 ;
        RECT 2319.5400 1985.2600 2321.1400 1985.7400 ;
        RECT 2319.5400 1990.7000 2321.1400 1991.1800 ;
        RECT 2319.5400 1996.1400 2321.1400 1996.6200 ;
        RECT 2319.5400 1974.3800 2321.1400 1974.8600 ;
        RECT 2319.5400 1979.8200 2321.1400 1980.3000 ;
        RECT 2319.5400 1958.0600 2321.1400 1958.5400 ;
        RECT 2319.5400 1963.5000 2321.1400 1963.9800 ;
        RECT 2319.5400 1968.9400 2321.1400 1969.4200 ;
        RECT 2374.2800 1941.7400 2375.8800 1942.2200 ;
        RECT 2374.2800 1947.1800 2375.8800 1947.6600 ;
        RECT 2374.2800 1952.6200 2375.8800 1953.1000 ;
        RECT 2364.5400 1941.7400 2366.1400 1942.2200 ;
        RECT 2364.5400 1947.1800 2366.1400 1947.6600 ;
        RECT 2364.5400 1952.6200 2366.1400 1953.1000 ;
        RECT 2374.2800 1930.8600 2375.8800 1931.3400 ;
        RECT 2374.2800 1936.3000 2375.8800 1936.7800 ;
        RECT 2364.5400 1930.8600 2366.1400 1931.3400 ;
        RECT 2364.5400 1936.3000 2366.1400 1936.7800 ;
        RECT 2374.2800 1914.5400 2375.8800 1915.0200 ;
        RECT 2374.2800 1919.9800 2375.8800 1920.4600 ;
        RECT 2374.2800 1925.4200 2375.8800 1925.9000 ;
        RECT 2364.5400 1914.5400 2366.1400 1915.0200 ;
        RECT 2364.5400 1919.9800 2366.1400 1920.4600 ;
        RECT 2364.5400 1925.4200 2366.1400 1925.9000 ;
        RECT 2374.2800 1903.6600 2375.8800 1904.1400 ;
        RECT 2374.2800 1909.1000 2375.8800 1909.5800 ;
        RECT 2364.5400 1903.6600 2366.1400 1904.1400 ;
        RECT 2364.5400 1909.1000 2366.1400 1909.5800 ;
        RECT 2319.5400 1941.7400 2321.1400 1942.2200 ;
        RECT 2319.5400 1947.1800 2321.1400 1947.6600 ;
        RECT 2319.5400 1952.6200 2321.1400 1953.1000 ;
        RECT 2319.5400 1930.8600 2321.1400 1931.3400 ;
        RECT 2319.5400 1936.3000 2321.1400 1936.7800 ;
        RECT 2319.5400 1914.5400 2321.1400 1915.0200 ;
        RECT 2319.5400 1919.9800 2321.1400 1920.4600 ;
        RECT 2319.5400 1925.4200 2321.1400 1925.9000 ;
        RECT 2319.5400 1903.6600 2321.1400 1904.1400 ;
        RECT 2319.5400 1909.1000 2321.1400 1909.5800 ;
        RECT 2274.5400 1985.2600 2276.1400 1985.7400 ;
        RECT 2274.5400 1990.7000 2276.1400 1991.1800 ;
        RECT 2274.5400 1996.1400 2276.1400 1996.6200 ;
        RECT 2229.5400 1985.2600 2231.1400 1985.7400 ;
        RECT 2229.5400 1990.7000 2231.1400 1991.1800 ;
        RECT 2229.5400 1996.1400 2231.1400 1996.6200 ;
        RECT 2274.5400 1974.3800 2276.1400 1974.8600 ;
        RECT 2274.5400 1979.8200 2276.1400 1980.3000 ;
        RECT 2274.5400 1958.0600 2276.1400 1958.5400 ;
        RECT 2274.5400 1963.5000 2276.1400 1963.9800 ;
        RECT 2274.5400 1968.9400 2276.1400 1969.4200 ;
        RECT 2229.5400 1974.3800 2231.1400 1974.8600 ;
        RECT 2229.5400 1979.8200 2231.1400 1980.3000 ;
        RECT 2229.5400 1958.0600 2231.1400 1958.5400 ;
        RECT 2229.5400 1963.5000 2231.1400 1963.9800 ;
        RECT 2229.5400 1968.9400 2231.1400 1969.4200 ;
        RECT 2184.5400 1985.2600 2186.1400 1985.7400 ;
        RECT 2184.5400 1990.7000 2186.1400 1991.1800 ;
        RECT 2176.7800 1985.2600 2178.3800 1985.7400 ;
        RECT 2176.7800 1990.7000 2178.3800 1991.1800 ;
        RECT 2176.7800 1996.1400 2178.3800 1996.6200 ;
        RECT 2184.5400 1996.1400 2186.1400 1996.6200 ;
        RECT 2184.5400 1974.3800 2186.1400 1974.8600 ;
        RECT 2184.5400 1979.8200 2186.1400 1980.3000 ;
        RECT 2176.7800 1974.3800 2178.3800 1974.8600 ;
        RECT 2176.7800 1979.8200 2178.3800 1980.3000 ;
        RECT 2184.5400 1958.0600 2186.1400 1958.5400 ;
        RECT 2184.5400 1963.5000 2186.1400 1963.9800 ;
        RECT 2176.7800 1958.0600 2178.3800 1958.5400 ;
        RECT 2176.7800 1963.5000 2178.3800 1963.9800 ;
        RECT 2176.7800 1968.9400 2178.3800 1969.4200 ;
        RECT 2184.5400 1968.9400 2186.1400 1969.4200 ;
        RECT 2274.5400 1941.7400 2276.1400 1942.2200 ;
        RECT 2274.5400 1947.1800 2276.1400 1947.6600 ;
        RECT 2274.5400 1952.6200 2276.1400 1953.1000 ;
        RECT 2274.5400 1930.8600 2276.1400 1931.3400 ;
        RECT 2274.5400 1936.3000 2276.1400 1936.7800 ;
        RECT 2229.5400 1941.7400 2231.1400 1942.2200 ;
        RECT 2229.5400 1947.1800 2231.1400 1947.6600 ;
        RECT 2229.5400 1952.6200 2231.1400 1953.1000 ;
        RECT 2229.5400 1930.8600 2231.1400 1931.3400 ;
        RECT 2229.5400 1936.3000 2231.1400 1936.7800 ;
        RECT 2274.5400 1914.5400 2276.1400 1915.0200 ;
        RECT 2274.5400 1919.9800 2276.1400 1920.4600 ;
        RECT 2274.5400 1925.4200 2276.1400 1925.9000 ;
        RECT 2274.5400 1903.6600 2276.1400 1904.1400 ;
        RECT 2274.5400 1909.1000 2276.1400 1909.5800 ;
        RECT 2229.5400 1914.5400 2231.1400 1915.0200 ;
        RECT 2229.5400 1919.9800 2231.1400 1920.4600 ;
        RECT 2229.5400 1925.4200 2231.1400 1925.9000 ;
        RECT 2229.5400 1903.6600 2231.1400 1904.1400 ;
        RECT 2229.5400 1909.1000 2231.1400 1909.5800 ;
        RECT 2184.5400 1941.7400 2186.1400 1942.2200 ;
        RECT 2184.5400 1947.1800 2186.1400 1947.6600 ;
        RECT 2184.5400 1952.6200 2186.1400 1953.1000 ;
        RECT 2176.7800 1941.7400 2178.3800 1942.2200 ;
        RECT 2176.7800 1947.1800 2178.3800 1947.6600 ;
        RECT 2176.7800 1952.6200 2178.3800 1953.1000 ;
        RECT 2184.5400 1930.8600 2186.1400 1931.3400 ;
        RECT 2184.5400 1936.3000 2186.1400 1936.7800 ;
        RECT 2176.7800 1930.8600 2178.3800 1931.3400 ;
        RECT 2176.7800 1936.3000 2178.3800 1936.7800 ;
        RECT 2184.5400 1914.5400 2186.1400 1915.0200 ;
        RECT 2184.5400 1919.9800 2186.1400 1920.4600 ;
        RECT 2184.5400 1925.4200 2186.1400 1925.9000 ;
        RECT 2176.7800 1914.5400 2178.3800 1915.0200 ;
        RECT 2176.7800 1919.9800 2178.3800 1920.4600 ;
        RECT 2176.7800 1925.4200 2178.3800 1925.9000 ;
        RECT 2184.5400 1903.6600 2186.1400 1904.1400 ;
        RECT 2184.5400 1909.1000 2186.1400 1909.5800 ;
        RECT 2176.7800 1903.6600 2178.3800 1904.1400 ;
        RECT 2176.7800 1909.1000 2178.3800 1909.5800 ;
        RECT 2374.2800 1887.3400 2375.8800 1887.8200 ;
        RECT 2374.2800 1892.7800 2375.8800 1893.2600 ;
        RECT 2374.2800 1898.2200 2375.8800 1898.7000 ;
        RECT 2364.5400 1887.3400 2366.1400 1887.8200 ;
        RECT 2364.5400 1892.7800 2366.1400 1893.2600 ;
        RECT 2364.5400 1898.2200 2366.1400 1898.7000 ;
        RECT 2374.2800 1876.4600 2375.8800 1876.9400 ;
        RECT 2374.2800 1881.9000 2375.8800 1882.3800 ;
        RECT 2364.5400 1876.4600 2366.1400 1876.9400 ;
        RECT 2364.5400 1881.9000 2366.1400 1882.3800 ;
        RECT 2374.2800 1860.1400 2375.8800 1860.6200 ;
        RECT 2374.2800 1865.5800 2375.8800 1866.0600 ;
        RECT 2374.2800 1871.0200 2375.8800 1871.5000 ;
        RECT 2364.5400 1860.1400 2366.1400 1860.6200 ;
        RECT 2364.5400 1865.5800 2366.1400 1866.0600 ;
        RECT 2364.5400 1871.0200 2366.1400 1871.5000 ;
        RECT 2374.2800 1849.2600 2375.8800 1849.7400 ;
        RECT 2374.2800 1854.7000 2375.8800 1855.1800 ;
        RECT 2364.5400 1849.2600 2366.1400 1849.7400 ;
        RECT 2364.5400 1854.7000 2366.1400 1855.1800 ;
        RECT 2319.5400 1887.3400 2321.1400 1887.8200 ;
        RECT 2319.5400 1892.7800 2321.1400 1893.2600 ;
        RECT 2319.5400 1898.2200 2321.1400 1898.7000 ;
        RECT 2319.5400 1876.4600 2321.1400 1876.9400 ;
        RECT 2319.5400 1881.9000 2321.1400 1882.3800 ;
        RECT 2319.5400 1860.1400 2321.1400 1860.6200 ;
        RECT 2319.5400 1865.5800 2321.1400 1866.0600 ;
        RECT 2319.5400 1871.0200 2321.1400 1871.5000 ;
        RECT 2319.5400 1849.2600 2321.1400 1849.7400 ;
        RECT 2319.5400 1854.7000 2321.1400 1855.1800 ;
        RECT 2374.2800 1832.9400 2375.8800 1833.4200 ;
        RECT 2374.2800 1838.3800 2375.8800 1838.8600 ;
        RECT 2374.2800 1843.8200 2375.8800 1844.3000 ;
        RECT 2364.5400 1832.9400 2366.1400 1833.4200 ;
        RECT 2364.5400 1838.3800 2366.1400 1838.8600 ;
        RECT 2364.5400 1843.8200 2366.1400 1844.3000 ;
        RECT 2374.2800 1822.0600 2375.8800 1822.5400 ;
        RECT 2374.2800 1827.5000 2375.8800 1827.9800 ;
        RECT 2364.5400 1822.0600 2366.1400 1822.5400 ;
        RECT 2364.5400 1827.5000 2366.1400 1827.9800 ;
        RECT 2374.2800 1805.7400 2375.8800 1806.2200 ;
        RECT 2374.2800 1811.1800 2375.8800 1811.6600 ;
        RECT 2374.2800 1816.6200 2375.8800 1817.1000 ;
        RECT 2364.5400 1805.7400 2366.1400 1806.2200 ;
        RECT 2364.5400 1811.1800 2366.1400 1811.6600 ;
        RECT 2364.5400 1816.6200 2366.1400 1817.1000 ;
        RECT 2364.5400 1800.3000 2366.1400 1800.7800 ;
        RECT 2374.2800 1800.3000 2375.8800 1800.7800 ;
        RECT 2319.5400 1832.9400 2321.1400 1833.4200 ;
        RECT 2319.5400 1838.3800 2321.1400 1838.8600 ;
        RECT 2319.5400 1843.8200 2321.1400 1844.3000 ;
        RECT 2319.5400 1822.0600 2321.1400 1822.5400 ;
        RECT 2319.5400 1827.5000 2321.1400 1827.9800 ;
        RECT 2319.5400 1805.7400 2321.1400 1806.2200 ;
        RECT 2319.5400 1811.1800 2321.1400 1811.6600 ;
        RECT 2319.5400 1816.6200 2321.1400 1817.1000 ;
        RECT 2319.5400 1800.3000 2321.1400 1800.7800 ;
        RECT 2274.5400 1887.3400 2276.1400 1887.8200 ;
        RECT 2274.5400 1892.7800 2276.1400 1893.2600 ;
        RECT 2274.5400 1898.2200 2276.1400 1898.7000 ;
        RECT 2274.5400 1876.4600 2276.1400 1876.9400 ;
        RECT 2274.5400 1881.9000 2276.1400 1882.3800 ;
        RECT 2229.5400 1887.3400 2231.1400 1887.8200 ;
        RECT 2229.5400 1892.7800 2231.1400 1893.2600 ;
        RECT 2229.5400 1898.2200 2231.1400 1898.7000 ;
        RECT 2229.5400 1876.4600 2231.1400 1876.9400 ;
        RECT 2229.5400 1881.9000 2231.1400 1882.3800 ;
        RECT 2274.5400 1860.1400 2276.1400 1860.6200 ;
        RECT 2274.5400 1865.5800 2276.1400 1866.0600 ;
        RECT 2274.5400 1871.0200 2276.1400 1871.5000 ;
        RECT 2274.5400 1849.2600 2276.1400 1849.7400 ;
        RECT 2274.5400 1854.7000 2276.1400 1855.1800 ;
        RECT 2229.5400 1860.1400 2231.1400 1860.6200 ;
        RECT 2229.5400 1865.5800 2231.1400 1866.0600 ;
        RECT 2229.5400 1871.0200 2231.1400 1871.5000 ;
        RECT 2229.5400 1849.2600 2231.1400 1849.7400 ;
        RECT 2229.5400 1854.7000 2231.1400 1855.1800 ;
        RECT 2184.5400 1887.3400 2186.1400 1887.8200 ;
        RECT 2184.5400 1892.7800 2186.1400 1893.2600 ;
        RECT 2184.5400 1898.2200 2186.1400 1898.7000 ;
        RECT 2176.7800 1887.3400 2178.3800 1887.8200 ;
        RECT 2176.7800 1892.7800 2178.3800 1893.2600 ;
        RECT 2176.7800 1898.2200 2178.3800 1898.7000 ;
        RECT 2184.5400 1876.4600 2186.1400 1876.9400 ;
        RECT 2184.5400 1881.9000 2186.1400 1882.3800 ;
        RECT 2176.7800 1876.4600 2178.3800 1876.9400 ;
        RECT 2176.7800 1881.9000 2178.3800 1882.3800 ;
        RECT 2184.5400 1860.1400 2186.1400 1860.6200 ;
        RECT 2184.5400 1865.5800 2186.1400 1866.0600 ;
        RECT 2184.5400 1871.0200 2186.1400 1871.5000 ;
        RECT 2176.7800 1860.1400 2178.3800 1860.6200 ;
        RECT 2176.7800 1865.5800 2178.3800 1866.0600 ;
        RECT 2176.7800 1871.0200 2178.3800 1871.5000 ;
        RECT 2184.5400 1849.2600 2186.1400 1849.7400 ;
        RECT 2184.5400 1854.7000 2186.1400 1855.1800 ;
        RECT 2176.7800 1849.2600 2178.3800 1849.7400 ;
        RECT 2176.7800 1854.7000 2178.3800 1855.1800 ;
        RECT 2274.5400 1832.9400 2276.1400 1833.4200 ;
        RECT 2274.5400 1838.3800 2276.1400 1838.8600 ;
        RECT 2274.5400 1843.8200 2276.1400 1844.3000 ;
        RECT 2274.5400 1822.0600 2276.1400 1822.5400 ;
        RECT 2274.5400 1827.5000 2276.1400 1827.9800 ;
        RECT 2229.5400 1832.9400 2231.1400 1833.4200 ;
        RECT 2229.5400 1838.3800 2231.1400 1838.8600 ;
        RECT 2229.5400 1843.8200 2231.1400 1844.3000 ;
        RECT 2229.5400 1822.0600 2231.1400 1822.5400 ;
        RECT 2229.5400 1827.5000 2231.1400 1827.9800 ;
        RECT 2274.5400 1805.7400 2276.1400 1806.2200 ;
        RECT 2274.5400 1811.1800 2276.1400 1811.6600 ;
        RECT 2274.5400 1816.6200 2276.1400 1817.1000 ;
        RECT 2274.5400 1800.3000 2276.1400 1800.7800 ;
        RECT 2229.5400 1805.7400 2231.1400 1806.2200 ;
        RECT 2229.5400 1811.1800 2231.1400 1811.6600 ;
        RECT 2229.5400 1816.6200 2231.1400 1817.1000 ;
        RECT 2229.5400 1800.3000 2231.1400 1800.7800 ;
        RECT 2184.5400 1832.9400 2186.1400 1833.4200 ;
        RECT 2184.5400 1838.3800 2186.1400 1838.8600 ;
        RECT 2184.5400 1843.8200 2186.1400 1844.3000 ;
        RECT 2176.7800 1832.9400 2178.3800 1833.4200 ;
        RECT 2176.7800 1838.3800 2178.3800 1838.8600 ;
        RECT 2176.7800 1843.8200 2178.3800 1844.3000 ;
        RECT 2184.5400 1822.0600 2186.1400 1822.5400 ;
        RECT 2184.5400 1827.5000 2186.1400 1827.9800 ;
        RECT 2176.7800 1822.0600 2178.3800 1822.5400 ;
        RECT 2176.7800 1827.5000 2178.3800 1827.9800 ;
        RECT 2184.5400 1805.7400 2186.1400 1806.2200 ;
        RECT 2184.5400 1811.1800 2186.1400 1811.6600 ;
        RECT 2184.5400 1816.6200 2186.1400 1817.1000 ;
        RECT 2176.7800 1805.7400 2178.3800 1806.2200 ;
        RECT 2176.7800 1811.1800 2178.3800 1811.6600 ;
        RECT 2176.7800 1816.6200 2178.3800 1817.1000 ;
        RECT 2176.7800 1800.3000 2178.3800 1800.7800 ;
        RECT 2184.5400 1800.3000 2186.1400 1800.7800 ;
        RECT 2171.2200 2002.6100 2381.4400 2004.2100 ;
        RECT 2171.2200 1796.1100 2381.4400 1797.7100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1790.6800 2178.3800 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 2008.7200 2178.3800 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1790.6800 2375.8800 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 2008.7200 2375.8800 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1796.1100 2172.8200 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1796.1100 2381.4400 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 2002.6100 2172.8200 2004.2100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 2002.6100 2381.4400 2004.2100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 1566.4700 2366.1400 1774.5700 ;
        RECT 2319.5400 1566.4700 2321.1400 1774.5700 ;
        RECT 2274.5400 1566.4700 2276.1400 1774.5700 ;
        RECT 2229.5400 1566.4700 2231.1400 1774.5700 ;
        RECT 2184.5400 1566.4700 2186.1400 1774.5700 ;
        RECT 2374.2800 1561.0400 2375.8800 1780.6800 ;
        RECT 2176.7800 1561.0400 2178.3800 1780.6800 ;
      LAYER met3 ;
        RECT 2374.2800 1755.6200 2375.8800 1756.1000 ;
        RECT 2374.2800 1761.0600 2375.8800 1761.5400 ;
        RECT 2364.5400 1755.6200 2366.1400 1756.1000 ;
        RECT 2364.5400 1761.0600 2366.1400 1761.5400 ;
        RECT 2364.5400 1766.5000 2366.1400 1766.9800 ;
        RECT 2374.2800 1766.5000 2375.8800 1766.9800 ;
        RECT 2374.2800 1744.7400 2375.8800 1745.2200 ;
        RECT 2374.2800 1750.1800 2375.8800 1750.6600 ;
        RECT 2364.5400 1744.7400 2366.1400 1745.2200 ;
        RECT 2364.5400 1750.1800 2366.1400 1750.6600 ;
        RECT 2374.2800 1728.4200 2375.8800 1728.9000 ;
        RECT 2374.2800 1733.8600 2375.8800 1734.3400 ;
        RECT 2364.5400 1728.4200 2366.1400 1728.9000 ;
        RECT 2364.5400 1733.8600 2366.1400 1734.3400 ;
        RECT 2364.5400 1739.3000 2366.1400 1739.7800 ;
        RECT 2374.2800 1739.3000 2375.8800 1739.7800 ;
        RECT 2319.5400 1755.6200 2321.1400 1756.1000 ;
        RECT 2319.5400 1761.0600 2321.1400 1761.5400 ;
        RECT 2319.5400 1766.5000 2321.1400 1766.9800 ;
        RECT 2319.5400 1744.7400 2321.1400 1745.2200 ;
        RECT 2319.5400 1750.1800 2321.1400 1750.6600 ;
        RECT 2319.5400 1728.4200 2321.1400 1728.9000 ;
        RECT 2319.5400 1733.8600 2321.1400 1734.3400 ;
        RECT 2319.5400 1739.3000 2321.1400 1739.7800 ;
        RECT 2374.2800 1712.1000 2375.8800 1712.5800 ;
        RECT 2374.2800 1717.5400 2375.8800 1718.0200 ;
        RECT 2374.2800 1722.9800 2375.8800 1723.4600 ;
        RECT 2364.5400 1712.1000 2366.1400 1712.5800 ;
        RECT 2364.5400 1717.5400 2366.1400 1718.0200 ;
        RECT 2364.5400 1722.9800 2366.1400 1723.4600 ;
        RECT 2374.2800 1701.2200 2375.8800 1701.7000 ;
        RECT 2374.2800 1706.6600 2375.8800 1707.1400 ;
        RECT 2364.5400 1701.2200 2366.1400 1701.7000 ;
        RECT 2364.5400 1706.6600 2366.1400 1707.1400 ;
        RECT 2374.2800 1684.9000 2375.8800 1685.3800 ;
        RECT 2374.2800 1690.3400 2375.8800 1690.8200 ;
        RECT 2374.2800 1695.7800 2375.8800 1696.2600 ;
        RECT 2364.5400 1684.9000 2366.1400 1685.3800 ;
        RECT 2364.5400 1690.3400 2366.1400 1690.8200 ;
        RECT 2364.5400 1695.7800 2366.1400 1696.2600 ;
        RECT 2374.2800 1674.0200 2375.8800 1674.5000 ;
        RECT 2374.2800 1679.4600 2375.8800 1679.9400 ;
        RECT 2364.5400 1674.0200 2366.1400 1674.5000 ;
        RECT 2364.5400 1679.4600 2366.1400 1679.9400 ;
        RECT 2319.5400 1712.1000 2321.1400 1712.5800 ;
        RECT 2319.5400 1717.5400 2321.1400 1718.0200 ;
        RECT 2319.5400 1722.9800 2321.1400 1723.4600 ;
        RECT 2319.5400 1701.2200 2321.1400 1701.7000 ;
        RECT 2319.5400 1706.6600 2321.1400 1707.1400 ;
        RECT 2319.5400 1684.9000 2321.1400 1685.3800 ;
        RECT 2319.5400 1690.3400 2321.1400 1690.8200 ;
        RECT 2319.5400 1695.7800 2321.1400 1696.2600 ;
        RECT 2319.5400 1674.0200 2321.1400 1674.5000 ;
        RECT 2319.5400 1679.4600 2321.1400 1679.9400 ;
        RECT 2274.5400 1755.6200 2276.1400 1756.1000 ;
        RECT 2274.5400 1761.0600 2276.1400 1761.5400 ;
        RECT 2274.5400 1766.5000 2276.1400 1766.9800 ;
        RECT 2229.5400 1755.6200 2231.1400 1756.1000 ;
        RECT 2229.5400 1761.0600 2231.1400 1761.5400 ;
        RECT 2229.5400 1766.5000 2231.1400 1766.9800 ;
        RECT 2274.5400 1744.7400 2276.1400 1745.2200 ;
        RECT 2274.5400 1750.1800 2276.1400 1750.6600 ;
        RECT 2274.5400 1728.4200 2276.1400 1728.9000 ;
        RECT 2274.5400 1733.8600 2276.1400 1734.3400 ;
        RECT 2274.5400 1739.3000 2276.1400 1739.7800 ;
        RECT 2229.5400 1744.7400 2231.1400 1745.2200 ;
        RECT 2229.5400 1750.1800 2231.1400 1750.6600 ;
        RECT 2229.5400 1728.4200 2231.1400 1728.9000 ;
        RECT 2229.5400 1733.8600 2231.1400 1734.3400 ;
        RECT 2229.5400 1739.3000 2231.1400 1739.7800 ;
        RECT 2184.5400 1755.6200 2186.1400 1756.1000 ;
        RECT 2184.5400 1761.0600 2186.1400 1761.5400 ;
        RECT 2176.7800 1755.6200 2178.3800 1756.1000 ;
        RECT 2176.7800 1761.0600 2178.3800 1761.5400 ;
        RECT 2176.7800 1766.5000 2178.3800 1766.9800 ;
        RECT 2184.5400 1766.5000 2186.1400 1766.9800 ;
        RECT 2184.5400 1744.7400 2186.1400 1745.2200 ;
        RECT 2184.5400 1750.1800 2186.1400 1750.6600 ;
        RECT 2176.7800 1744.7400 2178.3800 1745.2200 ;
        RECT 2176.7800 1750.1800 2178.3800 1750.6600 ;
        RECT 2184.5400 1728.4200 2186.1400 1728.9000 ;
        RECT 2184.5400 1733.8600 2186.1400 1734.3400 ;
        RECT 2176.7800 1728.4200 2178.3800 1728.9000 ;
        RECT 2176.7800 1733.8600 2178.3800 1734.3400 ;
        RECT 2176.7800 1739.3000 2178.3800 1739.7800 ;
        RECT 2184.5400 1739.3000 2186.1400 1739.7800 ;
        RECT 2274.5400 1712.1000 2276.1400 1712.5800 ;
        RECT 2274.5400 1717.5400 2276.1400 1718.0200 ;
        RECT 2274.5400 1722.9800 2276.1400 1723.4600 ;
        RECT 2274.5400 1701.2200 2276.1400 1701.7000 ;
        RECT 2274.5400 1706.6600 2276.1400 1707.1400 ;
        RECT 2229.5400 1712.1000 2231.1400 1712.5800 ;
        RECT 2229.5400 1717.5400 2231.1400 1718.0200 ;
        RECT 2229.5400 1722.9800 2231.1400 1723.4600 ;
        RECT 2229.5400 1701.2200 2231.1400 1701.7000 ;
        RECT 2229.5400 1706.6600 2231.1400 1707.1400 ;
        RECT 2274.5400 1684.9000 2276.1400 1685.3800 ;
        RECT 2274.5400 1690.3400 2276.1400 1690.8200 ;
        RECT 2274.5400 1695.7800 2276.1400 1696.2600 ;
        RECT 2274.5400 1674.0200 2276.1400 1674.5000 ;
        RECT 2274.5400 1679.4600 2276.1400 1679.9400 ;
        RECT 2229.5400 1684.9000 2231.1400 1685.3800 ;
        RECT 2229.5400 1690.3400 2231.1400 1690.8200 ;
        RECT 2229.5400 1695.7800 2231.1400 1696.2600 ;
        RECT 2229.5400 1674.0200 2231.1400 1674.5000 ;
        RECT 2229.5400 1679.4600 2231.1400 1679.9400 ;
        RECT 2184.5400 1712.1000 2186.1400 1712.5800 ;
        RECT 2184.5400 1717.5400 2186.1400 1718.0200 ;
        RECT 2184.5400 1722.9800 2186.1400 1723.4600 ;
        RECT 2176.7800 1712.1000 2178.3800 1712.5800 ;
        RECT 2176.7800 1717.5400 2178.3800 1718.0200 ;
        RECT 2176.7800 1722.9800 2178.3800 1723.4600 ;
        RECT 2184.5400 1701.2200 2186.1400 1701.7000 ;
        RECT 2184.5400 1706.6600 2186.1400 1707.1400 ;
        RECT 2176.7800 1701.2200 2178.3800 1701.7000 ;
        RECT 2176.7800 1706.6600 2178.3800 1707.1400 ;
        RECT 2184.5400 1684.9000 2186.1400 1685.3800 ;
        RECT 2184.5400 1690.3400 2186.1400 1690.8200 ;
        RECT 2184.5400 1695.7800 2186.1400 1696.2600 ;
        RECT 2176.7800 1684.9000 2178.3800 1685.3800 ;
        RECT 2176.7800 1690.3400 2178.3800 1690.8200 ;
        RECT 2176.7800 1695.7800 2178.3800 1696.2600 ;
        RECT 2184.5400 1674.0200 2186.1400 1674.5000 ;
        RECT 2184.5400 1679.4600 2186.1400 1679.9400 ;
        RECT 2176.7800 1674.0200 2178.3800 1674.5000 ;
        RECT 2176.7800 1679.4600 2178.3800 1679.9400 ;
        RECT 2374.2800 1657.7000 2375.8800 1658.1800 ;
        RECT 2374.2800 1663.1400 2375.8800 1663.6200 ;
        RECT 2374.2800 1668.5800 2375.8800 1669.0600 ;
        RECT 2364.5400 1657.7000 2366.1400 1658.1800 ;
        RECT 2364.5400 1663.1400 2366.1400 1663.6200 ;
        RECT 2364.5400 1668.5800 2366.1400 1669.0600 ;
        RECT 2374.2800 1646.8200 2375.8800 1647.3000 ;
        RECT 2374.2800 1652.2600 2375.8800 1652.7400 ;
        RECT 2364.5400 1646.8200 2366.1400 1647.3000 ;
        RECT 2364.5400 1652.2600 2366.1400 1652.7400 ;
        RECT 2374.2800 1630.5000 2375.8800 1630.9800 ;
        RECT 2374.2800 1635.9400 2375.8800 1636.4200 ;
        RECT 2374.2800 1641.3800 2375.8800 1641.8600 ;
        RECT 2364.5400 1630.5000 2366.1400 1630.9800 ;
        RECT 2364.5400 1635.9400 2366.1400 1636.4200 ;
        RECT 2364.5400 1641.3800 2366.1400 1641.8600 ;
        RECT 2374.2800 1619.6200 2375.8800 1620.1000 ;
        RECT 2374.2800 1625.0600 2375.8800 1625.5400 ;
        RECT 2364.5400 1619.6200 2366.1400 1620.1000 ;
        RECT 2364.5400 1625.0600 2366.1400 1625.5400 ;
        RECT 2319.5400 1657.7000 2321.1400 1658.1800 ;
        RECT 2319.5400 1663.1400 2321.1400 1663.6200 ;
        RECT 2319.5400 1668.5800 2321.1400 1669.0600 ;
        RECT 2319.5400 1646.8200 2321.1400 1647.3000 ;
        RECT 2319.5400 1652.2600 2321.1400 1652.7400 ;
        RECT 2319.5400 1630.5000 2321.1400 1630.9800 ;
        RECT 2319.5400 1635.9400 2321.1400 1636.4200 ;
        RECT 2319.5400 1641.3800 2321.1400 1641.8600 ;
        RECT 2319.5400 1619.6200 2321.1400 1620.1000 ;
        RECT 2319.5400 1625.0600 2321.1400 1625.5400 ;
        RECT 2374.2800 1603.3000 2375.8800 1603.7800 ;
        RECT 2374.2800 1608.7400 2375.8800 1609.2200 ;
        RECT 2374.2800 1614.1800 2375.8800 1614.6600 ;
        RECT 2364.5400 1603.3000 2366.1400 1603.7800 ;
        RECT 2364.5400 1608.7400 2366.1400 1609.2200 ;
        RECT 2364.5400 1614.1800 2366.1400 1614.6600 ;
        RECT 2374.2800 1592.4200 2375.8800 1592.9000 ;
        RECT 2374.2800 1597.8600 2375.8800 1598.3400 ;
        RECT 2364.5400 1592.4200 2366.1400 1592.9000 ;
        RECT 2364.5400 1597.8600 2366.1400 1598.3400 ;
        RECT 2374.2800 1576.1000 2375.8800 1576.5800 ;
        RECT 2374.2800 1581.5400 2375.8800 1582.0200 ;
        RECT 2374.2800 1586.9800 2375.8800 1587.4600 ;
        RECT 2364.5400 1576.1000 2366.1400 1576.5800 ;
        RECT 2364.5400 1581.5400 2366.1400 1582.0200 ;
        RECT 2364.5400 1586.9800 2366.1400 1587.4600 ;
        RECT 2364.5400 1570.6600 2366.1400 1571.1400 ;
        RECT 2374.2800 1570.6600 2375.8800 1571.1400 ;
        RECT 2319.5400 1603.3000 2321.1400 1603.7800 ;
        RECT 2319.5400 1608.7400 2321.1400 1609.2200 ;
        RECT 2319.5400 1614.1800 2321.1400 1614.6600 ;
        RECT 2319.5400 1592.4200 2321.1400 1592.9000 ;
        RECT 2319.5400 1597.8600 2321.1400 1598.3400 ;
        RECT 2319.5400 1576.1000 2321.1400 1576.5800 ;
        RECT 2319.5400 1581.5400 2321.1400 1582.0200 ;
        RECT 2319.5400 1586.9800 2321.1400 1587.4600 ;
        RECT 2319.5400 1570.6600 2321.1400 1571.1400 ;
        RECT 2274.5400 1657.7000 2276.1400 1658.1800 ;
        RECT 2274.5400 1663.1400 2276.1400 1663.6200 ;
        RECT 2274.5400 1668.5800 2276.1400 1669.0600 ;
        RECT 2274.5400 1646.8200 2276.1400 1647.3000 ;
        RECT 2274.5400 1652.2600 2276.1400 1652.7400 ;
        RECT 2229.5400 1657.7000 2231.1400 1658.1800 ;
        RECT 2229.5400 1663.1400 2231.1400 1663.6200 ;
        RECT 2229.5400 1668.5800 2231.1400 1669.0600 ;
        RECT 2229.5400 1646.8200 2231.1400 1647.3000 ;
        RECT 2229.5400 1652.2600 2231.1400 1652.7400 ;
        RECT 2274.5400 1630.5000 2276.1400 1630.9800 ;
        RECT 2274.5400 1635.9400 2276.1400 1636.4200 ;
        RECT 2274.5400 1641.3800 2276.1400 1641.8600 ;
        RECT 2274.5400 1619.6200 2276.1400 1620.1000 ;
        RECT 2274.5400 1625.0600 2276.1400 1625.5400 ;
        RECT 2229.5400 1630.5000 2231.1400 1630.9800 ;
        RECT 2229.5400 1635.9400 2231.1400 1636.4200 ;
        RECT 2229.5400 1641.3800 2231.1400 1641.8600 ;
        RECT 2229.5400 1619.6200 2231.1400 1620.1000 ;
        RECT 2229.5400 1625.0600 2231.1400 1625.5400 ;
        RECT 2184.5400 1657.7000 2186.1400 1658.1800 ;
        RECT 2184.5400 1663.1400 2186.1400 1663.6200 ;
        RECT 2184.5400 1668.5800 2186.1400 1669.0600 ;
        RECT 2176.7800 1657.7000 2178.3800 1658.1800 ;
        RECT 2176.7800 1663.1400 2178.3800 1663.6200 ;
        RECT 2176.7800 1668.5800 2178.3800 1669.0600 ;
        RECT 2184.5400 1646.8200 2186.1400 1647.3000 ;
        RECT 2184.5400 1652.2600 2186.1400 1652.7400 ;
        RECT 2176.7800 1646.8200 2178.3800 1647.3000 ;
        RECT 2176.7800 1652.2600 2178.3800 1652.7400 ;
        RECT 2184.5400 1630.5000 2186.1400 1630.9800 ;
        RECT 2184.5400 1635.9400 2186.1400 1636.4200 ;
        RECT 2184.5400 1641.3800 2186.1400 1641.8600 ;
        RECT 2176.7800 1630.5000 2178.3800 1630.9800 ;
        RECT 2176.7800 1635.9400 2178.3800 1636.4200 ;
        RECT 2176.7800 1641.3800 2178.3800 1641.8600 ;
        RECT 2184.5400 1619.6200 2186.1400 1620.1000 ;
        RECT 2184.5400 1625.0600 2186.1400 1625.5400 ;
        RECT 2176.7800 1619.6200 2178.3800 1620.1000 ;
        RECT 2176.7800 1625.0600 2178.3800 1625.5400 ;
        RECT 2274.5400 1603.3000 2276.1400 1603.7800 ;
        RECT 2274.5400 1608.7400 2276.1400 1609.2200 ;
        RECT 2274.5400 1614.1800 2276.1400 1614.6600 ;
        RECT 2274.5400 1592.4200 2276.1400 1592.9000 ;
        RECT 2274.5400 1597.8600 2276.1400 1598.3400 ;
        RECT 2229.5400 1603.3000 2231.1400 1603.7800 ;
        RECT 2229.5400 1608.7400 2231.1400 1609.2200 ;
        RECT 2229.5400 1614.1800 2231.1400 1614.6600 ;
        RECT 2229.5400 1592.4200 2231.1400 1592.9000 ;
        RECT 2229.5400 1597.8600 2231.1400 1598.3400 ;
        RECT 2274.5400 1576.1000 2276.1400 1576.5800 ;
        RECT 2274.5400 1581.5400 2276.1400 1582.0200 ;
        RECT 2274.5400 1586.9800 2276.1400 1587.4600 ;
        RECT 2274.5400 1570.6600 2276.1400 1571.1400 ;
        RECT 2229.5400 1576.1000 2231.1400 1576.5800 ;
        RECT 2229.5400 1581.5400 2231.1400 1582.0200 ;
        RECT 2229.5400 1586.9800 2231.1400 1587.4600 ;
        RECT 2229.5400 1570.6600 2231.1400 1571.1400 ;
        RECT 2184.5400 1603.3000 2186.1400 1603.7800 ;
        RECT 2184.5400 1608.7400 2186.1400 1609.2200 ;
        RECT 2184.5400 1614.1800 2186.1400 1614.6600 ;
        RECT 2176.7800 1603.3000 2178.3800 1603.7800 ;
        RECT 2176.7800 1608.7400 2178.3800 1609.2200 ;
        RECT 2176.7800 1614.1800 2178.3800 1614.6600 ;
        RECT 2184.5400 1592.4200 2186.1400 1592.9000 ;
        RECT 2184.5400 1597.8600 2186.1400 1598.3400 ;
        RECT 2176.7800 1592.4200 2178.3800 1592.9000 ;
        RECT 2176.7800 1597.8600 2178.3800 1598.3400 ;
        RECT 2184.5400 1576.1000 2186.1400 1576.5800 ;
        RECT 2184.5400 1581.5400 2186.1400 1582.0200 ;
        RECT 2184.5400 1586.9800 2186.1400 1587.4600 ;
        RECT 2176.7800 1576.1000 2178.3800 1576.5800 ;
        RECT 2176.7800 1581.5400 2178.3800 1582.0200 ;
        RECT 2176.7800 1586.9800 2178.3800 1587.4600 ;
        RECT 2176.7800 1570.6600 2178.3800 1571.1400 ;
        RECT 2184.5400 1570.6600 2186.1400 1571.1400 ;
        RECT 2171.2200 1772.9700 2381.4400 1774.5700 ;
        RECT 2171.2200 1566.4700 2381.4400 1568.0700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1561.0400 2178.3800 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1779.0800 2178.3800 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1561.0400 2375.8800 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1779.0800 2375.8800 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1566.4700 2172.8200 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1566.4700 2381.4400 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1772.9700 2172.8200 1774.5700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1772.9700 2381.4400 1774.5700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 1336.8300 2366.1400 1544.9300 ;
        RECT 2319.5400 1336.8300 2321.1400 1544.9300 ;
        RECT 2274.5400 1336.8300 2276.1400 1544.9300 ;
        RECT 2229.5400 1336.8300 2231.1400 1544.9300 ;
        RECT 2184.5400 1336.8300 2186.1400 1544.9300 ;
        RECT 2374.2800 1331.4000 2375.8800 1551.0400 ;
        RECT 2176.7800 1331.4000 2178.3800 1551.0400 ;
      LAYER met3 ;
        RECT 2374.2800 1525.9800 2375.8800 1526.4600 ;
        RECT 2374.2800 1531.4200 2375.8800 1531.9000 ;
        RECT 2364.5400 1525.9800 2366.1400 1526.4600 ;
        RECT 2364.5400 1531.4200 2366.1400 1531.9000 ;
        RECT 2364.5400 1536.8600 2366.1400 1537.3400 ;
        RECT 2374.2800 1536.8600 2375.8800 1537.3400 ;
        RECT 2374.2800 1515.1000 2375.8800 1515.5800 ;
        RECT 2374.2800 1520.5400 2375.8800 1521.0200 ;
        RECT 2364.5400 1515.1000 2366.1400 1515.5800 ;
        RECT 2364.5400 1520.5400 2366.1400 1521.0200 ;
        RECT 2374.2800 1498.7800 2375.8800 1499.2600 ;
        RECT 2374.2800 1504.2200 2375.8800 1504.7000 ;
        RECT 2364.5400 1498.7800 2366.1400 1499.2600 ;
        RECT 2364.5400 1504.2200 2366.1400 1504.7000 ;
        RECT 2364.5400 1509.6600 2366.1400 1510.1400 ;
        RECT 2374.2800 1509.6600 2375.8800 1510.1400 ;
        RECT 2319.5400 1525.9800 2321.1400 1526.4600 ;
        RECT 2319.5400 1531.4200 2321.1400 1531.9000 ;
        RECT 2319.5400 1536.8600 2321.1400 1537.3400 ;
        RECT 2319.5400 1515.1000 2321.1400 1515.5800 ;
        RECT 2319.5400 1520.5400 2321.1400 1521.0200 ;
        RECT 2319.5400 1498.7800 2321.1400 1499.2600 ;
        RECT 2319.5400 1504.2200 2321.1400 1504.7000 ;
        RECT 2319.5400 1509.6600 2321.1400 1510.1400 ;
        RECT 2374.2800 1482.4600 2375.8800 1482.9400 ;
        RECT 2374.2800 1487.9000 2375.8800 1488.3800 ;
        RECT 2374.2800 1493.3400 2375.8800 1493.8200 ;
        RECT 2364.5400 1482.4600 2366.1400 1482.9400 ;
        RECT 2364.5400 1487.9000 2366.1400 1488.3800 ;
        RECT 2364.5400 1493.3400 2366.1400 1493.8200 ;
        RECT 2374.2800 1471.5800 2375.8800 1472.0600 ;
        RECT 2374.2800 1477.0200 2375.8800 1477.5000 ;
        RECT 2364.5400 1471.5800 2366.1400 1472.0600 ;
        RECT 2364.5400 1477.0200 2366.1400 1477.5000 ;
        RECT 2374.2800 1455.2600 2375.8800 1455.7400 ;
        RECT 2374.2800 1460.7000 2375.8800 1461.1800 ;
        RECT 2374.2800 1466.1400 2375.8800 1466.6200 ;
        RECT 2364.5400 1455.2600 2366.1400 1455.7400 ;
        RECT 2364.5400 1460.7000 2366.1400 1461.1800 ;
        RECT 2364.5400 1466.1400 2366.1400 1466.6200 ;
        RECT 2374.2800 1444.3800 2375.8800 1444.8600 ;
        RECT 2374.2800 1449.8200 2375.8800 1450.3000 ;
        RECT 2364.5400 1444.3800 2366.1400 1444.8600 ;
        RECT 2364.5400 1449.8200 2366.1400 1450.3000 ;
        RECT 2319.5400 1482.4600 2321.1400 1482.9400 ;
        RECT 2319.5400 1487.9000 2321.1400 1488.3800 ;
        RECT 2319.5400 1493.3400 2321.1400 1493.8200 ;
        RECT 2319.5400 1471.5800 2321.1400 1472.0600 ;
        RECT 2319.5400 1477.0200 2321.1400 1477.5000 ;
        RECT 2319.5400 1455.2600 2321.1400 1455.7400 ;
        RECT 2319.5400 1460.7000 2321.1400 1461.1800 ;
        RECT 2319.5400 1466.1400 2321.1400 1466.6200 ;
        RECT 2319.5400 1444.3800 2321.1400 1444.8600 ;
        RECT 2319.5400 1449.8200 2321.1400 1450.3000 ;
        RECT 2274.5400 1525.9800 2276.1400 1526.4600 ;
        RECT 2274.5400 1531.4200 2276.1400 1531.9000 ;
        RECT 2274.5400 1536.8600 2276.1400 1537.3400 ;
        RECT 2229.5400 1525.9800 2231.1400 1526.4600 ;
        RECT 2229.5400 1531.4200 2231.1400 1531.9000 ;
        RECT 2229.5400 1536.8600 2231.1400 1537.3400 ;
        RECT 2274.5400 1515.1000 2276.1400 1515.5800 ;
        RECT 2274.5400 1520.5400 2276.1400 1521.0200 ;
        RECT 2274.5400 1498.7800 2276.1400 1499.2600 ;
        RECT 2274.5400 1504.2200 2276.1400 1504.7000 ;
        RECT 2274.5400 1509.6600 2276.1400 1510.1400 ;
        RECT 2229.5400 1515.1000 2231.1400 1515.5800 ;
        RECT 2229.5400 1520.5400 2231.1400 1521.0200 ;
        RECT 2229.5400 1498.7800 2231.1400 1499.2600 ;
        RECT 2229.5400 1504.2200 2231.1400 1504.7000 ;
        RECT 2229.5400 1509.6600 2231.1400 1510.1400 ;
        RECT 2184.5400 1525.9800 2186.1400 1526.4600 ;
        RECT 2184.5400 1531.4200 2186.1400 1531.9000 ;
        RECT 2176.7800 1525.9800 2178.3800 1526.4600 ;
        RECT 2176.7800 1531.4200 2178.3800 1531.9000 ;
        RECT 2176.7800 1536.8600 2178.3800 1537.3400 ;
        RECT 2184.5400 1536.8600 2186.1400 1537.3400 ;
        RECT 2184.5400 1515.1000 2186.1400 1515.5800 ;
        RECT 2184.5400 1520.5400 2186.1400 1521.0200 ;
        RECT 2176.7800 1515.1000 2178.3800 1515.5800 ;
        RECT 2176.7800 1520.5400 2178.3800 1521.0200 ;
        RECT 2184.5400 1498.7800 2186.1400 1499.2600 ;
        RECT 2184.5400 1504.2200 2186.1400 1504.7000 ;
        RECT 2176.7800 1498.7800 2178.3800 1499.2600 ;
        RECT 2176.7800 1504.2200 2178.3800 1504.7000 ;
        RECT 2176.7800 1509.6600 2178.3800 1510.1400 ;
        RECT 2184.5400 1509.6600 2186.1400 1510.1400 ;
        RECT 2274.5400 1482.4600 2276.1400 1482.9400 ;
        RECT 2274.5400 1487.9000 2276.1400 1488.3800 ;
        RECT 2274.5400 1493.3400 2276.1400 1493.8200 ;
        RECT 2274.5400 1471.5800 2276.1400 1472.0600 ;
        RECT 2274.5400 1477.0200 2276.1400 1477.5000 ;
        RECT 2229.5400 1482.4600 2231.1400 1482.9400 ;
        RECT 2229.5400 1487.9000 2231.1400 1488.3800 ;
        RECT 2229.5400 1493.3400 2231.1400 1493.8200 ;
        RECT 2229.5400 1471.5800 2231.1400 1472.0600 ;
        RECT 2229.5400 1477.0200 2231.1400 1477.5000 ;
        RECT 2274.5400 1455.2600 2276.1400 1455.7400 ;
        RECT 2274.5400 1460.7000 2276.1400 1461.1800 ;
        RECT 2274.5400 1466.1400 2276.1400 1466.6200 ;
        RECT 2274.5400 1444.3800 2276.1400 1444.8600 ;
        RECT 2274.5400 1449.8200 2276.1400 1450.3000 ;
        RECT 2229.5400 1455.2600 2231.1400 1455.7400 ;
        RECT 2229.5400 1460.7000 2231.1400 1461.1800 ;
        RECT 2229.5400 1466.1400 2231.1400 1466.6200 ;
        RECT 2229.5400 1444.3800 2231.1400 1444.8600 ;
        RECT 2229.5400 1449.8200 2231.1400 1450.3000 ;
        RECT 2184.5400 1482.4600 2186.1400 1482.9400 ;
        RECT 2184.5400 1487.9000 2186.1400 1488.3800 ;
        RECT 2184.5400 1493.3400 2186.1400 1493.8200 ;
        RECT 2176.7800 1482.4600 2178.3800 1482.9400 ;
        RECT 2176.7800 1487.9000 2178.3800 1488.3800 ;
        RECT 2176.7800 1493.3400 2178.3800 1493.8200 ;
        RECT 2184.5400 1471.5800 2186.1400 1472.0600 ;
        RECT 2184.5400 1477.0200 2186.1400 1477.5000 ;
        RECT 2176.7800 1471.5800 2178.3800 1472.0600 ;
        RECT 2176.7800 1477.0200 2178.3800 1477.5000 ;
        RECT 2184.5400 1455.2600 2186.1400 1455.7400 ;
        RECT 2184.5400 1460.7000 2186.1400 1461.1800 ;
        RECT 2184.5400 1466.1400 2186.1400 1466.6200 ;
        RECT 2176.7800 1455.2600 2178.3800 1455.7400 ;
        RECT 2176.7800 1460.7000 2178.3800 1461.1800 ;
        RECT 2176.7800 1466.1400 2178.3800 1466.6200 ;
        RECT 2184.5400 1444.3800 2186.1400 1444.8600 ;
        RECT 2184.5400 1449.8200 2186.1400 1450.3000 ;
        RECT 2176.7800 1444.3800 2178.3800 1444.8600 ;
        RECT 2176.7800 1449.8200 2178.3800 1450.3000 ;
        RECT 2374.2800 1428.0600 2375.8800 1428.5400 ;
        RECT 2374.2800 1433.5000 2375.8800 1433.9800 ;
        RECT 2374.2800 1438.9400 2375.8800 1439.4200 ;
        RECT 2364.5400 1428.0600 2366.1400 1428.5400 ;
        RECT 2364.5400 1433.5000 2366.1400 1433.9800 ;
        RECT 2364.5400 1438.9400 2366.1400 1439.4200 ;
        RECT 2374.2800 1417.1800 2375.8800 1417.6600 ;
        RECT 2374.2800 1422.6200 2375.8800 1423.1000 ;
        RECT 2364.5400 1417.1800 2366.1400 1417.6600 ;
        RECT 2364.5400 1422.6200 2366.1400 1423.1000 ;
        RECT 2374.2800 1400.8600 2375.8800 1401.3400 ;
        RECT 2374.2800 1406.3000 2375.8800 1406.7800 ;
        RECT 2374.2800 1411.7400 2375.8800 1412.2200 ;
        RECT 2364.5400 1400.8600 2366.1400 1401.3400 ;
        RECT 2364.5400 1406.3000 2366.1400 1406.7800 ;
        RECT 2364.5400 1411.7400 2366.1400 1412.2200 ;
        RECT 2374.2800 1389.9800 2375.8800 1390.4600 ;
        RECT 2374.2800 1395.4200 2375.8800 1395.9000 ;
        RECT 2364.5400 1389.9800 2366.1400 1390.4600 ;
        RECT 2364.5400 1395.4200 2366.1400 1395.9000 ;
        RECT 2319.5400 1428.0600 2321.1400 1428.5400 ;
        RECT 2319.5400 1433.5000 2321.1400 1433.9800 ;
        RECT 2319.5400 1438.9400 2321.1400 1439.4200 ;
        RECT 2319.5400 1417.1800 2321.1400 1417.6600 ;
        RECT 2319.5400 1422.6200 2321.1400 1423.1000 ;
        RECT 2319.5400 1400.8600 2321.1400 1401.3400 ;
        RECT 2319.5400 1406.3000 2321.1400 1406.7800 ;
        RECT 2319.5400 1411.7400 2321.1400 1412.2200 ;
        RECT 2319.5400 1389.9800 2321.1400 1390.4600 ;
        RECT 2319.5400 1395.4200 2321.1400 1395.9000 ;
        RECT 2374.2800 1373.6600 2375.8800 1374.1400 ;
        RECT 2374.2800 1379.1000 2375.8800 1379.5800 ;
        RECT 2374.2800 1384.5400 2375.8800 1385.0200 ;
        RECT 2364.5400 1373.6600 2366.1400 1374.1400 ;
        RECT 2364.5400 1379.1000 2366.1400 1379.5800 ;
        RECT 2364.5400 1384.5400 2366.1400 1385.0200 ;
        RECT 2374.2800 1362.7800 2375.8800 1363.2600 ;
        RECT 2374.2800 1368.2200 2375.8800 1368.7000 ;
        RECT 2364.5400 1362.7800 2366.1400 1363.2600 ;
        RECT 2364.5400 1368.2200 2366.1400 1368.7000 ;
        RECT 2374.2800 1346.4600 2375.8800 1346.9400 ;
        RECT 2374.2800 1351.9000 2375.8800 1352.3800 ;
        RECT 2374.2800 1357.3400 2375.8800 1357.8200 ;
        RECT 2364.5400 1346.4600 2366.1400 1346.9400 ;
        RECT 2364.5400 1351.9000 2366.1400 1352.3800 ;
        RECT 2364.5400 1357.3400 2366.1400 1357.8200 ;
        RECT 2364.5400 1341.0200 2366.1400 1341.5000 ;
        RECT 2374.2800 1341.0200 2375.8800 1341.5000 ;
        RECT 2319.5400 1373.6600 2321.1400 1374.1400 ;
        RECT 2319.5400 1379.1000 2321.1400 1379.5800 ;
        RECT 2319.5400 1384.5400 2321.1400 1385.0200 ;
        RECT 2319.5400 1362.7800 2321.1400 1363.2600 ;
        RECT 2319.5400 1368.2200 2321.1400 1368.7000 ;
        RECT 2319.5400 1346.4600 2321.1400 1346.9400 ;
        RECT 2319.5400 1351.9000 2321.1400 1352.3800 ;
        RECT 2319.5400 1357.3400 2321.1400 1357.8200 ;
        RECT 2319.5400 1341.0200 2321.1400 1341.5000 ;
        RECT 2274.5400 1428.0600 2276.1400 1428.5400 ;
        RECT 2274.5400 1433.5000 2276.1400 1433.9800 ;
        RECT 2274.5400 1438.9400 2276.1400 1439.4200 ;
        RECT 2274.5400 1417.1800 2276.1400 1417.6600 ;
        RECT 2274.5400 1422.6200 2276.1400 1423.1000 ;
        RECT 2229.5400 1428.0600 2231.1400 1428.5400 ;
        RECT 2229.5400 1433.5000 2231.1400 1433.9800 ;
        RECT 2229.5400 1438.9400 2231.1400 1439.4200 ;
        RECT 2229.5400 1417.1800 2231.1400 1417.6600 ;
        RECT 2229.5400 1422.6200 2231.1400 1423.1000 ;
        RECT 2274.5400 1400.8600 2276.1400 1401.3400 ;
        RECT 2274.5400 1406.3000 2276.1400 1406.7800 ;
        RECT 2274.5400 1411.7400 2276.1400 1412.2200 ;
        RECT 2274.5400 1389.9800 2276.1400 1390.4600 ;
        RECT 2274.5400 1395.4200 2276.1400 1395.9000 ;
        RECT 2229.5400 1400.8600 2231.1400 1401.3400 ;
        RECT 2229.5400 1406.3000 2231.1400 1406.7800 ;
        RECT 2229.5400 1411.7400 2231.1400 1412.2200 ;
        RECT 2229.5400 1389.9800 2231.1400 1390.4600 ;
        RECT 2229.5400 1395.4200 2231.1400 1395.9000 ;
        RECT 2184.5400 1428.0600 2186.1400 1428.5400 ;
        RECT 2184.5400 1433.5000 2186.1400 1433.9800 ;
        RECT 2184.5400 1438.9400 2186.1400 1439.4200 ;
        RECT 2176.7800 1428.0600 2178.3800 1428.5400 ;
        RECT 2176.7800 1433.5000 2178.3800 1433.9800 ;
        RECT 2176.7800 1438.9400 2178.3800 1439.4200 ;
        RECT 2184.5400 1417.1800 2186.1400 1417.6600 ;
        RECT 2184.5400 1422.6200 2186.1400 1423.1000 ;
        RECT 2176.7800 1417.1800 2178.3800 1417.6600 ;
        RECT 2176.7800 1422.6200 2178.3800 1423.1000 ;
        RECT 2184.5400 1400.8600 2186.1400 1401.3400 ;
        RECT 2184.5400 1406.3000 2186.1400 1406.7800 ;
        RECT 2184.5400 1411.7400 2186.1400 1412.2200 ;
        RECT 2176.7800 1400.8600 2178.3800 1401.3400 ;
        RECT 2176.7800 1406.3000 2178.3800 1406.7800 ;
        RECT 2176.7800 1411.7400 2178.3800 1412.2200 ;
        RECT 2184.5400 1389.9800 2186.1400 1390.4600 ;
        RECT 2184.5400 1395.4200 2186.1400 1395.9000 ;
        RECT 2176.7800 1389.9800 2178.3800 1390.4600 ;
        RECT 2176.7800 1395.4200 2178.3800 1395.9000 ;
        RECT 2274.5400 1373.6600 2276.1400 1374.1400 ;
        RECT 2274.5400 1379.1000 2276.1400 1379.5800 ;
        RECT 2274.5400 1384.5400 2276.1400 1385.0200 ;
        RECT 2274.5400 1362.7800 2276.1400 1363.2600 ;
        RECT 2274.5400 1368.2200 2276.1400 1368.7000 ;
        RECT 2229.5400 1373.6600 2231.1400 1374.1400 ;
        RECT 2229.5400 1379.1000 2231.1400 1379.5800 ;
        RECT 2229.5400 1384.5400 2231.1400 1385.0200 ;
        RECT 2229.5400 1362.7800 2231.1400 1363.2600 ;
        RECT 2229.5400 1368.2200 2231.1400 1368.7000 ;
        RECT 2274.5400 1346.4600 2276.1400 1346.9400 ;
        RECT 2274.5400 1351.9000 2276.1400 1352.3800 ;
        RECT 2274.5400 1357.3400 2276.1400 1357.8200 ;
        RECT 2274.5400 1341.0200 2276.1400 1341.5000 ;
        RECT 2229.5400 1346.4600 2231.1400 1346.9400 ;
        RECT 2229.5400 1351.9000 2231.1400 1352.3800 ;
        RECT 2229.5400 1357.3400 2231.1400 1357.8200 ;
        RECT 2229.5400 1341.0200 2231.1400 1341.5000 ;
        RECT 2184.5400 1373.6600 2186.1400 1374.1400 ;
        RECT 2184.5400 1379.1000 2186.1400 1379.5800 ;
        RECT 2184.5400 1384.5400 2186.1400 1385.0200 ;
        RECT 2176.7800 1373.6600 2178.3800 1374.1400 ;
        RECT 2176.7800 1379.1000 2178.3800 1379.5800 ;
        RECT 2176.7800 1384.5400 2178.3800 1385.0200 ;
        RECT 2184.5400 1362.7800 2186.1400 1363.2600 ;
        RECT 2184.5400 1368.2200 2186.1400 1368.7000 ;
        RECT 2176.7800 1362.7800 2178.3800 1363.2600 ;
        RECT 2176.7800 1368.2200 2178.3800 1368.7000 ;
        RECT 2184.5400 1346.4600 2186.1400 1346.9400 ;
        RECT 2184.5400 1351.9000 2186.1400 1352.3800 ;
        RECT 2184.5400 1357.3400 2186.1400 1357.8200 ;
        RECT 2176.7800 1346.4600 2178.3800 1346.9400 ;
        RECT 2176.7800 1351.9000 2178.3800 1352.3800 ;
        RECT 2176.7800 1357.3400 2178.3800 1357.8200 ;
        RECT 2176.7800 1341.0200 2178.3800 1341.5000 ;
        RECT 2184.5400 1341.0200 2186.1400 1341.5000 ;
        RECT 2171.2200 1543.3300 2381.4400 1544.9300 ;
        RECT 2171.2200 1336.8300 2381.4400 1338.4300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1331.4000 2178.3800 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1549.4400 2178.3800 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1331.4000 2375.8800 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1549.4400 2375.8800 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1336.8300 2172.8200 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1336.8300 2381.4400 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1543.3300 2172.8200 1544.9300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1543.3300 2381.4400 1544.9300 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 1107.1900 2366.1400 1315.2900 ;
        RECT 2319.5400 1107.1900 2321.1400 1315.2900 ;
        RECT 2274.5400 1107.1900 2276.1400 1315.2900 ;
        RECT 2229.5400 1107.1900 2231.1400 1315.2900 ;
        RECT 2184.5400 1107.1900 2186.1400 1315.2900 ;
        RECT 2374.2800 1101.7600 2375.8800 1321.4000 ;
        RECT 2176.7800 1101.7600 2178.3800 1321.4000 ;
      LAYER met3 ;
        RECT 2374.2800 1296.3400 2375.8800 1296.8200 ;
        RECT 2374.2800 1301.7800 2375.8800 1302.2600 ;
        RECT 2364.5400 1296.3400 2366.1400 1296.8200 ;
        RECT 2364.5400 1301.7800 2366.1400 1302.2600 ;
        RECT 2364.5400 1307.2200 2366.1400 1307.7000 ;
        RECT 2374.2800 1307.2200 2375.8800 1307.7000 ;
        RECT 2374.2800 1285.4600 2375.8800 1285.9400 ;
        RECT 2374.2800 1290.9000 2375.8800 1291.3800 ;
        RECT 2364.5400 1285.4600 2366.1400 1285.9400 ;
        RECT 2364.5400 1290.9000 2366.1400 1291.3800 ;
        RECT 2374.2800 1269.1400 2375.8800 1269.6200 ;
        RECT 2374.2800 1274.5800 2375.8800 1275.0600 ;
        RECT 2364.5400 1269.1400 2366.1400 1269.6200 ;
        RECT 2364.5400 1274.5800 2366.1400 1275.0600 ;
        RECT 2364.5400 1280.0200 2366.1400 1280.5000 ;
        RECT 2374.2800 1280.0200 2375.8800 1280.5000 ;
        RECT 2319.5400 1296.3400 2321.1400 1296.8200 ;
        RECT 2319.5400 1301.7800 2321.1400 1302.2600 ;
        RECT 2319.5400 1307.2200 2321.1400 1307.7000 ;
        RECT 2319.5400 1285.4600 2321.1400 1285.9400 ;
        RECT 2319.5400 1290.9000 2321.1400 1291.3800 ;
        RECT 2319.5400 1269.1400 2321.1400 1269.6200 ;
        RECT 2319.5400 1274.5800 2321.1400 1275.0600 ;
        RECT 2319.5400 1280.0200 2321.1400 1280.5000 ;
        RECT 2374.2800 1252.8200 2375.8800 1253.3000 ;
        RECT 2374.2800 1258.2600 2375.8800 1258.7400 ;
        RECT 2374.2800 1263.7000 2375.8800 1264.1800 ;
        RECT 2364.5400 1252.8200 2366.1400 1253.3000 ;
        RECT 2364.5400 1258.2600 2366.1400 1258.7400 ;
        RECT 2364.5400 1263.7000 2366.1400 1264.1800 ;
        RECT 2374.2800 1241.9400 2375.8800 1242.4200 ;
        RECT 2374.2800 1247.3800 2375.8800 1247.8600 ;
        RECT 2364.5400 1241.9400 2366.1400 1242.4200 ;
        RECT 2364.5400 1247.3800 2366.1400 1247.8600 ;
        RECT 2374.2800 1225.6200 2375.8800 1226.1000 ;
        RECT 2374.2800 1231.0600 2375.8800 1231.5400 ;
        RECT 2374.2800 1236.5000 2375.8800 1236.9800 ;
        RECT 2364.5400 1225.6200 2366.1400 1226.1000 ;
        RECT 2364.5400 1231.0600 2366.1400 1231.5400 ;
        RECT 2364.5400 1236.5000 2366.1400 1236.9800 ;
        RECT 2374.2800 1214.7400 2375.8800 1215.2200 ;
        RECT 2374.2800 1220.1800 2375.8800 1220.6600 ;
        RECT 2364.5400 1214.7400 2366.1400 1215.2200 ;
        RECT 2364.5400 1220.1800 2366.1400 1220.6600 ;
        RECT 2319.5400 1252.8200 2321.1400 1253.3000 ;
        RECT 2319.5400 1258.2600 2321.1400 1258.7400 ;
        RECT 2319.5400 1263.7000 2321.1400 1264.1800 ;
        RECT 2319.5400 1241.9400 2321.1400 1242.4200 ;
        RECT 2319.5400 1247.3800 2321.1400 1247.8600 ;
        RECT 2319.5400 1225.6200 2321.1400 1226.1000 ;
        RECT 2319.5400 1231.0600 2321.1400 1231.5400 ;
        RECT 2319.5400 1236.5000 2321.1400 1236.9800 ;
        RECT 2319.5400 1214.7400 2321.1400 1215.2200 ;
        RECT 2319.5400 1220.1800 2321.1400 1220.6600 ;
        RECT 2274.5400 1296.3400 2276.1400 1296.8200 ;
        RECT 2274.5400 1301.7800 2276.1400 1302.2600 ;
        RECT 2274.5400 1307.2200 2276.1400 1307.7000 ;
        RECT 2229.5400 1296.3400 2231.1400 1296.8200 ;
        RECT 2229.5400 1301.7800 2231.1400 1302.2600 ;
        RECT 2229.5400 1307.2200 2231.1400 1307.7000 ;
        RECT 2274.5400 1285.4600 2276.1400 1285.9400 ;
        RECT 2274.5400 1290.9000 2276.1400 1291.3800 ;
        RECT 2274.5400 1269.1400 2276.1400 1269.6200 ;
        RECT 2274.5400 1274.5800 2276.1400 1275.0600 ;
        RECT 2274.5400 1280.0200 2276.1400 1280.5000 ;
        RECT 2229.5400 1285.4600 2231.1400 1285.9400 ;
        RECT 2229.5400 1290.9000 2231.1400 1291.3800 ;
        RECT 2229.5400 1269.1400 2231.1400 1269.6200 ;
        RECT 2229.5400 1274.5800 2231.1400 1275.0600 ;
        RECT 2229.5400 1280.0200 2231.1400 1280.5000 ;
        RECT 2184.5400 1296.3400 2186.1400 1296.8200 ;
        RECT 2184.5400 1301.7800 2186.1400 1302.2600 ;
        RECT 2176.7800 1296.3400 2178.3800 1296.8200 ;
        RECT 2176.7800 1301.7800 2178.3800 1302.2600 ;
        RECT 2176.7800 1307.2200 2178.3800 1307.7000 ;
        RECT 2184.5400 1307.2200 2186.1400 1307.7000 ;
        RECT 2184.5400 1285.4600 2186.1400 1285.9400 ;
        RECT 2184.5400 1290.9000 2186.1400 1291.3800 ;
        RECT 2176.7800 1285.4600 2178.3800 1285.9400 ;
        RECT 2176.7800 1290.9000 2178.3800 1291.3800 ;
        RECT 2184.5400 1269.1400 2186.1400 1269.6200 ;
        RECT 2184.5400 1274.5800 2186.1400 1275.0600 ;
        RECT 2176.7800 1269.1400 2178.3800 1269.6200 ;
        RECT 2176.7800 1274.5800 2178.3800 1275.0600 ;
        RECT 2176.7800 1280.0200 2178.3800 1280.5000 ;
        RECT 2184.5400 1280.0200 2186.1400 1280.5000 ;
        RECT 2274.5400 1252.8200 2276.1400 1253.3000 ;
        RECT 2274.5400 1258.2600 2276.1400 1258.7400 ;
        RECT 2274.5400 1263.7000 2276.1400 1264.1800 ;
        RECT 2274.5400 1241.9400 2276.1400 1242.4200 ;
        RECT 2274.5400 1247.3800 2276.1400 1247.8600 ;
        RECT 2229.5400 1252.8200 2231.1400 1253.3000 ;
        RECT 2229.5400 1258.2600 2231.1400 1258.7400 ;
        RECT 2229.5400 1263.7000 2231.1400 1264.1800 ;
        RECT 2229.5400 1241.9400 2231.1400 1242.4200 ;
        RECT 2229.5400 1247.3800 2231.1400 1247.8600 ;
        RECT 2274.5400 1225.6200 2276.1400 1226.1000 ;
        RECT 2274.5400 1231.0600 2276.1400 1231.5400 ;
        RECT 2274.5400 1236.5000 2276.1400 1236.9800 ;
        RECT 2274.5400 1214.7400 2276.1400 1215.2200 ;
        RECT 2274.5400 1220.1800 2276.1400 1220.6600 ;
        RECT 2229.5400 1225.6200 2231.1400 1226.1000 ;
        RECT 2229.5400 1231.0600 2231.1400 1231.5400 ;
        RECT 2229.5400 1236.5000 2231.1400 1236.9800 ;
        RECT 2229.5400 1214.7400 2231.1400 1215.2200 ;
        RECT 2229.5400 1220.1800 2231.1400 1220.6600 ;
        RECT 2184.5400 1252.8200 2186.1400 1253.3000 ;
        RECT 2184.5400 1258.2600 2186.1400 1258.7400 ;
        RECT 2184.5400 1263.7000 2186.1400 1264.1800 ;
        RECT 2176.7800 1252.8200 2178.3800 1253.3000 ;
        RECT 2176.7800 1258.2600 2178.3800 1258.7400 ;
        RECT 2176.7800 1263.7000 2178.3800 1264.1800 ;
        RECT 2184.5400 1241.9400 2186.1400 1242.4200 ;
        RECT 2184.5400 1247.3800 2186.1400 1247.8600 ;
        RECT 2176.7800 1241.9400 2178.3800 1242.4200 ;
        RECT 2176.7800 1247.3800 2178.3800 1247.8600 ;
        RECT 2184.5400 1225.6200 2186.1400 1226.1000 ;
        RECT 2184.5400 1231.0600 2186.1400 1231.5400 ;
        RECT 2184.5400 1236.5000 2186.1400 1236.9800 ;
        RECT 2176.7800 1225.6200 2178.3800 1226.1000 ;
        RECT 2176.7800 1231.0600 2178.3800 1231.5400 ;
        RECT 2176.7800 1236.5000 2178.3800 1236.9800 ;
        RECT 2184.5400 1214.7400 2186.1400 1215.2200 ;
        RECT 2184.5400 1220.1800 2186.1400 1220.6600 ;
        RECT 2176.7800 1214.7400 2178.3800 1215.2200 ;
        RECT 2176.7800 1220.1800 2178.3800 1220.6600 ;
        RECT 2374.2800 1198.4200 2375.8800 1198.9000 ;
        RECT 2374.2800 1203.8600 2375.8800 1204.3400 ;
        RECT 2374.2800 1209.3000 2375.8800 1209.7800 ;
        RECT 2364.5400 1198.4200 2366.1400 1198.9000 ;
        RECT 2364.5400 1203.8600 2366.1400 1204.3400 ;
        RECT 2364.5400 1209.3000 2366.1400 1209.7800 ;
        RECT 2374.2800 1187.5400 2375.8800 1188.0200 ;
        RECT 2374.2800 1192.9800 2375.8800 1193.4600 ;
        RECT 2364.5400 1187.5400 2366.1400 1188.0200 ;
        RECT 2364.5400 1192.9800 2366.1400 1193.4600 ;
        RECT 2374.2800 1171.2200 2375.8800 1171.7000 ;
        RECT 2374.2800 1176.6600 2375.8800 1177.1400 ;
        RECT 2374.2800 1182.1000 2375.8800 1182.5800 ;
        RECT 2364.5400 1171.2200 2366.1400 1171.7000 ;
        RECT 2364.5400 1176.6600 2366.1400 1177.1400 ;
        RECT 2364.5400 1182.1000 2366.1400 1182.5800 ;
        RECT 2374.2800 1160.3400 2375.8800 1160.8200 ;
        RECT 2374.2800 1165.7800 2375.8800 1166.2600 ;
        RECT 2364.5400 1160.3400 2366.1400 1160.8200 ;
        RECT 2364.5400 1165.7800 2366.1400 1166.2600 ;
        RECT 2319.5400 1198.4200 2321.1400 1198.9000 ;
        RECT 2319.5400 1203.8600 2321.1400 1204.3400 ;
        RECT 2319.5400 1209.3000 2321.1400 1209.7800 ;
        RECT 2319.5400 1187.5400 2321.1400 1188.0200 ;
        RECT 2319.5400 1192.9800 2321.1400 1193.4600 ;
        RECT 2319.5400 1171.2200 2321.1400 1171.7000 ;
        RECT 2319.5400 1176.6600 2321.1400 1177.1400 ;
        RECT 2319.5400 1182.1000 2321.1400 1182.5800 ;
        RECT 2319.5400 1160.3400 2321.1400 1160.8200 ;
        RECT 2319.5400 1165.7800 2321.1400 1166.2600 ;
        RECT 2374.2800 1144.0200 2375.8800 1144.5000 ;
        RECT 2374.2800 1149.4600 2375.8800 1149.9400 ;
        RECT 2374.2800 1154.9000 2375.8800 1155.3800 ;
        RECT 2364.5400 1144.0200 2366.1400 1144.5000 ;
        RECT 2364.5400 1149.4600 2366.1400 1149.9400 ;
        RECT 2364.5400 1154.9000 2366.1400 1155.3800 ;
        RECT 2374.2800 1133.1400 2375.8800 1133.6200 ;
        RECT 2374.2800 1138.5800 2375.8800 1139.0600 ;
        RECT 2364.5400 1133.1400 2366.1400 1133.6200 ;
        RECT 2364.5400 1138.5800 2366.1400 1139.0600 ;
        RECT 2374.2800 1116.8200 2375.8800 1117.3000 ;
        RECT 2374.2800 1122.2600 2375.8800 1122.7400 ;
        RECT 2374.2800 1127.7000 2375.8800 1128.1800 ;
        RECT 2364.5400 1116.8200 2366.1400 1117.3000 ;
        RECT 2364.5400 1122.2600 2366.1400 1122.7400 ;
        RECT 2364.5400 1127.7000 2366.1400 1128.1800 ;
        RECT 2364.5400 1111.3800 2366.1400 1111.8600 ;
        RECT 2374.2800 1111.3800 2375.8800 1111.8600 ;
        RECT 2319.5400 1144.0200 2321.1400 1144.5000 ;
        RECT 2319.5400 1149.4600 2321.1400 1149.9400 ;
        RECT 2319.5400 1154.9000 2321.1400 1155.3800 ;
        RECT 2319.5400 1133.1400 2321.1400 1133.6200 ;
        RECT 2319.5400 1138.5800 2321.1400 1139.0600 ;
        RECT 2319.5400 1116.8200 2321.1400 1117.3000 ;
        RECT 2319.5400 1122.2600 2321.1400 1122.7400 ;
        RECT 2319.5400 1127.7000 2321.1400 1128.1800 ;
        RECT 2319.5400 1111.3800 2321.1400 1111.8600 ;
        RECT 2274.5400 1198.4200 2276.1400 1198.9000 ;
        RECT 2274.5400 1203.8600 2276.1400 1204.3400 ;
        RECT 2274.5400 1209.3000 2276.1400 1209.7800 ;
        RECT 2274.5400 1187.5400 2276.1400 1188.0200 ;
        RECT 2274.5400 1192.9800 2276.1400 1193.4600 ;
        RECT 2229.5400 1198.4200 2231.1400 1198.9000 ;
        RECT 2229.5400 1203.8600 2231.1400 1204.3400 ;
        RECT 2229.5400 1209.3000 2231.1400 1209.7800 ;
        RECT 2229.5400 1187.5400 2231.1400 1188.0200 ;
        RECT 2229.5400 1192.9800 2231.1400 1193.4600 ;
        RECT 2274.5400 1171.2200 2276.1400 1171.7000 ;
        RECT 2274.5400 1176.6600 2276.1400 1177.1400 ;
        RECT 2274.5400 1182.1000 2276.1400 1182.5800 ;
        RECT 2274.5400 1160.3400 2276.1400 1160.8200 ;
        RECT 2274.5400 1165.7800 2276.1400 1166.2600 ;
        RECT 2229.5400 1171.2200 2231.1400 1171.7000 ;
        RECT 2229.5400 1176.6600 2231.1400 1177.1400 ;
        RECT 2229.5400 1182.1000 2231.1400 1182.5800 ;
        RECT 2229.5400 1160.3400 2231.1400 1160.8200 ;
        RECT 2229.5400 1165.7800 2231.1400 1166.2600 ;
        RECT 2184.5400 1198.4200 2186.1400 1198.9000 ;
        RECT 2184.5400 1203.8600 2186.1400 1204.3400 ;
        RECT 2184.5400 1209.3000 2186.1400 1209.7800 ;
        RECT 2176.7800 1198.4200 2178.3800 1198.9000 ;
        RECT 2176.7800 1203.8600 2178.3800 1204.3400 ;
        RECT 2176.7800 1209.3000 2178.3800 1209.7800 ;
        RECT 2184.5400 1187.5400 2186.1400 1188.0200 ;
        RECT 2184.5400 1192.9800 2186.1400 1193.4600 ;
        RECT 2176.7800 1187.5400 2178.3800 1188.0200 ;
        RECT 2176.7800 1192.9800 2178.3800 1193.4600 ;
        RECT 2184.5400 1171.2200 2186.1400 1171.7000 ;
        RECT 2184.5400 1176.6600 2186.1400 1177.1400 ;
        RECT 2184.5400 1182.1000 2186.1400 1182.5800 ;
        RECT 2176.7800 1171.2200 2178.3800 1171.7000 ;
        RECT 2176.7800 1176.6600 2178.3800 1177.1400 ;
        RECT 2176.7800 1182.1000 2178.3800 1182.5800 ;
        RECT 2184.5400 1160.3400 2186.1400 1160.8200 ;
        RECT 2184.5400 1165.7800 2186.1400 1166.2600 ;
        RECT 2176.7800 1160.3400 2178.3800 1160.8200 ;
        RECT 2176.7800 1165.7800 2178.3800 1166.2600 ;
        RECT 2274.5400 1144.0200 2276.1400 1144.5000 ;
        RECT 2274.5400 1149.4600 2276.1400 1149.9400 ;
        RECT 2274.5400 1154.9000 2276.1400 1155.3800 ;
        RECT 2274.5400 1133.1400 2276.1400 1133.6200 ;
        RECT 2274.5400 1138.5800 2276.1400 1139.0600 ;
        RECT 2229.5400 1144.0200 2231.1400 1144.5000 ;
        RECT 2229.5400 1149.4600 2231.1400 1149.9400 ;
        RECT 2229.5400 1154.9000 2231.1400 1155.3800 ;
        RECT 2229.5400 1133.1400 2231.1400 1133.6200 ;
        RECT 2229.5400 1138.5800 2231.1400 1139.0600 ;
        RECT 2274.5400 1116.8200 2276.1400 1117.3000 ;
        RECT 2274.5400 1122.2600 2276.1400 1122.7400 ;
        RECT 2274.5400 1127.7000 2276.1400 1128.1800 ;
        RECT 2274.5400 1111.3800 2276.1400 1111.8600 ;
        RECT 2229.5400 1116.8200 2231.1400 1117.3000 ;
        RECT 2229.5400 1122.2600 2231.1400 1122.7400 ;
        RECT 2229.5400 1127.7000 2231.1400 1128.1800 ;
        RECT 2229.5400 1111.3800 2231.1400 1111.8600 ;
        RECT 2184.5400 1144.0200 2186.1400 1144.5000 ;
        RECT 2184.5400 1149.4600 2186.1400 1149.9400 ;
        RECT 2184.5400 1154.9000 2186.1400 1155.3800 ;
        RECT 2176.7800 1144.0200 2178.3800 1144.5000 ;
        RECT 2176.7800 1149.4600 2178.3800 1149.9400 ;
        RECT 2176.7800 1154.9000 2178.3800 1155.3800 ;
        RECT 2184.5400 1133.1400 2186.1400 1133.6200 ;
        RECT 2184.5400 1138.5800 2186.1400 1139.0600 ;
        RECT 2176.7800 1133.1400 2178.3800 1133.6200 ;
        RECT 2176.7800 1138.5800 2178.3800 1139.0600 ;
        RECT 2184.5400 1116.8200 2186.1400 1117.3000 ;
        RECT 2184.5400 1122.2600 2186.1400 1122.7400 ;
        RECT 2184.5400 1127.7000 2186.1400 1128.1800 ;
        RECT 2176.7800 1116.8200 2178.3800 1117.3000 ;
        RECT 2176.7800 1122.2600 2178.3800 1122.7400 ;
        RECT 2176.7800 1127.7000 2178.3800 1128.1800 ;
        RECT 2176.7800 1111.3800 2178.3800 1111.8600 ;
        RECT 2184.5400 1111.3800 2186.1400 1111.8600 ;
        RECT 2171.2200 1313.6900 2381.4400 1315.2900 ;
        RECT 2171.2200 1107.1900 2381.4400 1108.7900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1101.7600 2178.3800 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1319.8000 2178.3800 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1101.7600 2375.8800 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1319.8000 2375.8800 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1107.1900 2172.8200 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1107.1900 2381.4400 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1313.6900 2172.8200 1315.2900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1313.6900 2381.4400 1315.2900 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 877.5500 2366.1400 1085.6500 ;
        RECT 2319.5400 877.5500 2321.1400 1085.6500 ;
        RECT 2274.5400 877.5500 2276.1400 1085.6500 ;
        RECT 2229.5400 877.5500 2231.1400 1085.6500 ;
        RECT 2184.5400 877.5500 2186.1400 1085.6500 ;
        RECT 2374.2800 872.1200 2375.8800 1091.7600 ;
        RECT 2176.7800 872.1200 2178.3800 1091.7600 ;
      LAYER met3 ;
        RECT 2374.2800 1066.7000 2375.8800 1067.1800 ;
        RECT 2374.2800 1072.1400 2375.8800 1072.6200 ;
        RECT 2364.5400 1066.7000 2366.1400 1067.1800 ;
        RECT 2364.5400 1072.1400 2366.1400 1072.6200 ;
        RECT 2364.5400 1077.5800 2366.1400 1078.0600 ;
        RECT 2374.2800 1077.5800 2375.8800 1078.0600 ;
        RECT 2374.2800 1055.8200 2375.8800 1056.3000 ;
        RECT 2374.2800 1061.2600 2375.8800 1061.7400 ;
        RECT 2364.5400 1055.8200 2366.1400 1056.3000 ;
        RECT 2364.5400 1061.2600 2366.1400 1061.7400 ;
        RECT 2374.2800 1039.5000 2375.8800 1039.9800 ;
        RECT 2374.2800 1044.9400 2375.8800 1045.4200 ;
        RECT 2364.5400 1039.5000 2366.1400 1039.9800 ;
        RECT 2364.5400 1044.9400 2366.1400 1045.4200 ;
        RECT 2364.5400 1050.3800 2366.1400 1050.8600 ;
        RECT 2374.2800 1050.3800 2375.8800 1050.8600 ;
        RECT 2319.5400 1066.7000 2321.1400 1067.1800 ;
        RECT 2319.5400 1072.1400 2321.1400 1072.6200 ;
        RECT 2319.5400 1077.5800 2321.1400 1078.0600 ;
        RECT 2319.5400 1055.8200 2321.1400 1056.3000 ;
        RECT 2319.5400 1061.2600 2321.1400 1061.7400 ;
        RECT 2319.5400 1039.5000 2321.1400 1039.9800 ;
        RECT 2319.5400 1044.9400 2321.1400 1045.4200 ;
        RECT 2319.5400 1050.3800 2321.1400 1050.8600 ;
        RECT 2374.2800 1023.1800 2375.8800 1023.6600 ;
        RECT 2374.2800 1028.6200 2375.8800 1029.1000 ;
        RECT 2374.2800 1034.0600 2375.8800 1034.5400 ;
        RECT 2364.5400 1023.1800 2366.1400 1023.6600 ;
        RECT 2364.5400 1028.6200 2366.1400 1029.1000 ;
        RECT 2364.5400 1034.0600 2366.1400 1034.5400 ;
        RECT 2374.2800 1012.3000 2375.8800 1012.7800 ;
        RECT 2374.2800 1017.7400 2375.8800 1018.2200 ;
        RECT 2364.5400 1012.3000 2366.1400 1012.7800 ;
        RECT 2364.5400 1017.7400 2366.1400 1018.2200 ;
        RECT 2374.2800 995.9800 2375.8800 996.4600 ;
        RECT 2374.2800 1001.4200 2375.8800 1001.9000 ;
        RECT 2374.2800 1006.8600 2375.8800 1007.3400 ;
        RECT 2364.5400 995.9800 2366.1400 996.4600 ;
        RECT 2364.5400 1001.4200 2366.1400 1001.9000 ;
        RECT 2364.5400 1006.8600 2366.1400 1007.3400 ;
        RECT 2374.2800 985.1000 2375.8800 985.5800 ;
        RECT 2374.2800 990.5400 2375.8800 991.0200 ;
        RECT 2364.5400 985.1000 2366.1400 985.5800 ;
        RECT 2364.5400 990.5400 2366.1400 991.0200 ;
        RECT 2319.5400 1023.1800 2321.1400 1023.6600 ;
        RECT 2319.5400 1028.6200 2321.1400 1029.1000 ;
        RECT 2319.5400 1034.0600 2321.1400 1034.5400 ;
        RECT 2319.5400 1012.3000 2321.1400 1012.7800 ;
        RECT 2319.5400 1017.7400 2321.1400 1018.2200 ;
        RECT 2319.5400 995.9800 2321.1400 996.4600 ;
        RECT 2319.5400 1001.4200 2321.1400 1001.9000 ;
        RECT 2319.5400 1006.8600 2321.1400 1007.3400 ;
        RECT 2319.5400 985.1000 2321.1400 985.5800 ;
        RECT 2319.5400 990.5400 2321.1400 991.0200 ;
        RECT 2274.5400 1066.7000 2276.1400 1067.1800 ;
        RECT 2274.5400 1072.1400 2276.1400 1072.6200 ;
        RECT 2274.5400 1077.5800 2276.1400 1078.0600 ;
        RECT 2229.5400 1066.7000 2231.1400 1067.1800 ;
        RECT 2229.5400 1072.1400 2231.1400 1072.6200 ;
        RECT 2229.5400 1077.5800 2231.1400 1078.0600 ;
        RECT 2274.5400 1055.8200 2276.1400 1056.3000 ;
        RECT 2274.5400 1061.2600 2276.1400 1061.7400 ;
        RECT 2274.5400 1039.5000 2276.1400 1039.9800 ;
        RECT 2274.5400 1044.9400 2276.1400 1045.4200 ;
        RECT 2274.5400 1050.3800 2276.1400 1050.8600 ;
        RECT 2229.5400 1055.8200 2231.1400 1056.3000 ;
        RECT 2229.5400 1061.2600 2231.1400 1061.7400 ;
        RECT 2229.5400 1039.5000 2231.1400 1039.9800 ;
        RECT 2229.5400 1044.9400 2231.1400 1045.4200 ;
        RECT 2229.5400 1050.3800 2231.1400 1050.8600 ;
        RECT 2184.5400 1066.7000 2186.1400 1067.1800 ;
        RECT 2184.5400 1072.1400 2186.1400 1072.6200 ;
        RECT 2176.7800 1066.7000 2178.3800 1067.1800 ;
        RECT 2176.7800 1072.1400 2178.3800 1072.6200 ;
        RECT 2176.7800 1077.5800 2178.3800 1078.0600 ;
        RECT 2184.5400 1077.5800 2186.1400 1078.0600 ;
        RECT 2184.5400 1055.8200 2186.1400 1056.3000 ;
        RECT 2184.5400 1061.2600 2186.1400 1061.7400 ;
        RECT 2176.7800 1055.8200 2178.3800 1056.3000 ;
        RECT 2176.7800 1061.2600 2178.3800 1061.7400 ;
        RECT 2184.5400 1039.5000 2186.1400 1039.9800 ;
        RECT 2184.5400 1044.9400 2186.1400 1045.4200 ;
        RECT 2176.7800 1039.5000 2178.3800 1039.9800 ;
        RECT 2176.7800 1044.9400 2178.3800 1045.4200 ;
        RECT 2176.7800 1050.3800 2178.3800 1050.8600 ;
        RECT 2184.5400 1050.3800 2186.1400 1050.8600 ;
        RECT 2274.5400 1023.1800 2276.1400 1023.6600 ;
        RECT 2274.5400 1028.6200 2276.1400 1029.1000 ;
        RECT 2274.5400 1034.0600 2276.1400 1034.5400 ;
        RECT 2274.5400 1012.3000 2276.1400 1012.7800 ;
        RECT 2274.5400 1017.7400 2276.1400 1018.2200 ;
        RECT 2229.5400 1023.1800 2231.1400 1023.6600 ;
        RECT 2229.5400 1028.6200 2231.1400 1029.1000 ;
        RECT 2229.5400 1034.0600 2231.1400 1034.5400 ;
        RECT 2229.5400 1012.3000 2231.1400 1012.7800 ;
        RECT 2229.5400 1017.7400 2231.1400 1018.2200 ;
        RECT 2274.5400 995.9800 2276.1400 996.4600 ;
        RECT 2274.5400 1001.4200 2276.1400 1001.9000 ;
        RECT 2274.5400 1006.8600 2276.1400 1007.3400 ;
        RECT 2274.5400 985.1000 2276.1400 985.5800 ;
        RECT 2274.5400 990.5400 2276.1400 991.0200 ;
        RECT 2229.5400 995.9800 2231.1400 996.4600 ;
        RECT 2229.5400 1001.4200 2231.1400 1001.9000 ;
        RECT 2229.5400 1006.8600 2231.1400 1007.3400 ;
        RECT 2229.5400 985.1000 2231.1400 985.5800 ;
        RECT 2229.5400 990.5400 2231.1400 991.0200 ;
        RECT 2184.5400 1023.1800 2186.1400 1023.6600 ;
        RECT 2184.5400 1028.6200 2186.1400 1029.1000 ;
        RECT 2184.5400 1034.0600 2186.1400 1034.5400 ;
        RECT 2176.7800 1023.1800 2178.3800 1023.6600 ;
        RECT 2176.7800 1028.6200 2178.3800 1029.1000 ;
        RECT 2176.7800 1034.0600 2178.3800 1034.5400 ;
        RECT 2184.5400 1012.3000 2186.1400 1012.7800 ;
        RECT 2184.5400 1017.7400 2186.1400 1018.2200 ;
        RECT 2176.7800 1012.3000 2178.3800 1012.7800 ;
        RECT 2176.7800 1017.7400 2178.3800 1018.2200 ;
        RECT 2184.5400 995.9800 2186.1400 996.4600 ;
        RECT 2184.5400 1001.4200 2186.1400 1001.9000 ;
        RECT 2184.5400 1006.8600 2186.1400 1007.3400 ;
        RECT 2176.7800 995.9800 2178.3800 996.4600 ;
        RECT 2176.7800 1001.4200 2178.3800 1001.9000 ;
        RECT 2176.7800 1006.8600 2178.3800 1007.3400 ;
        RECT 2184.5400 985.1000 2186.1400 985.5800 ;
        RECT 2184.5400 990.5400 2186.1400 991.0200 ;
        RECT 2176.7800 985.1000 2178.3800 985.5800 ;
        RECT 2176.7800 990.5400 2178.3800 991.0200 ;
        RECT 2374.2800 968.7800 2375.8800 969.2600 ;
        RECT 2374.2800 974.2200 2375.8800 974.7000 ;
        RECT 2374.2800 979.6600 2375.8800 980.1400 ;
        RECT 2364.5400 968.7800 2366.1400 969.2600 ;
        RECT 2364.5400 974.2200 2366.1400 974.7000 ;
        RECT 2364.5400 979.6600 2366.1400 980.1400 ;
        RECT 2374.2800 957.9000 2375.8800 958.3800 ;
        RECT 2374.2800 963.3400 2375.8800 963.8200 ;
        RECT 2364.5400 957.9000 2366.1400 958.3800 ;
        RECT 2364.5400 963.3400 2366.1400 963.8200 ;
        RECT 2374.2800 941.5800 2375.8800 942.0600 ;
        RECT 2374.2800 947.0200 2375.8800 947.5000 ;
        RECT 2374.2800 952.4600 2375.8800 952.9400 ;
        RECT 2364.5400 941.5800 2366.1400 942.0600 ;
        RECT 2364.5400 947.0200 2366.1400 947.5000 ;
        RECT 2364.5400 952.4600 2366.1400 952.9400 ;
        RECT 2374.2800 930.7000 2375.8800 931.1800 ;
        RECT 2374.2800 936.1400 2375.8800 936.6200 ;
        RECT 2364.5400 930.7000 2366.1400 931.1800 ;
        RECT 2364.5400 936.1400 2366.1400 936.6200 ;
        RECT 2319.5400 968.7800 2321.1400 969.2600 ;
        RECT 2319.5400 974.2200 2321.1400 974.7000 ;
        RECT 2319.5400 979.6600 2321.1400 980.1400 ;
        RECT 2319.5400 957.9000 2321.1400 958.3800 ;
        RECT 2319.5400 963.3400 2321.1400 963.8200 ;
        RECT 2319.5400 941.5800 2321.1400 942.0600 ;
        RECT 2319.5400 947.0200 2321.1400 947.5000 ;
        RECT 2319.5400 952.4600 2321.1400 952.9400 ;
        RECT 2319.5400 930.7000 2321.1400 931.1800 ;
        RECT 2319.5400 936.1400 2321.1400 936.6200 ;
        RECT 2374.2800 914.3800 2375.8800 914.8600 ;
        RECT 2374.2800 919.8200 2375.8800 920.3000 ;
        RECT 2374.2800 925.2600 2375.8800 925.7400 ;
        RECT 2364.5400 914.3800 2366.1400 914.8600 ;
        RECT 2364.5400 919.8200 2366.1400 920.3000 ;
        RECT 2364.5400 925.2600 2366.1400 925.7400 ;
        RECT 2374.2800 903.5000 2375.8800 903.9800 ;
        RECT 2374.2800 908.9400 2375.8800 909.4200 ;
        RECT 2364.5400 903.5000 2366.1400 903.9800 ;
        RECT 2364.5400 908.9400 2366.1400 909.4200 ;
        RECT 2374.2800 887.1800 2375.8800 887.6600 ;
        RECT 2374.2800 892.6200 2375.8800 893.1000 ;
        RECT 2374.2800 898.0600 2375.8800 898.5400 ;
        RECT 2364.5400 887.1800 2366.1400 887.6600 ;
        RECT 2364.5400 892.6200 2366.1400 893.1000 ;
        RECT 2364.5400 898.0600 2366.1400 898.5400 ;
        RECT 2364.5400 881.7400 2366.1400 882.2200 ;
        RECT 2374.2800 881.7400 2375.8800 882.2200 ;
        RECT 2319.5400 914.3800 2321.1400 914.8600 ;
        RECT 2319.5400 919.8200 2321.1400 920.3000 ;
        RECT 2319.5400 925.2600 2321.1400 925.7400 ;
        RECT 2319.5400 903.5000 2321.1400 903.9800 ;
        RECT 2319.5400 908.9400 2321.1400 909.4200 ;
        RECT 2319.5400 887.1800 2321.1400 887.6600 ;
        RECT 2319.5400 892.6200 2321.1400 893.1000 ;
        RECT 2319.5400 898.0600 2321.1400 898.5400 ;
        RECT 2319.5400 881.7400 2321.1400 882.2200 ;
        RECT 2274.5400 968.7800 2276.1400 969.2600 ;
        RECT 2274.5400 974.2200 2276.1400 974.7000 ;
        RECT 2274.5400 979.6600 2276.1400 980.1400 ;
        RECT 2274.5400 957.9000 2276.1400 958.3800 ;
        RECT 2274.5400 963.3400 2276.1400 963.8200 ;
        RECT 2229.5400 968.7800 2231.1400 969.2600 ;
        RECT 2229.5400 974.2200 2231.1400 974.7000 ;
        RECT 2229.5400 979.6600 2231.1400 980.1400 ;
        RECT 2229.5400 957.9000 2231.1400 958.3800 ;
        RECT 2229.5400 963.3400 2231.1400 963.8200 ;
        RECT 2274.5400 941.5800 2276.1400 942.0600 ;
        RECT 2274.5400 947.0200 2276.1400 947.5000 ;
        RECT 2274.5400 952.4600 2276.1400 952.9400 ;
        RECT 2274.5400 930.7000 2276.1400 931.1800 ;
        RECT 2274.5400 936.1400 2276.1400 936.6200 ;
        RECT 2229.5400 941.5800 2231.1400 942.0600 ;
        RECT 2229.5400 947.0200 2231.1400 947.5000 ;
        RECT 2229.5400 952.4600 2231.1400 952.9400 ;
        RECT 2229.5400 930.7000 2231.1400 931.1800 ;
        RECT 2229.5400 936.1400 2231.1400 936.6200 ;
        RECT 2184.5400 968.7800 2186.1400 969.2600 ;
        RECT 2184.5400 974.2200 2186.1400 974.7000 ;
        RECT 2184.5400 979.6600 2186.1400 980.1400 ;
        RECT 2176.7800 968.7800 2178.3800 969.2600 ;
        RECT 2176.7800 974.2200 2178.3800 974.7000 ;
        RECT 2176.7800 979.6600 2178.3800 980.1400 ;
        RECT 2184.5400 957.9000 2186.1400 958.3800 ;
        RECT 2184.5400 963.3400 2186.1400 963.8200 ;
        RECT 2176.7800 957.9000 2178.3800 958.3800 ;
        RECT 2176.7800 963.3400 2178.3800 963.8200 ;
        RECT 2184.5400 941.5800 2186.1400 942.0600 ;
        RECT 2184.5400 947.0200 2186.1400 947.5000 ;
        RECT 2184.5400 952.4600 2186.1400 952.9400 ;
        RECT 2176.7800 941.5800 2178.3800 942.0600 ;
        RECT 2176.7800 947.0200 2178.3800 947.5000 ;
        RECT 2176.7800 952.4600 2178.3800 952.9400 ;
        RECT 2184.5400 930.7000 2186.1400 931.1800 ;
        RECT 2184.5400 936.1400 2186.1400 936.6200 ;
        RECT 2176.7800 930.7000 2178.3800 931.1800 ;
        RECT 2176.7800 936.1400 2178.3800 936.6200 ;
        RECT 2274.5400 914.3800 2276.1400 914.8600 ;
        RECT 2274.5400 919.8200 2276.1400 920.3000 ;
        RECT 2274.5400 925.2600 2276.1400 925.7400 ;
        RECT 2274.5400 903.5000 2276.1400 903.9800 ;
        RECT 2274.5400 908.9400 2276.1400 909.4200 ;
        RECT 2229.5400 914.3800 2231.1400 914.8600 ;
        RECT 2229.5400 919.8200 2231.1400 920.3000 ;
        RECT 2229.5400 925.2600 2231.1400 925.7400 ;
        RECT 2229.5400 903.5000 2231.1400 903.9800 ;
        RECT 2229.5400 908.9400 2231.1400 909.4200 ;
        RECT 2274.5400 887.1800 2276.1400 887.6600 ;
        RECT 2274.5400 892.6200 2276.1400 893.1000 ;
        RECT 2274.5400 898.0600 2276.1400 898.5400 ;
        RECT 2274.5400 881.7400 2276.1400 882.2200 ;
        RECT 2229.5400 887.1800 2231.1400 887.6600 ;
        RECT 2229.5400 892.6200 2231.1400 893.1000 ;
        RECT 2229.5400 898.0600 2231.1400 898.5400 ;
        RECT 2229.5400 881.7400 2231.1400 882.2200 ;
        RECT 2184.5400 914.3800 2186.1400 914.8600 ;
        RECT 2184.5400 919.8200 2186.1400 920.3000 ;
        RECT 2184.5400 925.2600 2186.1400 925.7400 ;
        RECT 2176.7800 914.3800 2178.3800 914.8600 ;
        RECT 2176.7800 919.8200 2178.3800 920.3000 ;
        RECT 2176.7800 925.2600 2178.3800 925.7400 ;
        RECT 2184.5400 903.5000 2186.1400 903.9800 ;
        RECT 2184.5400 908.9400 2186.1400 909.4200 ;
        RECT 2176.7800 903.5000 2178.3800 903.9800 ;
        RECT 2176.7800 908.9400 2178.3800 909.4200 ;
        RECT 2184.5400 887.1800 2186.1400 887.6600 ;
        RECT 2184.5400 892.6200 2186.1400 893.1000 ;
        RECT 2184.5400 898.0600 2186.1400 898.5400 ;
        RECT 2176.7800 887.1800 2178.3800 887.6600 ;
        RECT 2176.7800 892.6200 2178.3800 893.1000 ;
        RECT 2176.7800 898.0600 2178.3800 898.5400 ;
        RECT 2176.7800 881.7400 2178.3800 882.2200 ;
        RECT 2184.5400 881.7400 2186.1400 882.2200 ;
        RECT 2171.2200 1084.0500 2381.4400 1085.6500 ;
        RECT 2171.2200 877.5500 2381.4400 879.1500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 872.1200 2178.3800 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 1090.1600 2178.3800 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 872.1200 2375.8800 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 1090.1600 2375.8800 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 877.5500 2172.8200 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 877.5500 2381.4400 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 1084.0500 2172.8200 1085.6500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 1084.0500 2381.4400 1085.6500 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 647.9100 2366.1400 856.0100 ;
        RECT 2319.5400 647.9100 2321.1400 856.0100 ;
        RECT 2274.5400 647.9100 2276.1400 856.0100 ;
        RECT 2229.5400 647.9100 2231.1400 856.0100 ;
        RECT 2184.5400 647.9100 2186.1400 856.0100 ;
        RECT 2374.2800 642.4800 2375.8800 862.1200 ;
        RECT 2176.7800 642.4800 2178.3800 862.1200 ;
      LAYER met3 ;
        RECT 2374.2800 837.0600 2375.8800 837.5400 ;
        RECT 2374.2800 842.5000 2375.8800 842.9800 ;
        RECT 2364.5400 837.0600 2366.1400 837.5400 ;
        RECT 2364.5400 842.5000 2366.1400 842.9800 ;
        RECT 2364.5400 847.9400 2366.1400 848.4200 ;
        RECT 2374.2800 847.9400 2375.8800 848.4200 ;
        RECT 2374.2800 826.1800 2375.8800 826.6600 ;
        RECT 2374.2800 831.6200 2375.8800 832.1000 ;
        RECT 2364.5400 826.1800 2366.1400 826.6600 ;
        RECT 2364.5400 831.6200 2366.1400 832.1000 ;
        RECT 2374.2800 809.8600 2375.8800 810.3400 ;
        RECT 2374.2800 815.3000 2375.8800 815.7800 ;
        RECT 2364.5400 809.8600 2366.1400 810.3400 ;
        RECT 2364.5400 815.3000 2366.1400 815.7800 ;
        RECT 2364.5400 820.7400 2366.1400 821.2200 ;
        RECT 2374.2800 820.7400 2375.8800 821.2200 ;
        RECT 2319.5400 837.0600 2321.1400 837.5400 ;
        RECT 2319.5400 842.5000 2321.1400 842.9800 ;
        RECT 2319.5400 847.9400 2321.1400 848.4200 ;
        RECT 2319.5400 826.1800 2321.1400 826.6600 ;
        RECT 2319.5400 831.6200 2321.1400 832.1000 ;
        RECT 2319.5400 809.8600 2321.1400 810.3400 ;
        RECT 2319.5400 815.3000 2321.1400 815.7800 ;
        RECT 2319.5400 820.7400 2321.1400 821.2200 ;
        RECT 2374.2800 793.5400 2375.8800 794.0200 ;
        RECT 2374.2800 798.9800 2375.8800 799.4600 ;
        RECT 2374.2800 804.4200 2375.8800 804.9000 ;
        RECT 2364.5400 793.5400 2366.1400 794.0200 ;
        RECT 2364.5400 798.9800 2366.1400 799.4600 ;
        RECT 2364.5400 804.4200 2366.1400 804.9000 ;
        RECT 2374.2800 782.6600 2375.8800 783.1400 ;
        RECT 2374.2800 788.1000 2375.8800 788.5800 ;
        RECT 2364.5400 782.6600 2366.1400 783.1400 ;
        RECT 2364.5400 788.1000 2366.1400 788.5800 ;
        RECT 2374.2800 766.3400 2375.8800 766.8200 ;
        RECT 2374.2800 771.7800 2375.8800 772.2600 ;
        RECT 2374.2800 777.2200 2375.8800 777.7000 ;
        RECT 2364.5400 766.3400 2366.1400 766.8200 ;
        RECT 2364.5400 771.7800 2366.1400 772.2600 ;
        RECT 2364.5400 777.2200 2366.1400 777.7000 ;
        RECT 2374.2800 755.4600 2375.8800 755.9400 ;
        RECT 2374.2800 760.9000 2375.8800 761.3800 ;
        RECT 2364.5400 755.4600 2366.1400 755.9400 ;
        RECT 2364.5400 760.9000 2366.1400 761.3800 ;
        RECT 2319.5400 793.5400 2321.1400 794.0200 ;
        RECT 2319.5400 798.9800 2321.1400 799.4600 ;
        RECT 2319.5400 804.4200 2321.1400 804.9000 ;
        RECT 2319.5400 782.6600 2321.1400 783.1400 ;
        RECT 2319.5400 788.1000 2321.1400 788.5800 ;
        RECT 2319.5400 766.3400 2321.1400 766.8200 ;
        RECT 2319.5400 771.7800 2321.1400 772.2600 ;
        RECT 2319.5400 777.2200 2321.1400 777.7000 ;
        RECT 2319.5400 755.4600 2321.1400 755.9400 ;
        RECT 2319.5400 760.9000 2321.1400 761.3800 ;
        RECT 2274.5400 837.0600 2276.1400 837.5400 ;
        RECT 2274.5400 842.5000 2276.1400 842.9800 ;
        RECT 2274.5400 847.9400 2276.1400 848.4200 ;
        RECT 2229.5400 837.0600 2231.1400 837.5400 ;
        RECT 2229.5400 842.5000 2231.1400 842.9800 ;
        RECT 2229.5400 847.9400 2231.1400 848.4200 ;
        RECT 2274.5400 826.1800 2276.1400 826.6600 ;
        RECT 2274.5400 831.6200 2276.1400 832.1000 ;
        RECT 2274.5400 809.8600 2276.1400 810.3400 ;
        RECT 2274.5400 815.3000 2276.1400 815.7800 ;
        RECT 2274.5400 820.7400 2276.1400 821.2200 ;
        RECT 2229.5400 826.1800 2231.1400 826.6600 ;
        RECT 2229.5400 831.6200 2231.1400 832.1000 ;
        RECT 2229.5400 809.8600 2231.1400 810.3400 ;
        RECT 2229.5400 815.3000 2231.1400 815.7800 ;
        RECT 2229.5400 820.7400 2231.1400 821.2200 ;
        RECT 2184.5400 837.0600 2186.1400 837.5400 ;
        RECT 2184.5400 842.5000 2186.1400 842.9800 ;
        RECT 2176.7800 837.0600 2178.3800 837.5400 ;
        RECT 2176.7800 842.5000 2178.3800 842.9800 ;
        RECT 2176.7800 847.9400 2178.3800 848.4200 ;
        RECT 2184.5400 847.9400 2186.1400 848.4200 ;
        RECT 2184.5400 826.1800 2186.1400 826.6600 ;
        RECT 2184.5400 831.6200 2186.1400 832.1000 ;
        RECT 2176.7800 826.1800 2178.3800 826.6600 ;
        RECT 2176.7800 831.6200 2178.3800 832.1000 ;
        RECT 2184.5400 809.8600 2186.1400 810.3400 ;
        RECT 2184.5400 815.3000 2186.1400 815.7800 ;
        RECT 2176.7800 809.8600 2178.3800 810.3400 ;
        RECT 2176.7800 815.3000 2178.3800 815.7800 ;
        RECT 2176.7800 820.7400 2178.3800 821.2200 ;
        RECT 2184.5400 820.7400 2186.1400 821.2200 ;
        RECT 2274.5400 793.5400 2276.1400 794.0200 ;
        RECT 2274.5400 798.9800 2276.1400 799.4600 ;
        RECT 2274.5400 804.4200 2276.1400 804.9000 ;
        RECT 2274.5400 782.6600 2276.1400 783.1400 ;
        RECT 2274.5400 788.1000 2276.1400 788.5800 ;
        RECT 2229.5400 793.5400 2231.1400 794.0200 ;
        RECT 2229.5400 798.9800 2231.1400 799.4600 ;
        RECT 2229.5400 804.4200 2231.1400 804.9000 ;
        RECT 2229.5400 782.6600 2231.1400 783.1400 ;
        RECT 2229.5400 788.1000 2231.1400 788.5800 ;
        RECT 2274.5400 766.3400 2276.1400 766.8200 ;
        RECT 2274.5400 771.7800 2276.1400 772.2600 ;
        RECT 2274.5400 777.2200 2276.1400 777.7000 ;
        RECT 2274.5400 755.4600 2276.1400 755.9400 ;
        RECT 2274.5400 760.9000 2276.1400 761.3800 ;
        RECT 2229.5400 766.3400 2231.1400 766.8200 ;
        RECT 2229.5400 771.7800 2231.1400 772.2600 ;
        RECT 2229.5400 777.2200 2231.1400 777.7000 ;
        RECT 2229.5400 755.4600 2231.1400 755.9400 ;
        RECT 2229.5400 760.9000 2231.1400 761.3800 ;
        RECT 2184.5400 793.5400 2186.1400 794.0200 ;
        RECT 2184.5400 798.9800 2186.1400 799.4600 ;
        RECT 2184.5400 804.4200 2186.1400 804.9000 ;
        RECT 2176.7800 793.5400 2178.3800 794.0200 ;
        RECT 2176.7800 798.9800 2178.3800 799.4600 ;
        RECT 2176.7800 804.4200 2178.3800 804.9000 ;
        RECT 2184.5400 782.6600 2186.1400 783.1400 ;
        RECT 2184.5400 788.1000 2186.1400 788.5800 ;
        RECT 2176.7800 782.6600 2178.3800 783.1400 ;
        RECT 2176.7800 788.1000 2178.3800 788.5800 ;
        RECT 2184.5400 766.3400 2186.1400 766.8200 ;
        RECT 2184.5400 771.7800 2186.1400 772.2600 ;
        RECT 2184.5400 777.2200 2186.1400 777.7000 ;
        RECT 2176.7800 766.3400 2178.3800 766.8200 ;
        RECT 2176.7800 771.7800 2178.3800 772.2600 ;
        RECT 2176.7800 777.2200 2178.3800 777.7000 ;
        RECT 2184.5400 755.4600 2186.1400 755.9400 ;
        RECT 2184.5400 760.9000 2186.1400 761.3800 ;
        RECT 2176.7800 755.4600 2178.3800 755.9400 ;
        RECT 2176.7800 760.9000 2178.3800 761.3800 ;
        RECT 2374.2800 739.1400 2375.8800 739.6200 ;
        RECT 2374.2800 744.5800 2375.8800 745.0600 ;
        RECT 2374.2800 750.0200 2375.8800 750.5000 ;
        RECT 2364.5400 739.1400 2366.1400 739.6200 ;
        RECT 2364.5400 744.5800 2366.1400 745.0600 ;
        RECT 2364.5400 750.0200 2366.1400 750.5000 ;
        RECT 2374.2800 728.2600 2375.8800 728.7400 ;
        RECT 2374.2800 733.7000 2375.8800 734.1800 ;
        RECT 2364.5400 728.2600 2366.1400 728.7400 ;
        RECT 2364.5400 733.7000 2366.1400 734.1800 ;
        RECT 2374.2800 711.9400 2375.8800 712.4200 ;
        RECT 2374.2800 717.3800 2375.8800 717.8600 ;
        RECT 2374.2800 722.8200 2375.8800 723.3000 ;
        RECT 2364.5400 711.9400 2366.1400 712.4200 ;
        RECT 2364.5400 717.3800 2366.1400 717.8600 ;
        RECT 2364.5400 722.8200 2366.1400 723.3000 ;
        RECT 2374.2800 701.0600 2375.8800 701.5400 ;
        RECT 2374.2800 706.5000 2375.8800 706.9800 ;
        RECT 2364.5400 701.0600 2366.1400 701.5400 ;
        RECT 2364.5400 706.5000 2366.1400 706.9800 ;
        RECT 2319.5400 739.1400 2321.1400 739.6200 ;
        RECT 2319.5400 744.5800 2321.1400 745.0600 ;
        RECT 2319.5400 750.0200 2321.1400 750.5000 ;
        RECT 2319.5400 728.2600 2321.1400 728.7400 ;
        RECT 2319.5400 733.7000 2321.1400 734.1800 ;
        RECT 2319.5400 711.9400 2321.1400 712.4200 ;
        RECT 2319.5400 717.3800 2321.1400 717.8600 ;
        RECT 2319.5400 722.8200 2321.1400 723.3000 ;
        RECT 2319.5400 701.0600 2321.1400 701.5400 ;
        RECT 2319.5400 706.5000 2321.1400 706.9800 ;
        RECT 2374.2800 684.7400 2375.8800 685.2200 ;
        RECT 2374.2800 690.1800 2375.8800 690.6600 ;
        RECT 2374.2800 695.6200 2375.8800 696.1000 ;
        RECT 2364.5400 684.7400 2366.1400 685.2200 ;
        RECT 2364.5400 690.1800 2366.1400 690.6600 ;
        RECT 2364.5400 695.6200 2366.1400 696.1000 ;
        RECT 2374.2800 673.8600 2375.8800 674.3400 ;
        RECT 2374.2800 679.3000 2375.8800 679.7800 ;
        RECT 2364.5400 673.8600 2366.1400 674.3400 ;
        RECT 2364.5400 679.3000 2366.1400 679.7800 ;
        RECT 2374.2800 657.5400 2375.8800 658.0200 ;
        RECT 2374.2800 662.9800 2375.8800 663.4600 ;
        RECT 2374.2800 668.4200 2375.8800 668.9000 ;
        RECT 2364.5400 657.5400 2366.1400 658.0200 ;
        RECT 2364.5400 662.9800 2366.1400 663.4600 ;
        RECT 2364.5400 668.4200 2366.1400 668.9000 ;
        RECT 2364.5400 652.1000 2366.1400 652.5800 ;
        RECT 2374.2800 652.1000 2375.8800 652.5800 ;
        RECT 2319.5400 684.7400 2321.1400 685.2200 ;
        RECT 2319.5400 690.1800 2321.1400 690.6600 ;
        RECT 2319.5400 695.6200 2321.1400 696.1000 ;
        RECT 2319.5400 673.8600 2321.1400 674.3400 ;
        RECT 2319.5400 679.3000 2321.1400 679.7800 ;
        RECT 2319.5400 657.5400 2321.1400 658.0200 ;
        RECT 2319.5400 662.9800 2321.1400 663.4600 ;
        RECT 2319.5400 668.4200 2321.1400 668.9000 ;
        RECT 2319.5400 652.1000 2321.1400 652.5800 ;
        RECT 2274.5400 739.1400 2276.1400 739.6200 ;
        RECT 2274.5400 744.5800 2276.1400 745.0600 ;
        RECT 2274.5400 750.0200 2276.1400 750.5000 ;
        RECT 2274.5400 728.2600 2276.1400 728.7400 ;
        RECT 2274.5400 733.7000 2276.1400 734.1800 ;
        RECT 2229.5400 739.1400 2231.1400 739.6200 ;
        RECT 2229.5400 744.5800 2231.1400 745.0600 ;
        RECT 2229.5400 750.0200 2231.1400 750.5000 ;
        RECT 2229.5400 728.2600 2231.1400 728.7400 ;
        RECT 2229.5400 733.7000 2231.1400 734.1800 ;
        RECT 2274.5400 711.9400 2276.1400 712.4200 ;
        RECT 2274.5400 717.3800 2276.1400 717.8600 ;
        RECT 2274.5400 722.8200 2276.1400 723.3000 ;
        RECT 2274.5400 701.0600 2276.1400 701.5400 ;
        RECT 2274.5400 706.5000 2276.1400 706.9800 ;
        RECT 2229.5400 711.9400 2231.1400 712.4200 ;
        RECT 2229.5400 717.3800 2231.1400 717.8600 ;
        RECT 2229.5400 722.8200 2231.1400 723.3000 ;
        RECT 2229.5400 701.0600 2231.1400 701.5400 ;
        RECT 2229.5400 706.5000 2231.1400 706.9800 ;
        RECT 2184.5400 739.1400 2186.1400 739.6200 ;
        RECT 2184.5400 744.5800 2186.1400 745.0600 ;
        RECT 2184.5400 750.0200 2186.1400 750.5000 ;
        RECT 2176.7800 739.1400 2178.3800 739.6200 ;
        RECT 2176.7800 744.5800 2178.3800 745.0600 ;
        RECT 2176.7800 750.0200 2178.3800 750.5000 ;
        RECT 2184.5400 728.2600 2186.1400 728.7400 ;
        RECT 2184.5400 733.7000 2186.1400 734.1800 ;
        RECT 2176.7800 728.2600 2178.3800 728.7400 ;
        RECT 2176.7800 733.7000 2178.3800 734.1800 ;
        RECT 2184.5400 711.9400 2186.1400 712.4200 ;
        RECT 2184.5400 717.3800 2186.1400 717.8600 ;
        RECT 2184.5400 722.8200 2186.1400 723.3000 ;
        RECT 2176.7800 711.9400 2178.3800 712.4200 ;
        RECT 2176.7800 717.3800 2178.3800 717.8600 ;
        RECT 2176.7800 722.8200 2178.3800 723.3000 ;
        RECT 2184.5400 701.0600 2186.1400 701.5400 ;
        RECT 2184.5400 706.5000 2186.1400 706.9800 ;
        RECT 2176.7800 701.0600 2178.3800 701.5400 ;
        RECT 2176.7800 706.5000 2178.3800 706.9800 ;
        RECT 2274.5400 684.7400 2276.1400 685.2200 ;
        RECT 2274.5400 690.1800 2276.1400 690.6600 ;
        RECT 2274.5400 695.6200 2276.1400 696.1000 ;
        RECT 2274.5400 673.8600 2276.1400 674.3400 ;
        RECT 2274.5400 679.3000 2276.1400 679.7800 ;
        RECT 2229.5400 684.7400 2231.1400 685.2200 ;
        RECT 2229.5400 690.1800 2231.1400 690.6600 ;
        RECT 2229.5400 695.6200 2231.1400 696.1000 ;
        RECT 2229.5400 673.8600 2231.1400 674.3400 ;
        RECT 2229.5400 679.3000 2231.1400 679.7800 ;
        RECT 2274.5400 657.5400 2276.1400 658.0200 ;
        RECT 2274.5400 662.9800 2276.1400 663.4600 ;
        RECT 2274.5400 668.4200 2276.1400 668.9000 ;
        RECT 2274.5400 652.1000 2276.1400 652.5800 ;
        RECT 2229.5400 657.5400 2231.1400 658.0200 ;
        RECT 2229.5400 662.9800 2231.1400 663.4600 ;
        RECT 2229.5400 668.4200 2231.1400 668.9000 ;
        RECT 2229.5400 652.1000 2231.1400 652.5800 ;
        RECT 2184.5400 684.7400 2186.1400 685.2200 ;
        RECT 2184.5400 690.1800 2186.1400 690.6600 ;
        RECT 2184.5400 695.6200 2186.1400 696.1000 ;
        RECT 2176.7800 684.7400 2178.3800 685.2200 ;
        RECT 2176.7800 690.1800 2178.3800 690.6600 ;
        RECT 2176.7800 695.6200 2178.3800 696.1000 ;
        RECT 2184.5400 673.8600 2186.1400 674.3400 ;
        RECT 2184.5400 679.3000 2186.1400 679.7800 ;
        RECT 2176.7800 673.8600 2178.3800 674.3400 ;
        RECT 2176.7800 679.3000 2178.3800 679.7800 ;
        RECT 2184.5400 657.5400 2186.1400 658.0200 ;
        RECT 2184.5400 662.9800 2186.1400 663.4600 ;
        RECT 2184.5400 668.4200 2186.1400 668.9000 ;
        RECT 2176.7800 657.5400 2178.3800 658.0200 ;
        RECT 2176.7800 662.9800 2178.3800 663.4600 ;
        RECT 2176.7800 668.4200 2178.3800 668.9000 ;
        RECT 2176.7800 652.1000 2178.3800 652.5800 ;
        RECT 2184.5400 652.1000 2186.1400 652.5800 ;
        RECT 2171.2200 854.4100 2381.4400 856.0100 ;
        RECT 2171.2200 647.9100 2381.4400 649.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 642.4800 2178.3800 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 860.5200 2178.3800 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 642.4800 2375.8800 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 860.5200 2375.8800 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 647.9100 2172.8200 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 647.9100 2381.4400 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 854.4100 2172.8200 856.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 854.4100 2381.4400 856.0100 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'LUT4AB'
    PORT
      LAYER met4 ;
        RECT 2364.5400 418.2700 2366.1400 626.3700 ;
        RECT 2319.5400 418.2700 2321.1400 626.3700 ;
        RECT 2274.5400 418.2700 2276.1400 626.3700 ;
        RECT 2229.5400 418.2700 2231.1400 626.3700 ;
        RECT 2184.5400 418.2700 2186.1400 626.3700 ;
        RECT 2374.2800 412.8400 2375.8800 632.4800 ;
        RECT 2176.7800 412.8400 2178.3800 632.4800 ;
      LAYER met3 ;
        RECT 2374.2800 607.4200 2375.8800 607.9000 ;
        RECT 2374.2800 612.8600 2375.8800 613.3400 ;
        RECT 2364.5400 607.4200 2366.1400 607.9000 ;
        RECT 2364.5400 612.8600 2366.1400 613.3400 ;
        RECT 2364.5400 618.3000 2366.1400 618.7800 ;
        RECT 2374.2800 618.3000 2375.8800 618.7800 ;
        RECT 2374.2800 596.5400 2375.8800 597.0200 ;
        RECT 2374.2800 601.9800 2375.8800 602.4600 ;
        RECT 2364.5400 596.5400 2366.1400 597.0200 ;
        RECT 2364.5400 601.9800 2366.1400 602.4600 ;
        RECT 2374.2800 580.2200 2375.8800 580.7000 ;
        RECT 2374.2800 585.6600 2375.8800 586.1400 ;
        RECT 2364.5400 580.2200 2366.1400 580.7000 ;
        RECT 2364.5400 585.6600 2366.1400 586.1400 ;
        RECT 2364.5400 591.1000 2366.1400 591.5800 ;
        RECT 2374.2800 591.1000 2375.8800 591.5800 ;
        RECT 2319.5400 607.4200 2321.1400 607.9000 ;
        RECT 2319.5400 612.8600 2321.1400 613.3400 ;
        RECT 2319.5400 618.3000 2321.1400 618.7800 ;
        RECT 2319.5400 596.5400 2321.1400 597.0200 ;
        RECT 2319.5400 601.9800 2321.1400 602.4600 ;
        RECT 2319.5400 580.2200 2321.1400 580.7000 ;
        RECT 2319.5400 585.6600 2321.1400 586.1400 ;
        RECT 2319.5400 591.1000 2321.1400 591.5800 ;
        RECT 2374.2800 563.9000 2375.8800 564.3800 ;
        RECT 2374.2800 569.3400 2375.8800 569.8200 ;
        RECT 2374.2800 574.7800 2375.8800 575.2600 ;
        RECT 2364.5400 563.9000 2366.1400 564.3800 ;
        RECT 2364.5400 569.3400 2366.1400 569.8200 ;
        RECT 2364.5400 574.7800 2366.1400 575.2600 ;
        RECT 2374.2800 553.0200 2375.8800 553.5000 ;
        RECT 2374.2800 558.4600 2375.8800 558.9400 ;
        RECT 2364.5400 553.0200 2366.1400 553.5000 ;
        RECT 2364.5400 558.4600 2366.1400 558.9400 ;
        RECT 2374.2800 536.7000 2375.8800 537.1800 ;
        RECT 2374.2800 542.1400 2375.8800 542.6200 ;
        RECT 2374.2800 547.5800 2375.8800 548.0600 ;
        RECT 2364.5400 536.7000 2366.1400 537.1800 ;
        RECT 2364.5400 542.1400 2366.1400 542.6200 ;
        RECT 2364.5400 547.5800 2366.1400 548.0600 ;
        RECT 2374.2800 525.8200 2375.8800 526.3000 ;
        RECT 2374.2800 531.2600 2375.8800 531.7400 ;
        RECT 2364.5400 525.8200 2366.1400 526.3000 ;
        RECT 2364.5400 531.2600 2366.1400 531.7400 ;
        RECT 2319.5400 563.9000 2321.1400 564.3800 ;
        RECT 2319.5400 569.3400 2321.1400 569.8200 ;
        RECT 2319.5400 574.7800 2321.1400 575.2600 ;
        RECT 2319.5400 553.0200 2321.1400 553.5000 ;
        RECT 2319.5400 558.4600 2321.1400 558.9400 ;
        RECT 2319.5400 536.7000 2321.1400 537.1800 ;
        RECT 2319.5400 542.1400 2321.1400 542.6200 ;
        RECT 2319.5400 547.5800 2321.1400 548.0600 ;
        RECT 2319.5400 525.8200 2321.1400 526.3000 ;
        RECT 2319.5400 531.2600 2321.1400 531.7400 ;
        RECT 2274.5400 607.4200 2276.1400 607.9000 ;
        RECT 2274.5400 612.8600 2276.1400 613.3400 ;
        RECT 2274.5400 618.3000 2276.1400 618.7800 ;
        RECT 2229.5400 607.4200 2231.1400 607.9000 ;
        RECT 2229.5400 612.8600 2231.1400 613.3400 ;
        RECT 2229.5400 618.3000 2231.1400 618.7800 ;
        RECT 2274.5400 596.5400 2276.1400 597.0200 ;
        RECT 2274.5400 601.9800 2276.1400 602.4600 ;
        RECT 2274.5400 580.2200 2276.1400 580.7000 ;
        RECT 2274.5400 585.6600 2276.1400 586.1400 ;
        RECT 2274.5400 591.1000 2276.1400 591.5800 ;
        RECT 2229.5400 596.5400 2231.1400 597.0200 ;
        RECT 2229.5400 601.9800 2231.1400 602.4600 ;
        RECT 2229.5400 580.2200 2231.1400 580.7000 ;
        RECT 2229.5400 585.6600 2231.1400 586.1400 ;
        RECT 2229.5400 591.1000 2231.1400 591.5800 ;
        RECT 2184.5400 607.4200 2186.1400 607.9000 ;
        RECT 2184.5400 612.8600 2186.1400 613.3400 ;
        RECT 2176.7800 607.4200 2178.3800 607.9000 ;
        RECT 2176.7800 612.8600 2178.3800 613.3400 ;
        RECT 2176.7800 618.3000 2178.3800 618.7800 ;
        RECT 2184.5400 618.3000 2186.1400 618.7800 ;
        RECT 2184.5400 596.5400 2186.1400 597.0200 ;
        RECT 2184.5400 601.9800 2186.1400 602.4600 ;
        RECT 2176.7800 596.5400 2178.3800 597.0200 ;
        RECT 2176.7800 601.9800 2178.3800 602.4600 ;
        RECT 2184.5400 580.2200 2186.1400 580.7000 ;
        RECT 2184.5400 585.6600 2186.1400 586.1400 ;
        RECT 2176.7800 580.2200 2178.3800 580.7000 ;
        RECT 2176.7800 585.6600 2178.3800 586.1400 ;
        RECT 2176.7800 591.1000 2178.3800 591.5800 ;
        RECT 2184.5400 591.1000 2186.1400 591.5800 ;
        RECT 2274.5400 563.9000 2276.1400 564.3800 ;
        RECT 2274.5400 569.3400 2276.1400 569.8200 ;
        RECT 2274.5400 574.7800 2276.1400 575.2600 ;
        RECT 2274.5400 553.0200 2276.1400 553.5000 ;
        RECT 2274.5400 558.4600 2276.1400 558.9400 ;
        RECT 2229.5400 563.9000 2231.1400 564.3800 ;
        RECT 2229.5400 569.3400 2231.1400 569.8200 ;
        RECT 2229.5400 574.7800 2231.1400 575.2600 ;
        RECT 2229.5400 553.0200 2231.1400 553.5000 ;
        RECT 2229.5400 558.4600 2231.1400 558.9400 ;
        RECT 2274.5400 536.7000 2276.1400 537.1800 ;
        RECT 2274.5400 542.1400 2276.1400 542.6200 ;
        RECT 2274.5400 547.5800 2276.1400 548.0600 ;
        RECT 2274.5400 525.8200 2276.1400 526.3000 ;
        RECT 2274.5400 531.2600 2276.1400 531.7400 ;
        RECT 2229.5400 536.7000 2231.1400 537.1800 ;
        RECT 2229.5400 542.1400 2231.1400 542.6200 ;
        RECT 2229.5400 547.5800 2231.1400 548.0600 ;
        RECT 2229.5400 525.8200 2231.1400 526.3000 ;
        RECT 2229.5400 531.2600 2231.1400 531.7400 ;
        RECT 2184.5400 563.9000 2186.1400 564.3800 ;
        RECT 2184.5400 569.3400 2186.1400 569.8200 ;
        RECT 2184.5400 574.7800 2186.1400 575.2600 ;
        RECT 2176.7800 563.9000 2178.3800 564.3800 ;
        RECT 2176.7800 569.3400 2178.3800 569.8200 ;
        RECT 2176.7800 574.7800 2178.3800 575.2600 ;
        RECT 2184.5400 553.0200 2186.1400 553.5000 ;
        RECT 2184.5400 558.4600 2186.1400 558.9400 ;
        RECT 2176.7800 553.0200 2178.3800 553.5000 ;
        RECT 2176.7800 558.4600 2178.3800 558.9400 ;
        RECT 2184.5400 536.7000 2186.1400 537.1800 ;
        RECT 2184.5400 542.1400 2186.1400 542.6200 ;
        RECT 2184.5400 547.5800 2186.1400 548.0600 ;
        RECT 2176.7800 536.7000 2178.3800 537.1800 ;
        RECT 2176.7800 542.1400 2178.3800 542.6200 ;
        RECT 2176.7800 547.5800 2178.3800 548.0600 ;
        RECT 2184.5400 525.8200 2186.1400 526.3000 ;
        RECT 2184.5400 531.2600 2186.1400 531.7400 ;
        RECT 2176.7800 525.8200 2178.3800 526.3000 ;
        RECT 2176.7800 531.2600 2178.3800 531.7400 ;
        RECT 2374.2800 509.5000 2375.8800 509.9800 ;
        RECT 2374.2800 514.9400 2375.8800 515.4200 ;
        RECT 2374.2800 520.3800 2375.8800 520.8600 ;
        RECT 2364.5400 509.5000 2366.1400 509.9800 ;
        RECT 2364.5400 514.9400 2366.1400 515.4200 ;
        RECT 2364.5400 520.3800 2366.1400 520.8600 ;
        RECT 2374.2800 498.6200 2375.8800 499.1000 ;
        RECT 2374.2800 504.0600 2375.8800 504.5400 ;
        RECT 2364.5400 498.6200 2366.1400 499.1000 ;
        RECT 2364.5400 504.0600 2366.1400 504.5400 ;
        RECT 2374.2800 482.3000 2375.8800 482.7800 ;
        RECT 2374.2800 487.7400 2375.8800 488.2200 ;
        RECT 2374.2800 493.1800 2375.8800 493.6600 ;
        RECT 2364.5400 482.3000 2366.1400 482.7800 ;
        RECT 2364.5400 487.7400 2366.1400 488.2200 ;
        RECT 2364.5400 493.1800 2366.1400 493.6600 ;
        RECT 2374.2800 471.4200 2375.8800 471.9000 ;
        RECT 2374.2800 476.8600 2375.8800 477.3400 ;
        RECT 2364.5400 471.4200 2366.1400 471.9000 ;
        RECT 2364.5400 476.8600 2366.1400 477.3400 ;
        RECT 2319.5400 509.5000 2321.1400 509.9800 ;
        RECT 2319.5400 514.9400 2321.1400 515.4200 ;
        RECT 2319.5400 520.3800 2321.1400 520.8600 ;
        RECT 2319.5400 498.6200 2321.1400 499.1000 ;
        RECT 2319.5400 504.0600 2321.1400 504.5400 ;
        RECT 2319.5400 482.3000 2321.1400 482.7800 ;
        RECT 2319.5400 487.7400 2321.1400 488.2200 ;
        RECT 2319.5400 493.1800 2321.1400 493.6600 ;
        RECT 2319.5400 471.4200 2321.1400 471.9000 ;
        RECT 2319.5400 476.8600 2321.1400 477.3400 ;
        RECT 2374.2800 455.1000 2375.8800 455.5800 ;
        RECT 2374.2800 460.5400 2375.8800 461.0200 ;
        RECT 2374.2800 465.9800 2375.8800 466.4600 ;
        RECT 2364.5400 455.1000 2366.1400 455.5800 ;
        RECT 2364.5400 460.5400 2366.1400 461.0200 ;
        RECT 2364.5400 465.9800 2366.1400 466.4600 ;
        RECT 2374.2800 444.2200 2375.8800 444.7000 ;
        RECT 2374.2800 449.6600 2375.8800 450.1400 ;
        RECT 2364.5400 444.2200 2366.1400 444.7000 ;
        RECT 2364.5400 449.6600 2366.1400 450.1400 ;
        RECT 2374.2800 427.9000 2375.8800 428.3800 ;
        RECT 2374.2800 433.3400 2375.8800 433.8200 ;
        RECT 2374.2800 438.7800 2375.8800 439.2600 ;
        RECT 2364.5400 427.9000 2366.1400 428.3800 ;
        RECT 2364.5400 433.3400 2366.1400 433.8200 ;
        RECT 2364.5400 438.7800 2366.1400 439.2600 ;
        RECT 2364.5400 422.4600 2366.1400 422.9400 ;
        RECT 2374.2800 422.4600 2375.8800 422.9400 ;
        RECT 2319.5400 455.1000 2321.1400 455.5800 ;
        RECT 2319.5400 460.5400 2321.1400 461.0200 ;
        RECT 2319.5400 465.9800 2321.1400 466.4600 ;
        RECT 2319.5400 444.2200 2321.1400 444.7000 ;
        RECT 2319.5400 449.6600 2321.1400 450.1400 ;
        RECT 2319.5400 427.9000 2321.1400 428.3800 ;
        RECT 2319.5400 433.3400 2321.1400 433.8200 ;
        RECT 2319.5400 438.7800 2321.1400 439.2600 ;
        RECT 2319.5400 422.4600 2321.1400 422.9400 ;
        RECT 2274.5400 509.5000 2276.1400 509.9800 ;
        RECT 2274.5400 514.9400 2276.1400 515.4200 ;
        RECT 2274.5400 520.3800 2276.1400 520.8600 ;
        RECT 2274.5400 498.6200 2276.1400 499.1000 ;
        RECT 2274.5400 504.0600 2276.1400 504.5400 ;
        RECT 2229.5400 509.5000 2231.1400 509.9800 ;
        RECT 2229.5400 514.9400 2231.1400 515.4200 ;
        RECT 2229.5400 520.3800 2231.1400 520.8600 ;
        RECT 2229.5400 498.6200 2231.1400 499.1000 ;
        RECT 2229.5400 504.0600 2231.1400 504.5400 ;
        RECT 2274.5400 482.3000 2276.1400 482.7800 ;
        RECT 2274.5400 487.7400 2276.1400 488.2200 ;
        RECT 2274.5400 493.1800 2276.1400 493.6600 ;
        RECT 2274.5400 471.4200 2276.1400 471.9000 ;
        RECT 2274.5400 476.8600 2276.1400 477.3400 ;
        RECT 2229.5400 482.3000 2231.1400 482.7800 ;
        RECT 2229.5400 487.7400 2231.1400 488.2200 ;
        RECT 2229.5400 493.1800 2231.1400 493.6600 ;
        RECT 2229.5400 471.4200 2231.1400 471.9000 ;
        RECT 2229.5400 476.8600 2231.1400 477.3400 ;
        RECT 2184.5400 509.5000 2186.1400 509.9800 ;
        RECT 2184.5400 514.9400 2186.1400 515.4200 ;
        RECT 2184.5400 520.3800 2186.1400 520.8600 ;
        RECT 2176.7800 509.5000 2178.3800 509.9800 ;
        RECT 2176.7800 514.9400 2178.3800 515.4200 ;
        RECT 2176.7800 520.3800 2178.3800 520.8600 ;
        RECT 2184.5400 498.6200 2186.1400 499.1000 ;
        RECT 2184.5400 504.0600 2186.1400 504.5400 ;
        RECT 2176.7800 498.6200 2178.3800 499.1000 ;
        RECT 2176.7800 504.0600 2178.3800 504.5400 ;
        RECT 2184.5400 482.3000 2186.1400 482.7800 ;
        RECT 2184.5400 487.7400 2186.1400 488.2200 ;
        RECT 2184.5400 493.1800 2186.1400 493.6600 ;
        RECT 2176.7800 482.3000 2178.3800 482.7800 ;
        RECT 2176.7800 487.7400 2178.3800 488.2200 ;
        RECT 2176.7800 493.1800 2178.3800 493.6600 ;
        RECT 2184.5400 471.4200 2186.1400 471.9000 ;
        RECT 2184.5400 476.8600 2186.1400 477.3400 ;
        RECT 2176.7800 471.4200 2178.3800 471.9000 ;
        RECT 2176.7800 476.8600 2178.3800 477.3400 ;
        RECT 2274.5400 455.1000 2276.1400 455.5800 ;
        RECT 2274.5400 460.5400 2276.1400 461.0200 ;
        RECT 2274.5400 465.9800 2276.1400 466.4600 ;
        RECT 2274.5400 444.2200 2276.1400 444.7000 ;
        RECT 2274.5400 449.6600 2276.1400 450.1400 ;
        RECT 2229.5400 455.1000 2231.1400 455.5800 ;
        RECT 2229.5400 460.5400 2231.1400 461.0200 ;
        RECT 2229.5400 465.9800 2231.1400 466.4600 ;
        RECT 2229.5400 444.2200 2231.1400 444.7000 ;
        RECT 2229.5400 449.6600 2231.1400 450.1400 ;
        RECT 2274.5400 427.9000 2276.1400 428.3800 ;
        RECT 2274.5400 433.3400 2276.1400 433.8200 ;
        RECT 2274.5400 438.7800 2276.1400 439.2600 ;
        RECT 2274.5400 422.4600 2276.1400 422.9400 ;
        RECT 2229.5400 427.9000 2231.1400 428.3800 ;
        RECT 2229.5400 433.3400 2231.1400 433.8200 ;
        RECT 2229.5400 438.7800 2231.1400 439.2600 ;
        RECT 2229.5400 422.4600 2231.1400 422.9400 ;
        RECT 2184.5400 455.1000 2186.1400 455.5800 ;
        RECT 2184.5400 460.5400 2186.1400 461.0200 ;
        RECT 2184.5400 465.9800 2186.1400 466.4600 ;
        RECT 2176.7800 455.1000 2178.3800 455.5800 ;
        RECT 2176.7800 460.5400 2178.3800 461.0200 ;
        RECT 2176.7800 465.9800 2178.3800 466.4600 ;
        RECT 2184.5400 444.2200 2186.1400 444.7000 ;
        RECT 2184.5400 449.6600 2186.1400 450.1400 ;
        RECT 2176.7800 444.2200 2178.3800 444.7000 ;
        RECT 2176.7800 449.6600 2178.3800 450.1400 ;
        RECT 2184.5400 427.9000 2186.1400 428.3800 ;
        RECT 2184.5400 433.3400 2186.1400 433.8200 ;
        RECT 2184.5400 438.7800 2186.1400 439.2600 ;
        RECT 2176.7800 427.9000 2178.3800 428.3800 ;
        RECT 2176.7800 433.3400 2178.3800 433.8200 ;
        RECT 2176.7800 438.7800 2178.3800 439.2600 ;
        RECT 2176.7800 422.4600 2178.3800 422.9400 ;
        RECT 2184.5400 422.4600 2186.1400 422.9400 ;
        RECT 2171.2200 624.7700 2381.4400 626.3700 ;
        RECT 2171.2200 418.2700 2381.4400 419.8700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 412.8400 2178.3800 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2176.7800 630.8800 2178.3800 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 412.8400 2375.8800 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2374.2800 630.8800 2375.8800 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 418.2700 2172.8200 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 418.2700 2381.4400 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2171.2200 624.7700 2172.8200 626.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2379.8400 624.7700 2381.4400 626.3700 ;
    END
# end of P/G pin shape extracted from block 'LUT4AB'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 183.2000 2436.0200 402.8400 ;
        RECT 2397.0000 183.2000 2398.6000 402.8400 ;
      LAYER met3 ;
        RECT 2434.4200 377.7800 2436.0200 378.2600 ;
        RECT 2434.4200 383.2200 2436.0200 383.7000 ;
        RECT 2434.4200 388.6600 2436.0200 389.1400 ;
        RECT 2434.4200 366.9000 2436.0200 367.3800 ;
        RECT 2434.4200 372.3400 2436.0200 372.8200 ;
        RECT 2434.4200 350.5800 2436.0200 351.0600 ;
        RECT 2434.4200 356.0200 2436.0200 356.5000 ;
        RECT 2434.4200 361.4600 2436.0200 361.9400 ;
        RECT 2434.4200 334.2600 2436.0200 334.7400 ;
        RECT 2434.4200 339.7000 2436.0200 340.1800 ;
        RECT 2434.4200 345.1400 2436.0200 345.6200 ;
        RECT 2434.4200 323.3800 2436.0200 323.8600 ;
        RECT 2434.4200 328.8200 2436.0200 329.3000 ;
        RECT 2434.4200 307.0600 2436.0200 307.5400 ;
        RECT 2434.4200 312.5000 2436.0200 312.9800 ;
        RECT 2434.4200 317.9400 2436.0200 318.4200 ;
        RECT 2434.4200 296.1800 2436.0200 296.6600 ;
        RECT 2434.4200 301.6200 2436.0200 302.1000 ;
        RECT 2397.0000 377.7800 2398.6000 378.2600 ;
        RECT 2397.0000 383.2200 2398.6000 383.7000 ;
        RECT 2397.0000 388.6600 2398.6000 389.1400 ;
        RECT 2397.0000 366.9000 2398.6000 367.3800 ;
        RECT 2397.0000 372.3400 2398.6000 372.8200 ;
        RECT 2397.0000 350.5800 2398.6000 351.0600 ;
        RECT 2397.0000 356.0200 2398.6000 356.5000 ;
        RECT 2397.0000 361.4600 2398.6000 361.9400 ;
        RECT 2397.0000 334.2600 2398.6000 334.7400 ;
        RECT 2397.0000 339.7000 2398.6000 340.1800 ;
        RECT 2397.0000 345.1400 2398.6000 345.6200 ;
        RECT 2397.0000 323.3800 2398.6000 323.8600 ;
        RECT 2397.0000 328.8200 2398.6000 329.3000 ;
        RECT 2397.0000 307.0600 2398.6000 307.5400 ;
        RECT 2397.0000 312.5000 2398.6000 312.9800 ;
        RECT 2397.0000 317.9400 2398.6000 318.4200 ;
        RECT 2397.0000 296.1800 2398.6000 296.6600 ;
        RECT 2397.0000 301.6200 2398.6000 302.1000 ;
        RECT 2434.4200 279.8600 2436.0200 280.3400 ;
        RECT 2434.4200 285.3000 2436.0200 285.7800 ;
        RECT 2434.4200 290.7400 2436.0200 291.2200 ;
        RECT 2434.4200 268.9800 2436.0200 269.4600 ;
        RECT 2434.4200 274.4200 2436.0200 274.9000 ;
        RECT 2434.4200 252.6600 2436.0200 253.1400 ;
        RECT 2434.4200 258.1000 2436.0200 258.5800 ;
        RECT 2434.4200 263.5400 2436.0200 264.0200 ;
        RECT 2434.4200 241.7800 2436.0200 242.2600 ;
        RECT 2434.4200 247.2200 2436.0200 247.7000 ;
        RECT 2434.4200 225.4600 2436.0200 225.9400 ;
        RECT 2434.4200 230.9000 2436.0200 231.3800 ;
        RECT 2434.4200 236.3400 2436.0200 236.8200 ;
        RECT 2434.4200 214.5800 2436.0200 215.0600 ;
        RECT 2434.4200 220.0200 2436.0200 220.5000 ;
        RECT 2434.4200 198.2600 2436.0200 198.7400 ;
        RECT 2434.4200 203.7000 2436.0200 204.1800 ;
        RECT 2434.4200 209.1400 2436.0200 209.6200 ;
        RECT 2434.4200 192.8200 2436.0200 193.3000 ;
        RECT 2397.0000 279.8600 2398.6000 280.3400 ;
        RECT 2397.0000 285.3000 2398.6000 285.7800 ;
        RECT 2397.0000 290.7400 2398.6000 291.2200 ;
        RECT 2397.0000 268.9800 2398.6000 269.4600 ;
        RECT 2397.0000 274.4200 2398.6000 274.9000 ;
        RECT 2397.0000 252.6600 2398.6000 253.1400 ;
        RECT 2397.0000 258.1000 2398.6000 258.5800 ;
        RECT 2397.0000 263.5400 2398.6000 264.0200 ;
        RECT 2397.0000 241.7800 2398.6000 242.2600 ;
        RECT 2397.0000 247.2200 2398.6000 247.7000 ;
        RECT 2397.0000 225.4600 2398.6000 225.9400 ;
        RECT 2397.0000 230.9000 2398.6000 231.3800 ;
        RECT 2397.0000 236.3400 2398.6000 236.8200 ;
        RECT 2397.0000 214.5800 2398.6000 215.0600 ;
        RECT 2397.0000 220.0200 2398.6000 220.5000 ;
        RECT 2397.0000 198.2600 2398.6000 198.7400 ;
        RECT 2397.0000 203.7000 2398.6000 204.1800 ;
        RECT 2397.0000 209.1400 2398.6000 209.6200 ;
        RECT 2397.0000 192.8200 2398.6000 193.3000 ;
        RECT 2391.4400 395.1300 2441.5800 396.7300 ;
        RECT 2391.4400 188.6300 2441.5800 190.2300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 183.2000 2398.6000 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 401.2400 2398.6000 402.8400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 183.2000 2436.0200 184.8000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 401.2400 2436.0200 402.8400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 188.6300 2393.0400 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 188.6300 2441.5800 190.2300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 395.1300 2393.0400 396.7300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 395.1300 2441.5800 396.7300 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 2249.9600 2436.0200 2469.6000 ;
        RECT 2397.0000 2249.9600 2398.6000 2469.6000 ;
      LAYER met3 ;
        RECT 2434.4200 2444.5400 2436.0200 2445.0200 ;
        RECT 2434.4200 2449.9800 2436.0200 2450.4600 ;
        RECT 2434.4200 2455.4200 2436.0200 2455.9000 ;
        RECT 2434.4200 2433.6600 2436.0200 2434.1400 ;
        RECT 2434.4200 2439.1000 2436.0200 2439.5800 ;
        RECT 2434.4200 2417.3400 2436.0200 2417.8200 ;
        RECT 2434.4200 2422.7800 2436.0200 2423.2600 ;
        RECT 2434.4200 2428.2200 2436.0200 2428.7000 ;
        RECT 2434.4200 2401.0200 2436.0200 2401.5000 ;
        RECT 2434.4200 2406.4600 2436.0200 2406.9400 ;
        RECT 2434.4200 2411.9000 2436.0200 2412.3800 ;
        RECT 2434.4200 2390.1400 2436.0200 2390.6200 ;
        RECT 2434.4200 2395.5800 2436.0200 2396.0600 ;
        RECT 2434.4200 2373.8200 2436.0200 2374.3000 ;
        RECT 2434.4200 2379.2600 2436.0200 2379.7400 ;
        RECT 2434.4200 2384.7000 2436.0200 2385.1800 ;
        RECT 2434.4200 2362.9400 2436.0200 2363.4200 ;
        RECT 2434.4200 2368.3800 2436.0200 2368.8600 ;
        RECT 2397.0000 2444.5400 2398.6000 2445.0200 ;
        RECT 2397.0000 2449.9800 2398.6000 2450.4600 ;
        RECT 2397.0000 2455.4200 2398.6000 2455.9000 ;
        RECT 2397.0000 2433.6600 2398.6000 2434.1400 ;
        RECT 2397.0000 2439.1000 2398.6000 2439.5800 ;
        RECT 2397.0000 2417.3400 2398.6000 2417.8200 ;
        RECT 2397.0000 2422.7800 2398.6000 2423.2600 ;
        RECT 2397.0000 2428.2200 2398.6000 2428.7000 ;
        RECT 2397.0000 2401.0200 2398.6000 2401.5000 ;
        RECT 2397.0000 2406.4600 2398.6000 2406.9400 ;
        RECT 2397.0000 2411.9000 2398.6000 2412.3800 ;
        RECT 2397.0000 2390.1400 2398.6000 2390.6200 ;
        RECT 2397.0000 2395.5800 2398.6000 2396.0600 ;
        RECT 2397.0000 2373.8200 2398.6000 2374.3000 ;
        RECT 2397.0000 2379.2600 2398.6000 2379.7400 ;
        RECT 2397.0000 2384.7000 2398.6000 2385.1800 ;
        RECT 2397.0000 2362.9400 2398.6000 2363.4200 ;
        RECT 2397.0000 2368.3800 2398.6000 2368.8600 ;
        RECT 2434.4200 2346.6200 2436.0200 2347.1000 ;
        RECT 2434.4200 2352.0600 2436.0200 2352.5400 ;
        RECT 2434.4200 2357.5000 2436.0200 2357.9800 ;
        RECT 2434.4200 2335.7400 2436.0200 2336.2200 ;
        RECT 2434.4200 2341.1800 2436.0200 2341.6600 ;
        RECT 2434.4200 2319.4200 2436.0200 2319.9000 ;
        RECT 2434.4200 2324.8600 2436.0200 2325.3400 ;
        RECT 2434.4200 2330.3000 2436.0200 2330.7800 ;
        RECT 2434.4200 2308.5400 2436.0200 2309.0200 ;
        RECT 2434.4200 2313.9800 2436.0200 2314.4600 ;
        RECT 2434.4200 2292.2200 2436.0200 2292.7000 ;
        RECT 2434.4200 2297.6600 2436.0200 2298.1400 ;
        RECT 2434.4200 2303.1000 2436.0200 2303.5800 ;
        RECT 2434.4200 2281.3400 2436.0200 2281.8200 ;
        RECT 2434.4200 2286.7800 2436.0200 2287.2600 ;
        RECT 2434.4200 2265.0200 2436.0200 2265.5000 ;
        RECT 2434.4200 2270.4600 2436.0200 2270.9400 ;
        RECT 2434.4200 2275.9000 2436.0200 2276.3800 ;
        RECT 2434.4200 2259.5800 2436.0200 2260.0600 ;
        RECT 2397.0000 2346.6200 2398.6000 2347.1000 ;
        RECT 2397.0000 2352.0600 2398.6000 2352.5400 ;
        RECT 2397.0000 2357.5000 2398.6000 2357.9800 ;
        RECT 2397.0000 2335.7400 2398.6000 2336.2200 ;
        RECT 2397.0000 2341.1800 2398.6000 2341.6600 ;
        RECT 2397.0000 2319.4200 2398.6000 2319.9000 ;
        RECT 2397.0000 2324.8600 2398.6000 2325.3400 ;
        RECT 2397.0000 2330.3000 2398.6000 2330.7800 ;
        RECT 2397.0000 2308.5400 2398.6000 2309.0200 ;
        RECT 2397.0000 2313.9800 2398.6000 2314.4600 ;
        RECT 2397.0000 2292.2200 2398.6000 2292.7000 ;
        RECT 2397.0000 2297.6600 2398.6000 2298.1400 ;
        RECT 2397.0000 2303.1000 2398.6000 2303.5800 ;
        RECT 2397.0000 2281.3400 2398.6000 2281.8200 ;
        RECT 2397.0000 2286.7800 2398.6000 2287.2600 ;
        RECT 2397.0000 2265.0200 2398.6000 2265.5000 ;
        RECT 2397.0000 2270.4600 2398.6000 2270.9400 ;
        RECT 2397.0000 2275.9000 2398.6000 2276.3800 ;
        RECT 2397.0000 2259.5800 2398.6000 2260.0600 ;
        RECT 2391.4400 2461.8900 2441.5800 2463.4900 ;
        RECT 2391.4400 2255.3900 2441.5800 2256.9900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 2249.9600 2398.6000 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 2468.0000 2398.6000 2469.6000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 2249.9600 2436.0200 2251.5600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 2468.0000 2436.0200 2469.6000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2255.3900 2393.0400 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2255.3900 2441.5800 2256.9900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2461.8900 2393.0400 2463.4900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2461.8900 2441.5800 2463.4900 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 2020.3200 2436.0200 2239.9600 ;
        RECT 2397.0000 2020.3200 2398.6000 2239.9600 ;
      LAYER met3 ;
        RECT 2434.4200 2214.9000 2436.0200 2215.3800 ;
        RECT 2434.4200 2220.3400 2436.0200 2220.8200 ;
        RECT 2434.4200 2225.7800 2436.0200 2226.2600 ;
        RECT 2434.4200 2204.0200 2436.0200 2204.5000 ;
        RECT 2434.4200 2209.4600 2436.0200 2209.9400 ;
        RECT 2434.4200 2187.7000 2436.0200 2188.1800 ;
        RECT 2434.4200 2193.1400 2436.0200 2193.6200 ;
        RECT 2434.4200 2198.5800 2436.0200 2199.0600 ;
        RECT 2434.4200 2171.3800 2436.0200 2171.8600 ;
        RECT 2434.4200 2176.8200 2436.0200 2177.3000 ;
        RECT 2434.4200 2182.2600 2436.0200 2182.7400 ;
        RECT 2434.4200 2160.5000 2436.0200 2160.9800 ;
        RECT 2434.4200 2165.9400 2436.0200 2166.4200 ;
        RECT 2434.4200 2144.1800 2436.0200 2144.6600 ;
        RECT 2434.4200 2149.6200 2436.0200 2150.1000 ;
        RECT 2434.4200 2155.0600 2436.0200 2155.5400 ;
        RECT 2434.4200 2133.3000 2436.0200 2133.7800 ;
        RECT 2434.4200 2138.7400 2436.0200 2139.2200 ;
        RECT 2397.0000 2214.9000 2398.6000 2215.3800 ;
        RECT 2397.0000 2220.3400 2398.6000 2220.8200 ;
        RECT 2397.0000 2225.7800 2398.6000 2226.2600 ;
        RECT 2397.0000 2204.0200 2398.6000 2204.5000 ;
        RECT 2397.0000 2209.4600 2398.6000 2209.9400 ;
        RECT 2397.0000 2187.7000 2398.6000 2188.1800 ;
        RECT 2397.0000 2193.1400 2398.6000 2193.6200 ;
        RECT 2397.0000 2198.5800 2398.6000 2199.0600 ;
        RECT 2397.0000 2171.3800 2398.6000 2171.8600 ;
        RECT 2397.0000 2176.8200 2398.6000 2177.3000 ;
        RECT 2397.0000 2182.2600 2398.6000 2182.7400 ;
        RECT 2397.0000 2160.5000 2398.6000 2160.9800 ;
        RECT 2397.0000 2165.9400 2398.6000 2166.4200 ;
        RECT 2397.0000 2144.1800 2398.6000 2144.6600 ;
        RECT 2397.0000 2149.6200 2398.6000 2150.1000 ;
        RECT 2397.0000 2155.0600 2398.6000 2155.5400 ;
        RECT 2397.0000 2133.3000 2398.6000 2133.7800 ;
        RECT 2397.0000 2138.7400 2398.6000 2139.2200 ;
        RECT 2434.4200 2116.9800 2436.0200 2117.4600 ;
        RECT 2434.4200 2122.4200 2436.0200 2122.9000 ;
        RECT 2434.4200 2127.8600 2436.0200 2128.3400 ;
        RECT 2434.4200 2106.1000 2436.0200 2106.5800 ;
        RECT 2434.4200 2111.5400 2436.0200 2112.0200 ;
        RECT 2434.4200 2089.7800 2436.0200 2090.2600 ;
        RECT 2434.4200 2095.2200 2436.0200 2095.7000 ;
        RECT 2434.4200 2100.6600 2436.0200 2101.1400 ;
        RECT 2434.4200 2078.9000 2436.0200 2079.3800 ;
        RECT 2434.4200 2084.3400 2436.0200 2084.8200 ;
        RECT 2434.4200 2062.5800 2436.0200 2063.0600 ;
        RECT 2434.4200 2068.0200 2436.0200 2068.5000 ;
        RECT 2434.4200 2073.4600 2436.0200 2073.9400 ;
        RECT 2434.4200 2051.7000 2436.0200 2052.1800 ;
        RECT 2434.4200 2057.1400 2436.0200 2057.6200 ;
        RECT 2434.4200 2035.3800 2436.0200 2035.8600 ;
        RECT 2434.4200 2040.8200 2436.0200 2041.3000 ;
        RECT 2434.4200 2046.2600 2436.0200 2046.7400 ;
        RECT 2434.4200 2029.9400 2436.0200 2030.4200 ;
        RECT 2397.0000 2116.9800 2398.6000 2117.4600 ;
        RECT 2397.0000 2122.4200 2398.6000 2122.9000 ;
        RECT 2397.0000 2127.8600 2398.6000 2128.3400 ;
        RECT 2397.0000 2106.1000 2398.6000 2106.5800 ;
        RECT 2397.0000 2111.5400 2398.6000 2112.0200 ;
        RECT 2397.0000 2089.7800 2398.6000 2090.2600 ;
        RECT 2397.0000 2095.2200 2398.6000 2095.7000 ;
        RECT 2397.0000 2100.6600 2398.6000 2101.1400 ;
        RECT 2397.0000 2078.9000 2398.6000 2079.3800 ;
        RECT 2397.0000 2084.3400 2398.6000 2084.8200 ;
        RECT 2397.0000 2062.5800 2398.6000 2063.0600 ;
        RECT 2397.0000 2068.0200 2398.6000 2068.5000 ;
        RECT 2397.0000 2073.4600 2398.6000 2073.9400 ;
        RECT 2397.0000 2051.7000 2398.6000 2052.1800 ;
        RECT 2397.0000 2057.1400 2398.6000 2057.6200 ;
        RECT 2397.0000 2035.3800 2398.6000 2035.8600 ;
        RECT 2397.0000 2040.8200 2398.6000 2041.3000 ;
        RECT 2397.0000 2046.2600 2398.6000 2046.7400 ;
        RECT 2397.0000 2029.9400 2398.6000 2030.4200 ;
        RECT 2391.4400 2232.2500 2441.5800 2233.8500 ;
        RECT 2391.4400 2025.7500 2441.5800 2027.3500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 2020.3200 2398.6000 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 2238.3600 2398.6000 2239.9600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 2020.3200 2436.0200 2021.9200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 2238.3600 2436.0200 2239.9600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2025.7500 2393.0400 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2025.7500 2441.5800 2027.3500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2232.2500 2393.0400 2233.8500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2232.2500 2441.5800 2233.8500 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 1790.6800 2436.0200 2010.3200 ;
        RECT 2397.0000 1790.6800 2398.6000 2010.3200 ;
      LAYER met3 ;
        RECT 2434.4200 1985.2600 2436.0200 1985.7400 ;
        RECT 2434.4200 1990.7000 2436.0200 1991.1800 ;
        RECT 2434.4200 1996.1400 2436.0200 1996.6200 ;
        RECT 2434.4200 1974.3800 2436.0200 1974.8600 ;
        RECT 2434.4200 1979.8200 2436.0200 1980.3000 ;
        RECT 2434.4200 1958.0600 2436.0200 1958.5400 ;
        RECT 2434.4200 1963.5000 2436.0200 1963.9800 ;
        RECT 2434.4200 1968.9400 2436.0200 1969.4200 ;
        RECT 2434.4200 1941.7400 2436.0200 1942.2200 ;
        RECT 2434.4200 1947.1800 2436.0200 1947.6600 ;
        RECT 2434.4200 1952.6200 2436.0200 1953.1000 ;
        RECT 2434.4200 1930.8600 2436.0200 1931.3400 ;
        RECT 2434.4200 1936.3000 2436.0200 1936.7800 ;
        RECT 2434.4200 1914.5400 2436.0200 1915.0200 ;
        RECT 2434.4200 1919.9800 2436.0200 1920.4600 ;
        RECT 2434.4200 1925.4200 2436.0200 1925.9000 ;
        RECT 2434.4200 1903.6600 2436.0200 1904.1400 ;
        RECT 2434.4200 1909.1000 2436.0200 1909.5800 ;
        RECT 2397.0000 1985.2600 2398.6000 1985.7400 ;
        RECT 2397.0000 1990.7000 2398.6000 1991.1800 ;
        RECT 2397.0000 1996.1400 2398.6000 1996.6200 ;
        RECT 2397.0000 1974.3800 2398.6000 1974.8600 ;
        RECT 2397.0000 1979.8200 2398.6000 1980.3000 ;
        RECT 2397.0000 1958.0600 2398.6000 1958.5400 ;
        RECT 2397.0000 1963.5000 2398.6000 1963.9800 ;
        RECT 2397.0000 1968.9400 2398.6000 1969.4200 ;
        RECT 2397.0000 1941.7400 2398.6000 1942.2200 ;
        RECT 2397.0000 1947.1800 2398.6000 1947.6600 ;
        RECT 2397.0000 1952.6200 2398.6000 1953.1000 ;
        RECT 2397.0000 1930.8600 2398.6000 1931.3400 ;
        RECT 2397.0000 1936.3000 2398.6000 1936.7800 ;
        RECT 2397.0000 1914.5400 2398.6000 1915.0200 ;
        RECT 2397.0000 1919.9800 2398.6000 1920.4600 ;
        RECT 2397.0000 1925.4200 2398.6000 1925.9000 ;
        RECT 2397.0000 1903.6600 2398.6000 1904.1400 ;
        RECT 2397.0000 1909.1000 2398.6000 1909.5800 ;
        RECT 2434.4200 1887.3400 2436.0200 1887.8200 ;
        RECT 2434.4200 1892.7800 2436.0200 1893.2600 ;
        RECT 2434.4200 1898.2200 2436.0200 1898.7000 ;
        RECT 2434.4200 1876.4600 2436.0200 1876.9400 ;
        RECT 2434.4200 1881.9000 2436.0200 1882.3800 ;
        RECT 2434.4200 1860.1400 2436.0200 1860.6200 ;
        RECT 2434.4200 1865.5800 2436.0200 1866.0600 ;
        RECT 2434.4200 1871.0200 2436.0200 1871.5000 ;
        RECT 2434.4200 1849.2600 2436.0200 1849.7400 ;
        RECT 2434.4200 1854.7000 2436.0200 1855.1800 ;
        RECT 2434.4200 1832.9400 2436.0200 1833.4200 ;
        RECT 2434.4200 1838.3800 2436.0200 1838.8600 ;
        RECT 2434.4200 1843.8200 2436.0200 1844.3000 ;
        RECT 2434.4200 1822.0600 2436.0200 1822.5400 ;
        RECT 2434.4200 1827.5000 2436.0200 1827.9800 ;
        RECT 2434.4200 1805.7400 2436.0200 1806.2200 ;
        RECT 2434.4200 1811.1800 2436.0200 1811.6600 ;
        RECT 2434.4200 1816.6200 2436.0200 1817.1000 ;
        RECT 2434.4200 1800.3000 2436.0200 1800.7800 ;
        RECT 2397.0000 1887.3400 2398.6000 1887.8200 ;
        RECT 2397.0000 1892.7800 2398.6000 1893.2600 ;
        RECT 2397.0000 1898.2200 2398.6000 1898.7000 ;
        RECT 2397.0000 1876.4600 2398.6000 1876.9400 ;
        RECT 2397.0000 1881.9000 2398.6000 1882.3800 ;
        RECT 2397.0000 1860.1400 2398.6000 1860.6200 ;
        RECT 2397.0000 1865.5800 2398.6000 1866.0600 ;
        RECT 2397.0000 1871.0200 2398.6000 1871.5000 ;
        RECT 2397.0000 1849.2600 2398.6000 1849.7400 ;
        RECT 2397.0000 1854.7000 2398.6000 1855.1800 ;
        RECT 2397.0000 1832.9400 2398.6000 1833.4200 ;
        RECT 2397.0000 1838.3800 2398.6000 1838.8600 ;
        RECT 2397.0000 1843.8200 2398.6000 1844.3000 ;
        RECT 2397.0000 1822.0600 2398.6000 1822.5400 ;
        RECT 2397.0000 1827.5000 2398.6000 1827.9800 ;
        RECT 2397.0000 1805.7400 2398.6000 1806.2200 ;
        RECT 2397.0000 1811.1800 2398.6000 1811.6600 ;
        RECT 2397.0000 1816.6200 2398.6000 1817.1000 ;
        RECT 2397.0000 1800.3000 2398.6000 1800.7800 ;
        RECT 2391.4400 2002.6100 2441.5800 2004.2100 ;
        RECT 2391.4400 1796.1100 2441.5800 1797.7100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1790.6800 2398.6000 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 2008.7200 2398.6000 2010.3200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1790.6800 2436.0200 1792.2800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 2008.7200 2436.0200 2010.3200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1796.1100 2393.0400 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1796.1100 2441.5800 1797.7100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 2002.6100 2393.0400 2004.2100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 2002.6100 2441.5800 2004.2100 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 1561.0400 2436.0200 1780.6800 ;
        RECT 2397.0000 1561.0400 2398.6000 1780.6800 ;
      LAYER met3 ;
        RECT 2434.4200 1755.6200 2436.0200 1756.1000 ;
        RECT 2434.4200 1761.0600 2436.0200 1761.5400 ;
        RECT 2434.4200 1766.5000 2436.0200 1766.9800 ;
        RECT 2434.4200 1744.7400 2436.0200 1745.2200 ;
        RECT 2434.4200 1750.1800 2436.0200 1750.6600 ;
        RECT 2434.4200 1728.4200 2436.0200 1728.9000 ;
        RECT 2434.4200 1733.8600 2436.0200 1734.3400 ;
        RECT 2434.4200 1739.3000 2436.0200 1739.7800 ;
        RECT 2434.4200 1712.1000 2436.0200 1712.5800 ;
        RECT 2434.4200 1717.5400 2436.0200 1718.0200 ;
        RECT 2434.4200 1722.9800 2436.0200 1723.4600 ;
        RECT 2434.4200 1701.2200 2436.0200 1701.7000 ;
        RECT 2434.4200 1706.6600 2436.0200 1707.1400 ;
        RECT 2434.4200 1684.9000 2436.0200 1685.3800 ;
        RECT 2434.4200 1690.3400 2436.0200 1690.8200 ;
        RECT 2434.4200 1695.7800 2436.0200 1696.2600 ;
        RECT 2434.4200 1674.0200 2436.0200 1674.5000 ;
        RECT 2434.4200 1679.4600 2436.0200 1679.9400 ;
        RECT 2397.0000 1755.6200 2398.6000 1756.1000 ;
        RECT 2397.0000 1761.0600 2398.6000 1761.5400 ;
        RECT 2397.0000 1766.5000 2398.6000 1766.9800 ;
        RECT 2397.0000 1744.7400 2398.6000 1745.2200 ;
        RECT 2397.0000 1750.1800 2398.6000 1750.6600 ;
        RECT 2397.0000 1728.4200 2398.6000 1728.9000 ;
        RECT 2397.0000 1733.8600 2398.6000 1734.3400 ;
        RECT 2397.0000 1739.3000 2398.6000 1739.7800 ;
        RECT 2397.0000 1712.1000 2398.6000 1712.5800 ;
        RECT 2397.0000 1717.5400 2398.6000 1718.0200 ;
        RECT 2397.0000 1722.9800 2398.6000 1723.4600 ;
        RECT 2397.0000 1701.2200 2398.6000 1701.7000 ;
        RECT 2397.0000 1706.6600 2398.6000 1707.1400 ;
        RECT 2397.0000 1684.9000 2398.6000 1685.3800 ;
        RECT 2397.0000 1690.3400 2398.6000 1690.8200 ;
        RECT 2397.0000 1695.7800 2398.6000 1696.2600 ;
        RECT 2397.0000 1674.0200 2398.6000 1674.5000 ;
        RECT 2397.0000 1679.4600 2398.6000 1679.9400 ;
        RECT 2434.4200 1657.7000 2436.0200 1658.1800 ;
        RECT 2434.4200 1663.1400 2436.0200 1663.6200 ;
        RECT 2434.4200 1668.5800 2436.0200 1669.0600 ;
        RECT 2434.4200 1646.8200 2436.0200 1647.3000 ;
        RECT 2434.4200 1652.2600 2436.0200 1652.7400 ;
        RECT 2434.4200 1630.5000 2436.0200 1630.9800 ;
        RECT 2434.4200 1635.9400 2436.0200 1636.4200 ;
        RECT 2434.4200 1641.3800 2436.0200 1641.8600 ;
        RECT 2434.4200 1619.6200 2436.0200 1620.1000 ;
        RECT 2434.4200 1625.0600 2436.0200 1625.5400 ;
        RECT 2434.4200 1603.3000 2436.0200 1603.7800 ;
        RECT 2434.4200 1608.7400 2436.0200 1609.2200 ;
        RECT 2434.4200 1614.1800 2436.0200 1614.6600 ;
        RECT 2434.4200 1592.4200 2436.0200 1592.9000 ;
        RECT 2434.4200 1597.8600 2436.0200 1598.3400 ;
        RECT 2434.4200 1576.1000 2436.0200 1576.5800 ;
        RECT 2434.4200 1581.5400 2436.0200 1582.0200 ;
        RECT 2434.4200 1586.9800 2436.0200 1587.4600 ;
        RECT 2434.4200 1570.6600 2436.0200 1571.1400 ;
        RECT 2397.0000 1657.7000 2398.6000 1658.1800 ;
        RECT 2397.0000 1663.1400 2398.6000 1663.6200 ;
        RECT 2397.0000 1668.5800 2398.6000 1669.0600 ;
        RECT 2397.0000 1646.8200 2398.6000 1647.3000 ;
        RECT 2397.0000 1652.2600 2398.6000 1652.7400 ;
        RECT 2397.0000 1630.5000 2398.6000 1630.9800 ;
        RECT 2397.0000 1635.9400 2398.6000 1636.4200 ;
        RECT 2397.0000 1641.3800 2398.6000 1641.8600 ;
        RECT 2397.0000 1619.6200 2398.6000 1620.1000 ;
        RECT 2397.0000 1625.0600 2398.6000 1625.5400 ;
        RECT 2397.0000 1603.3000 2398.6000 1603.7800 ;
        RECT 2397.0000 1608.7400 2398.6000 1609.2200 ;
        RECT 2397.0000 1614.1800 2398.6000 1614.6600 ;
        RECT 2397.0000 1592.4200 2398.6000 1592.9000 ;
        RECT 2397.0000 1597.8600 2398.6000 1598.3400 ;
        RECT 2397.0000 1576.1000 2398.6000 1576.5800 ;
        RECT 2397.0000 1581.5400 2398.6000 1582.0200 ;
        RECT 2397.0000 1586.9800 2398.6000 1587.4600 ;
        RECT 2397.0000 1570.6600 2398.6000 1571.1400 ;
        RECT 2391.4400 1772.9700 2441.5800 1774.5700 ;
        RECT 2391.4400 1566.4700 2441.5800 1568.0700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1561.0400 2398.6000 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1779.0800 2398.6000 1780.6800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1561.0400 2436.0200 1562.6400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1779.0800 2436.0200 1780.6800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1566.4700 2393.0400 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1566.4700 2441.5800 1568.0700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1772.9700 2393.0400 1774.5700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1772.9700 2441.5800 1774.5700 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 1331.4000 2436.0200 1551.0400 ;
        RECT 2397.0000 1331.4000 2398.6000 1551.0400 ;
      LAYER met3 ;
        RECT 2434.4200 1525.9800 2436.0200 1526.4600 ;
        RECT 2434.4200 1531.4200 2436.0200 1531.9000 ;
        RECT 2434.4200 1536.8600 2436.0200 1537.3400 ;
        RECT 2434.4200 1515.1000 2436.0200 1515.5800 ;
        RECT 2434.4200 1520.5400 2436.0200 1521.0200 ;
        RECT 2434.4200 1498.7800 2436.0200 1499.2600 ;
        RECT 2434.4200 1504.2200 2436.0200 1504.7000 ;
        RECT 2434.4200 1509.6600 2436.0200 1510.1400 ;
        RECT 2434.4200 1482.4600 2436.0200 1482.9400 ;
        RECT 2434.4200 1487.9000 2436.0200 1488.3800 ;
        RECT 2434.4200 1493.3400 2436.0200 1493.8200 ;
        RECT 2434.4200 1471.5800 2436.0200 1472.0600 ;
        RECT 2434.4200 1477.0200 2436.0200 1477.5000 ;
        RECT 2434.4200 1455.2600 2436.0200 1455.7400 ;
        RECT 2434.4200 1460.7000 2436.0200 1461.1800 ;
        RECT 2434.4200 1466.1400 2436.0200 1466.6200 ;
        RECT 2434.4200 1444.3800 2436.0200 1444.8600 ;
        RECT 2434.4200 1449.8200 2436.0200 1450.3000 ;
        RECT 2397.0000 1525.9800 2398.6000 1526.4600 ;
        RECT 2397.0000 1531.4200 2398.6000 1531.9000 ;
        RECT 2397.0000 1536.8600 2398.6000 1537.3400 ;
        RECT 2397.0000 1515.1000 2398.6000 1515.5800 ;
        RECT 2397.0000 1520.5400 2398.6000 1521.0200 ;
        RECT 2397.0000 1498.7800 2398.6000 1499.2600 ;
        RECT 2397.0000 1504.2200 2398.6000 1504.7000 ;
        RECT 2397.0000 1509.6600 2398.6000 1510.1400 ;
        RECT 2397.0000 1482.4600 2398.6000 1482.9400 ;
        RECT 2397.0000 1487.9000 2398.6000 1488.3800 ;
        RECT 2397.0000 1493.3400 2398.6000 1493.8200 ;
        RECT 2397.0000 1471.5800 2398.6000 1472.0600 ;
        RECT 2397.0000 1477.0200 2398.6000 1477.5000 ;
        RECT 2397.0000 1455.2600 2398.6000 1455.7400 ;
        RECT 2397.0000 1460.7000 2398.6000 1461.1800 ;
        RECT 2397.0000 1466.1400 2398.6000 1466.6200 ;
        RECT 2397.0000 1444.3800 2398.6000 1444.8600 ;
        RECT 2397.0000 1449.8200 2398.6000 1450.3000 ;
        RECT 2434.4200 1428.0600 2436.0200 1428.5400 ;
        RECT 2434.4200 1433.5000 2436.0200 1433.9800 ;
        RECT 2434.4200 1438.9400 2436.0200 1439.4200 ;
        RECT 2434.4200 1417.1800 2436.0200 1417.6600 ;
        RECT 2434.4200 1422.6200 2436.0200 1423.1000 ;
        RECT 2434.4200 1400.8600 2436.0200 1401.3400 ;
        RECT 2434.4200 1406.3000 2436.0200 1406.7800 ;
        RECT 2434.4200 1411.7400 2436.0200 1412.2200 ;
        RECT 2434.4200 1389.9800 2436.0200 1390.4600 ;
        RECT 2434.4200 1395.4200 2436.0200 1395.9000 ;
        RECT 2434.4200 1373.6600 2436.0200 1374.1400 ;
        RECT 2434.4200 1379.1000 2436.0200 1379.5800 ;
        RECT 2434.4200 1384.5400 2436.0200 1385.0200 ;
        RECT 2434.4200 1362.7800 2436.0200 1363.2600 ;
        RECT 2434.4200 1368.2200 2436.0200 1368.7000 ;
        RECT 2434.4200 1346.4600 2436.0200 1346.9400 ;
        RECT 2434.4200 1351.9000 2436.0200 1352.3800 ;
        RECT 2434.4200 1357.3400 2436.0200 1357.8200 ;
        RECT 2434.4200 1341.0200 2436.0200 1341.5000 ;
        RECT 2397.0000 1428.0600 2398.6000 1428.5400 ;
        RECT 2397.0000 1433.5000 2398.6000 1433.9800 ;
        RECT 2397.0000 1438.9400 2398.6000 1439.4200 ;
        RECT 2397.0000 1417.1800 2398.6000 1417.6600 ;
        RECT 2397.0000 1422.6200 2398.6000 1423.1000 ;
        RECT 2397.0000 1400.8600 2398.6000 1401.3400 ;
        RECT 2397.0000 1406.3000 2398.6000 1406.7800 ;
        RECT 2397.0000 1411.7400 2398.6000 1412.2200 ;
        RECT 2397.0000 1389.9800 2398.6000 1390.4600 ;
        RECT 2397.0000 1395.4200 2398.6000 1395.9000 ;
        RECT 2397.0000 1373.6600 2398.6000 1374.1400 ;
        RECT 2397.0000 1379.1000 2398.6000 1379.5800 ;
        RECT 2397.0000 1384.5400 2398.6000 1385.0200 ;
        RECT 2397.0000 1362.7800 2398.6000 1363.2600 ;
        RECT 2397.0000 1368.2200 2398.6000 1368.7000 ;
        RECT 2397.0000 1346.4600 2398.6000 1346.9400 ;
        RECT 2397.0000 1351.9000 2398.6000 1352.3800 ;
        RECT 2397.0000 1357.3400 2398.6000 1357.8200 ;
        RECT 2397.0000 1341.0200 2398.6000 1341.5000 ;
        RECT 2391.4400 1543.3300 2441.5800 1544.9300 ;
        RECT 2391.4400 1336.8300 2441.5800 1338.4300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1331.4000 2398.6000 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1549.4400 2398.6000 1551.0400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1331.4000 2436.0200 1333.0000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1549.4400 2436.0200 1551.0400 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1336.8300 2393.0400 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1336.8300 2441.5800 1338.4300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1543.3300 2393.0400 1544.9300 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1543.3300 2441.5800 1544.9300 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 1101.7600 2436.0200 1321.4000 ;
        RECT 2397.0000 1101.7600 2398.6000 1321.4000 ;
      LAYER met3 ;
        RECT 2434.4200 1296.3400 2436.0200 1296.8200 ;
        RECT 2434.4200 1301.7800 2436.0200 1302.2600 ;
        RECT 2434.4200 1307.2200 2436.0200 1307.7000 ;
        RECT 2434.4200 1285.4600 2436.0200 1285.9400 ;
        RECT 2434.4200 1290.9000 2436.0200 1291.3800 ;
        RECT 2434.4200 1269.1400 2436.0200 1269.6200 ;
        RECT 2434.4200 1274.5800 2436.0200 1275.0600 ;
        RECT 2434.4200 1280.0200 2436.0200 1280.5000 ;
        RECT 2434.4200 1252.8200 2436.0200 1253.3000 ;
        RECT 2434.4200 1258.2600 2436.0200 1258.7400 ;
        RECT 2434.4200 1263.7000 2436.0200 1264.1800 ;
        RECT 2434.4200 1241.9400 2436.0200 1242.4200 ;
        RECT 2434.4200 1247.3800 2436.0200 1247.8600 ;
        RECT 2434.4200 1225.6200 2436.0200 1226.1000 ;
        RECT 2434.4200 1231.0600 2436.0200 1231.5400 ;
        RECT 2434.4200 1236.5000 2436.0200 1236.9800 ;
        RECT 2434.4200 1214.7400 2436.0200 1215.2200 ;
        RECT 2434.4200 1220.1800 2436.0200 1220.6600 ;
        RECT 2397.0000 1296.3400 2398.6000 1296.8200 ;
        RECT 2397.0000 1301.7800 2398.6000 1302.2600 ;
        RECT 2397.0000 1307.2200 2398.6000 1307.7000 ;
        RECT 2397.0000 1285.4600 2398.6000 1285.9400 ;
        RECT 2397.0000 1290.9000 2398.6000 1291.3800 ;
        RECT 2397.0000 1269.1400 2398.6000 1269.6200 ;
        RECT 2397.0000 1274.5800 2398.6000 1275.0600 ;
        RECT 2397.0000 1280.0200 2398.6000 1280.5000 ;
        RECT 2397.0000 1252.8200 2398.6000 1253.3000 ;
        RECT 2397.0000 1258.2600 2398.6000 1258.7400 ;
        RECT 2397.0000 1263.7000 2398.6000 1264.1800 ;
        RECT 2397.0000 1241.9400 2398.6000 1242.4200 ;
        RECT 2397.0000 1247.3800 2398.6000 1247.8600 ;
        RECT 2397.0000 1225.6200 2398.6000 1226.1000 ;
        RECT 2397.0000 1231.0600 2398.6000 1231.5400 ;
        RECT 2397.0000 1236.5000 2398.6000 1236.9800 ;
        RECT 2397.0000 1214.7400 2398.6000 1215.2200 ;
        RECT 2397.0000 1220.1800 2398.6000 1220.6600 ;
        RECT 2434.4200 1198.4200 2436.0200 1198.9000 ;
        RECT 2434.4200 1203.8600 2436.0200 1204.3400 ;
        RECT 2434.4200 1209.3000 2436.0200 1209.7800 ;
        RECT 2434.4200 1187.5400 2436.0200 1188.0200 ;
        RECT 2434.4200 1192.9800 2436.0200 1193.4600 ;
        RECT 2434.4200 1171.2200 2436.0200 1171.7000 ;
        RECT 2434.4200 1176.6600 2436.0200 1177.1400 ;
        RECT 2434.4200 1182.1000 2436.0200 1182.5800 ;
        RECT 2434.4200 1160.3400 2436.0200 1160.8200 ;
        RECT 2434.4200 1165.7800 2436.0200 1166.2600 ;
        RECT 2434.4200 1144.0200 2436.0200 1144.5000 ;
        RECT 2434.4200 1149.4600 2436.0200 1149.9400 ;
        RECT 2434.4200 1154.9000 2436.0200 1155.3800 ;
        RECT 2434.4200 1133.1400 2436.0200 1133.6200 ;
        RECT 2434.4200 1138.5800 2436.0200 1139.0600 ;
        RECT 2434.4200 1116.8200 2436.0200 1117.3000 ;
        RECT 2434.4200 1122.2600 2436.0200 1122.7400 ;
        RECT 2434.4200 1127.7000 2436.0200 1128.1800 ;
        RECT 2434.4200 1111.3800 2436.0200 1111.8600 ;
        RECT 2397.0000 1198.4200 2398.6000 1198.9000 ;
        RECT 2397.0000 1203.8600 2398.6000 1204.3400 ;
        RECT 2397.0000 1209.3000 2398.6000 1209.7800 ;
        RECT 2397.0000 1187.5400 2398.6000 1188.0200 ;
        RECT 2397.0000 1192.9800 2398.6000 1193.4600 ;
        RECT 2397.0000 1171.2200 2398.6000 1171.7000 ;
        RECT 2397.0000 1176.6600 2398.6000 1177.1400 ;
        RECT 2397.0000 1182.1000 2398.6000 1182.5800 ;
        RECT 2397.0000 1160.3400 2398.6000 1160.8200 ;
        RECT 2397.0000 1165.7800 2398.6000 1166.2600 ;
        RECT 2397.0000 1144.0200 2398.6000 1144.5000 ;
        RECT 2397.0000 1149.4600 2398.6000 1149.9400 ;
        RECT 2397.0000 1154.9000 2398.6000 1155.3800 ;
        RECT 2397.0000 1133.1400 2398.6000 1133.6200 ;
        RECT 2397.0000 1138.5800 2398.6000 1139.0600 ;
        RECT 2397.0000 1116.8200 2398.6000 1117.3000 ;
        RECT 2397.0000 1122.2600 2398.6000 1122.7400 ;
        RECT 2397.0000 1127.7000 2398.6000 1128.1800 ;
        RECT 2397.0000 1111.3800 2398.6000 1111.8600 ;
        RECT 2391.4400 1313.6900 2441.5800 1315.2900 ;
        RECT 2391.4400 1107.1900 2441.5800 1108.7900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1101.7600 2398.6000 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1319.8000 2398.6000 1321.4000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1101.7600 2436.0200 1103.3600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1319.8000 2436.0200 1321.4000 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1107.1900 2393.0400 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1107.1900 2441.5800 1108.7900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1313.6900 2393.0400 1315.2900 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1313.6900 2441.5800 1315.2900 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 872.1200 2436.0200 1091.7600 ;
        RECT 2397.0000 872.1200 2398.6000 1091.7600 ;
      LAYER met3 ;
        RECT 2434.4200 1066.7000 2436.0200 1067.1800 ;
        RECT 2434.4200 1072.1400 2436.0200 1072.6200 ;
        RECT 2434.4200 1077.5800 2436.0200 1078.0600 ;
        RECT 2434.4200 1055.8200 2436.0200 1056.3000 ;
        RECT 2434.4200 1061.2600 2436.0200 1061.7400 ;
        RECT 2434.4200 1039.5000 2436.0200 1039.9800 ;
        RECT 2434.4200 1044.9400 2436.0200 1045.4200 ;
        RECT 2434.4200 1050.3800 2436.0200 1050.8600 ;
        RECT 2434.4200 1023.1800 2436.0200 1023.6600 ;
        RECT 2434.4200 1028.6200 2436.0200 1029.1000 ;
        RECT 2434.4200 1034.0600 2436.0200 1034.5400 ;
        RECT 2434.4200 1012.3000 2436.0200 1012.7800 ;
        RECT 2434.4200 1017.7400 2436.0200 1018.2200 ;
        RECT 2434.4200 995.9800 2436.0200 996.4600 ;
        RECT 2434.4200 1001.4200 2436.0200 1001.9000 ;
        RECT 2434.4200 1006.8600 2436.0200 1007.3400 ;
        RECT 2434.4200 985.1000 2436.0200 985.5800 ;
        RECT 2434.4200 990.5400 2436.0200 991.0200 ;
        RECT 2397.0000 1066.7000 2398.6000 1067.1800 ;
        RECT 2397.0000 1072.1400 2398.6000 1072.6200 ;
        RECT 2397.0000 1077.5800 2398.6000 1078.0600 ;
        RECT 2397.0000 1055.8200 2398.6000 1056.3000 ;
        RECT 2397.0000 1061.2600 2398.6000 1061.7400 ;
        RECT 2397.0000 1039.5000 2398.6000 1039.9800 ;
        RECT 2397.0000 1044.9400 2398.6000 1045.4200 ;
        RECT 2397.0000 1050.3800 2398.6000 1050.8600 ;
        RECT 2397.0000 1023.1800 2398.6000 1023.6600 ;
        RECT 2397.0000 1028.6200 2398.6000 1029.1000 ;
        RECT 2397.0000 1034.0600 2398.6000 1034.5400 ;
        RECT 2397.0000 1012.3000 2398.6000 1012.7800 ;
        RECT 2397.0000 1017.7400 2398.6000 1018.2200 ;
        RECT 2397.0000 995.9800 2398.6000 996.4600 ;
        RECT 2397.0000 1001.4200 2398.6000 1001.9000 ;
        RECT 2397.0000 1006.8600 2398.6000 1007.3400 ;
        RECT 2397.0000 985.1000 2398.6000 985.5800 ;
        RECT 2397.0000 990.5400 2398.6000 991.0200 ;
        RECT 2434.4200 968.7800 2436.0200 969.2600 ;
        RECT 2434.4200 974.2200 2436.0200 974.7000 ;
        RECT 2434.4200 979.6600 2436.0200 980.1400 ;
        RECT 2434.4200 957.9000 2436.0200 958.3800 ;
        RECT 2434.4200 963.3400 2436.0200 963.8200 ;
        RECT 2434.4200 941.5800 2436.0200 942.0600 ;
        RECT 2434.4200 947.0200 2436.0200 947.5000 ;
        RECT 2434.4200 952.4600 2436.0200 952.9400 ;
        RECT 2434.4200 930.7000 2436.0200 931.1800 ;
        RECT 2434.4200 936.1400 2436.0200 936.6200 ;
        RECT 2434.4200 914.3800 2436.0200 914.8600 ;
        RECT 2434.4200 919.8200 2436.0200 920.3000 ;
        RECT 2434.4200 925.2600 2436.0200 925.7400 ;
        RECT 2434.4200 903.5000 2436.0200 903.9800 ;
        RECT 2434.4200 908.9400 2436.0200 909.4200 ;
        RECT 2434.4200 887.1800 2436.0200 887.6600 ;
        RECT 2434.4200 892.6200 2436.0200 893.1000 ;
        RECT 2434.4200 898.0600 2436.0200 898.5400 ;
        RECT 2434.4200 881.7400 2436.0200 882.2200 ;
        RECT 2397.0000 968.7800 2398.6000 969.2600 ;
        RECT 2397.0000 974.2200 2398.6000 974.7000 ;
        RECT 2397.0000 979.6600 2398.6000 980.1400 ;
        RECT 2397.0000 957.9000 2398.6000 958.3800 ;
        RECT 2397.0000 963.3400 2398.6000 963.8200 ;
        RECT 2397.0000 941.5800 2398.6000 942.0600 ;
        RECT 2397.0000 947.0200 2398.6000 947.5000 ;
        RECT 2397.0000 952.4600 2398.6000 952.9400 ;
        RECT 2397.0000 930.7000 2398.6000 931.1800 ;
        RECT 2397.0000 936.1400 2398.6000 936.6200 ;
        RECT 2397.0000 914.3800 2398.6000 914.8600 ;
        RECT 2397.0000 919.8200 2398.6000 920.3000 ;
        RECT 2397.0000 925.2600 2398.6000 925.7400 ;
        RECT 2397.0000 903.5000 2398.6000 903.9800 ;
        RECT 2397.0000 908.9400 2398.6000 909.4200 ;
        RECT 2397.0000 887.1800 2398.6000 887.6600 ;
        RECT 2397.0000 892.6200 2398.6000 893.1000 ;
        RECT 2397.0000 898.0600 2398.6000 898.5400 ;
        RECT 2397.0000 881.7400 2398.6000 882.2200 ;
        RECT 2391.4400 1084.0500 2441.5800 1085.6500 ;
        RECT 2391.4400 877.5500 2441.5800 879.1500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 872.1200 2398.6000 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 1090.1600 2398.6000 1091.7600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 872.1200 2436.0200 873.7200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 1090.1600 2436.0200 1091.7600 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 877.5500 2393.0400 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 877.5500 2441.5800 879.1500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 1084.0500 2393.0400 1085.6500 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 1084.0500 2441.5800 1085.6500 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 642.4800 2436.0200 862.1200 ;
        RECT 2397.0000 642.4800 2398.6000 862.1200 ;
      LAYER met3 ;
        RECT 2434.4200 837.0600 2436.0200 837.5400 ;
        RECT 2434.4200 842.5000 2436.0200 842.9800 ;
        RECT 2434.4200 847.9400 2436.0200 848.4200 ;
        RECT 2434.4200 826.1800 2436.0200 826.6600 ;
        RECT 2434.4200 831.6200 2436.0200 832.1000 ;
        RECT 2434.4200 809.8600 2436.0200 810.3400 ;
        RECT 2434.4200 815.3000 2436.0200 815.7800 ;
        RECT 2434.4200 820.7400 2436.0200 821.2200 ;
        RECT 2434.4200 793.5400 2436.0200 794.0200 ;
        RECT 2434.4200 798.9800 2436.0200 799.4600 ;
        RECT 2434.4200 804.4200 2436.0200 804.9000 ;
        RECT 2434.4200 782.6600 2436.0200 783.1400 ;
        RECT 2434.4200 788.1000 2436.0200 788.5800 ;
        RECT 2434.4200 766.3400 2436.0200 766.8200 ;
        RECT 2434.4200 771.7800 2436.0200 772.2600 ;
        RECT 2434.4200 777.2200 2436.0200 777.7000 ;
        RECT 2434.4200 755.4600 2436.0200 755.9400 ;
        RECT 2434.4200 760.9000 2436.0200 761.3800 ;
        RECT 2397.0000 837.0600 2398.6000 837.5400 ;
        RECT 2397.0000 842.5000 2398.6000 842.9800 ;
        RECT 2397.0000 847.9400 2398.6000 848.4200 ;
        RECT 2397.0000 826.1800 2398.6000 826.6600 ;
        RECT 2397.0000 831.6200 2398.6000 832.1000 ;
        RECT 2397.0000 809.8600 2398.6000 810.3400 ;
        RECT 2397.0000 815.3000 2398.6000 815.7800 ;
        RECT 2397.0000 820.7400 2398.6000 821.2200 ;
        RECT 2397.0000 793.5400 2398.6000 794.0200 ;
        RECT 2397.0000 798.9800 2398.6000 799.4600 ;
        RECT 2397.0000 804.4200 2398.6000 804.9000 ;
        RECT 2397.0000 782.6600 2398.6000 783.1400 ;
        RECT 2397.0000 788.1000 2398.6000 788.5800 ;
        RECT 2397.0000 766.3400 2398.6000 766.8200 ;
        RECT 2397.0000 771.7800 2398.6000 772.2600 ;
        RECT 2397.0000 777.2200 2398.6000 777.7000 ;
        RECT 2397.0000 755.4600 2398.6000 755.9400 ;
        RECT 2397.0000 760.9000 2398.6000 761.3800 ;
        RECT 2434.4200 739.1400 2436.0200 739.6200 ;
        RECT 2434.4200 744.5800 2436.0200 745.0600 ;
        RECT 2434.4200 750.0200 2436.0200 750.5000 ;
        RECT 2434.4200 728.2600 2436.0200 728.7400 ;
        RECT 2434.4200 733.7000 2436.0200 734.1800 ;
        RECT 2434.4200 711.9400 2436.0200 712.4200 ;
        RECT 2434.4200 717.3800 2436.0200 717.8600 ;
        RECT 2434.4200 722.8200 2436.0200 723.3000 ;
        RECT 2434.4200 701.0600 2436.0200 701.5400 ;
        RECT 2434.4200 706.5000 2436.0200 706.9800 ;
        RECT 2434.4200 684.7400 2436.0200 685.2200 ;
        RECT 2434.4200 690.1800 2436.0200 690.6600 ;
        RECT 2434.4200 695.6200 2436.0200 696.1000 ;
        RECT 2434.4200 673.8600 2436.0200 674.3400 ;
        RECT 2434.4200 679.3000 2436.0200 679.7800 ;
        RECT 2434.4200 657.5400 2436.0200 658.0200 ;
        RECT 2434.4200 662.9800 2436.0200 663.4600 ;
        RECT 2434.4200 668.4200 2436.0200 668.9000 ;
        RECT 2434.4200 652.1000 2436.0200 652.5800 ;
        RECT 2397.0000 739.1400 2398.6000 739.6200 ;
        RECT 2397.0000 744.5800 2398.6000 745.0600 ;
        RECT 2397.0000 750.0200 2398.6000 750.5000 ;
        RECT 2397.0000 728.2600 2398.6000 728.7400 ;
        RECT 2397.0000 733.7000 2398.6000 734.1800 ;
        RECT 2397.0000 711.9400 2398.6000 712.4200 ;
        RECT 2397.0000 717.3800 2398.6000 717.8600 ;
        RECT 2397.0000 722.8200 2398.6000 723.3000 ;
        RECT 2397.0000 701.0600 2398.6000 701.5400 ;
        RECT 2397.0000 706.5000 2398.6000 706.9800 ;
        RECT 2397.0000 684.7400 2398.6000 685.2200 ;
        RECT 2397.0000 690.1800 2398.6000 690.6600 ;
        RECT 2397.0000 695.6200 2398.6000 696.1000 ;
        RECT 2397.0000 673.8600 2398.6000 674.3400 ;
        RECT 2397.0000 679.3000 2398.6000 679.7800 ;
        RECT 2397.0000 657.5400 2398.6000 658.0200 ;
        RECT 2397.0000 662.9800 2398.6000 663.4600 ;
        RECT 2397.0000 668.4200 2398.6000 668.9000 ;
        RECT 2397.0000 652.1000 2398.6000 652.5800 ;
        RECT 2391.4400 854.4100 2441.5800 856.0100 ;
        RECT 2391.4400 647.9100 2441.5800 649.5100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 642.4800 2398.6000 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 860.5200 2398.6000 862.1200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 642.4800 2436.0200 644.0800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 860.5200 2436.0200 862.1200 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 647.9100 2393.0400 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 647.9100 2441.5800 649.5100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 854.4100 2393.0400 856.0100 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 854.4100 2441.5800 856.0100 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'E_CPU_IO'
    PORT
      LAYER met4 ;
        RECT 2434.4200 412.8400 2436.0200 632.4800 ;
        RECT 2397.0000 412.8400 2398.6000 632.4800 ;
      LAYER met3 ;
        RECT 2434.4200 607.4200 2436.0200 607.9000 ;
        RECT 2434.4200 612.8600 2436.0200 613.3400 ;
        RECT 2434.4200 618.3000 2436.0200 618.7800 ;
        RECT 2434.4200 596.5400 2436.0200 597.0200 ;
        RECT 2434.4200 601.9800 2436.0200 602.4600 ;
        RECT 2434.4200 580.2200 2436.0200 580.7000 ;
        RECT 2434.4200 585.6600 2436.0200 586.1400 ;
        RECT 2434.4200 591.1000 2436.0200 591.5800 ;
        RECT 2434.4200 563.9000 2436.0200 564.3800 ;
        RECT 2434.4200 569.3400 2436.0200 569.8200 ;
        RECT 2434.4200 574.7800 2436.0200 575.2600 ;
        RECT 2434.4200 553.0200 2436.0200 553.5000 ;
        RECT 2434.4200 558.4600 2436.0200 558.9400 ;
        RECT 2434.4200 536.7000 2436.0200 537.1800 ;
        RECT 2434.4200 542.1400 2436.0200 542.6200 ;
        RECT 2434.4200 547.5800 2436.0200 548.0600 ;
        RECT 2434.4200 525.8200 2436.0200 526.3000 ;
        RECT 2434.4200 531.2600 2436.0200 531.7400 ;
        RECT 2397.0000 607.4200 2398.6000 607.9000 ;
        RECT 2397.0000 612.8600 2398.6000 613.3400 ;
        RECT 2397.0000 618.3000 2398.6000 618.7800 ;
        RECT 2397.0000 596.5400 2398.6000 597.0200 ;
        RECT 2397.0000 601.9800 2398.6000 602.4600 ;
        RECT 2397.0000 580.2200 2398.6000 580.7000 ;
        RECT 2397.0000 585.6600 2398.6000 586.1400 ;
        RECT 2397.0000 591.1000 2398.6000 591.5800 ;
        RECT 2397.0000 563.9000 2398.6000 564.3800 ;
        RECT 2397.0000 569.3400 2398.6000 569.8200 ;
        RECT 2397.0000 574.7800 2398.6000 575.2600 ;
        RECT 2397.0000 553.0200 2398.6000 553.5000 ;
        RECT 2397.0000 558.4600 2398.6000 558.9400 ;
        RECT 2397.0000 536.7000 2398.6000 537.1800 ;
        RECT 2397.0000 542.1400 2398.6000 542.6200 ;
        RECT 2397.0000 547.5800 2398.6000 548.0600 ;
        RECT 2397.0000 525.8200 2398.6000 526.3000 ;
        RECT 2397.0000 531.2600 2398.6000 531.7400 ;
        RECT 2434.4200 509.5000 2436.0200 509.9800 ;
        RECT 2434.4200 514.9400 2436.0200 515.4200 ;
        RECT 2434.4200 520.3800 2436.0200 520.8600 ;
        RECT 2434.4200 498.6200 2436.0200 499.1000 ;
        RECT 2434.4200 504.0600 2436.0200 504.5400 ;
        RECT 2434.4200 482.3000 2436.0200 482.7800 ;
        RECT 2434.4200 487.7400 2436.0200 488.2200 ;
        RECT 2434.4200 493.1800 2436.0200 493.6600 ;
        RECT 2434.4200 471.4200 2436.0200 471.9000 ;
        RECT 2434.4200 476.8600 2436.0200 477.3400 ;
        RECT 2434.4200 455.1000 2436.0200 455.5800 ;
        RECT 2434.4200 460.5400 2436.0200 461.0200 ;
        RECT 2434.4200 465.9800 2436.0200 466.4600 ;
        RECT 2434.4200 444.2200 2436.0200 444.7000 ;
        RECT 2434.4200 449.6600 2436.0200 450.1400 ;
        RECT 2434.4200 427.9000 2436.0200 428.3800 ;
        RECT 2434.4200 433.3400 2436.0200 433.8200 ;
        RECT 2434.4200 438.7800 2436.0200 439.2600 ;
        RECT 2434.4200 422.4600 2436.0200 422.9400 ;
        RECT 2397.0000 509.5000 2398.6000 509.9800 ;
        RECT 2397.0000 514.9400 2398.6000 515.4200 ;
        RECT 2397.0000 520.3800 2398.6000 520.8600 ;
        RECT 2397.0000 498.6200 2398.6000 499.1000 ;
        RECT 2397.0000 504.0600 2398.6000 504.5400 ;
        RECT 2397.0000 482.3000 2398.6000 482.7800 ;
        RECT 2397.0000 487.7400 2398.6000 488.2200 ;
        RECT 2397.0000 493.1800 2398.6000 493.6600 ;
        RECT 2397.0000 471.4200 2398.6000 471.9000 ;
        RECT 2397.0000 476.8600 2398.6000 477.3400 ;
        RECT 2397.0000 455.1000 2398.6000 455.5800 ;
        RECT 2397.0000 460.5400 2398.6000 461.0200 ;
        RECT 2397.0000 465.9800 2398.6000 466.4600 ;
        RECT 2397.0000 444.2200 2398.6000 444.7000 ;
        RECT 2397.0000 449.6600 2398.6000 450.1400 ;
        RECT 2397.0000 427.9000 2398.6000 428.3800 ;
        RECT 2397.0000 433.3400 2398.6000 433.8200 ;
        RECT 2397.0000 438.7800 2398.6000 439.2600 ;
        RECT 2397.0000 422.4600 2398.6000 422.9400 ;
        RECT 2391.4400 624.7700 2441.5800 626.3700 ;
        RECT 2391.4400 418.2700 2441.5800 419.8700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 412.8400 2398.6000 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2397.0000 630.8800 2398.6000 632.4800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 412.8400 2436.0200 414.4400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2434.4200 630.8800 2436.0200 632.4800 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 418.2700 2393.0400 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 418.2700 2441.5800 419.8700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2391.4400 624.7700 2393.0400 626.3700 ;
    END
    PORT
      LAYER met3 ;
        RECT 2439.9800 624.7700 2441.5800 626.3700 ;
    END
# end of P/G pin shape extracted from block 'E_CPU_IO'


# P/G pin shape extracted from block 'wb_mem_split'
    PORT
      LAYER met4 ;
        RECT 521.1600 505.3800 649.4800 506.9800 ;
    END
# end of P/G pin shape extracted from block 'wb_mem_split'

  END vccd1
  OBS
    LAYER li1 ;
      RECT 0.0000 0.0000 3370.4200 2569.7200 ;
    LAYER met1 ;
      RECT 0.0000 0.0000 3370.4200 2569.7200 ;
    LAYER met2 ;
      RECT 0.0000 0.6250 3370.4200 2569.7200 ;
      RECT 3000.1000 0.0000 3370.4200 0.6250 ;
      RECT 2924.2000 0.0000 2999.6800 0.6250 ;
      RECT 2847.8400 0.0000 2923.7800 0.6250 ;
      RECT 2771.4800 0.0000 2847.4200 0.6250 ;
      RECT 2695.1200 0.0000 2771.0600 0.6250 ;
      RECT 2618.7600 0.0000 2694.7000 0.6250 ;
      RECT 2542.4000 0.0000 2618.3400 0.6250 ;
      RECT 2466.0400 0.0000 2541.9800 0.6250 ;
      RECT 2389.6800 0.0000 2465.6200 0.6250 ;
      RECT 2313.3200 0.0000 2389.2600 0.6250 ;
      RECT 2237.4200 0.0000 2312.9000 0.6250 ;
      RECT 2161.0600 0.0000 2237.0000 0.6250 ;
      RECT 2084.7000 0.0000 2160.6400 0.6250 ;
      RECT 2008.3400 0.0000 2084.2800 0.6250 ;
      RECT 1931.9800 0.0000 2007.9200 0.6250 ;
      RECT 1855.6200 0.0000 1931.5600 0.6250 ;
      RECT 1779.2600 0.0000 1855.2000 0.6250 ;
      RECT 1702.9000 0.0000 1778.8400 0.6250 ;
      RECT 1626.5400 0.0000 1702.4800 0.6250 ;
      RECT 1550.1800 0.0000 1626.1200 0.6250 ;
      RECT 1474.2800 0.0000 1549.7600 0.6250 ;
      RECT 1397.9200 0.0000 1473.8600 0.6250 ;
      RECT 1321.5600 0.0000 1397.5000 0.6250 ;
      RECT 1245.2000 0.0000 1321.1400 0.6250 ;
      RECT 1168.8400 0.0000 1244.7800 0.6250 ;
      RECT 1092.4800 0.0000 1168.4200 0.6250 ;
      RECT 1016.1200 0.0000 1092.0600 0.6250 ;
      RECT 939.7600 0.0000 1015.7000 0.6250 ;
      RECT 863.4000 0.0000 939.3400 0.6250 ;
      RECT 787.5000 0.0000 862.9800 0.6250 ;
      RECT 711.1400 0.0000 787.0800 0.6250 ;
      RECT 668.3600 0.0000 710.7200 0.6250 ;
      RECT 649.0400 0.0000 667.9400 0.6250 ;
      RECT 634.7800 0.0000 648.6200 0.6250 ;
      RECT 558.4200 0.0000 634.3600 0.6250 ;
      RECT 518.8600 0.0000 558.0000 0.6250 ;
      RECT 505.9800 0.0000 518.4400 0.6250 ;
      RECT 482.0600 0.0000 505.5600 0.6250 ;
      RECT 405.7000 0.0000 481.6400 0.6250 ;
      RECT 329.3400 0.0000 405.2800 0.6250 ;
      RECT 252.9800 0.0000 328.9200 0.6250 ;
      RECT 176.6200 0.0000 252.5600 0.6250 ;
      RECT 100.7200 0.0000 176.2000 0.6250 ;
      RECT 0.0000 0.0000 100.3000 0.6250 ;
    LAYER met3 ;
      RECT 0.0000 2568.0200 3370.4200 2569.7200 ;
      RECT 3368.7200 2564.4200 3370.4200 2568.0200 ;
      RECT 0.0000 2564.4200 1.7000 2568.0200 ;
      RECT 0.0000 2564.1200 3370.4200 2564.4200 ;
      RECT 1065.0600 2564.0200 3370.4200 2564.1200 ;
      RECT 0.0000 2564.0200 1062.5200 2564.1200 ;
      RECT 3364.7200 2560.4200 3370.4200 2564.0200 ;
      RECT 0.0000 2560.4200 5.7000 2564.0200 ;
      RECT 1065.0600 2559.0400 3370.4200 2560.4200 ;
      RECT 0.0000 2559.0400 1062.5200 2560.4200 ;
      RECT 1065.0600 2558.7200 1065.5600 2559.0400 ;
      RECT 1057.5000 2558.7200 1062.5200 2559.0400 ;
      RECT 3364.7200 2557.9600 3370.4200 2559.0400 ;
      RECT 3307.6200 2557.9600 3361.1200 2559.0400 ;
      RECT 2494.8200 2557.9600 3305.4200 2559.0400 ;
      RECT 2449.0800 2557.9600 2492.6200 2559.0400 ;
      RECT 2438.9200 2557.9600 2446.8800 2559.0400 ;
      RECT 2388.9400 2557.9600 2436.7200 2559.0400 ;
      RECT 2378.6800 2557.9600 2386.7400 2559.0400 ;
      RECT 2176.1800 2557.9600 2376.4800 2559.0400 ;
      RECT 2168.7200 2557.9600 2173.9800 2559.0400 ;
      RECT 2158.4600 2557.9600 2166.5200 2559.0400 ;
      RECT 1955.9600 2557.9600 2156.2600 2559.0400 ;
      RECT 1948.5000 2557.9600 1953.7600 2559.0400 ;
      RECT 1938.2400 2557.9600 1946.3000 2559.0400 ;
      RECT 1735.7400 2557.9600 1936.0400 2559.0400 ;
      RECT 1728.2800 2557.9600 1733.5400 2559.0400 ;
      RECT 1718.0200 2557.9600 1726.0800 2559.0400 ;
      RECT 1515.5200 2557.9600 1715.8200 2559.0400 ;
      RECT 1508.0600 2557.9600 1513.3200 2559.0400 ;
      RECT 1497.8000 2557.9600 1505.8600 2559.0400 ;
      RECT 1295.3000 2557.9600 1495.6000 2559.0400 ;
      RECT 1287.9800 2557.9600 1293.1000 2559.0400 ;
      RECT 1277.5800 2557.9600 1285.6400 2559.0400 ;
      RECT 1075.0800 2557.9600 1275.3800 2559.0400 ;
      RECT 1067.7600 2557.9600 1072.8800 2559.0400 ;
      RECT 1057.5000 2557.9600 1065.5600 2558.7200 ;
      RECT 1015.0800 2557.9600 1055.3000 2559.0400 ;
      RECT 1004.8200 2557.9600 1012.8800 2559.0400 ;
      RECT 9.3000 2557.9600 1002.6200 2559.0400 ;
      RECT 0.0000 2557.9600 5.7000 2559.0400 ;
      RECT 0.0000 2556.3200 3370.4200 2557.9600 ;
      RECT 3368.7200 2555.2400 3370.4200 2556.3200 ;
      RECT 3305.0200 2555.2400 3365.1200 2556.3200 ;
      RECT 2497.4200 2555.2400 3302.8200 2556.3200 ;
      RECT 2446.4800 2555.2400 2495.2200 2556.3200 ;
      RECT 2436.3200 2555.2400 2444.2800 2556.3200 ;
      RECT 2398.9000 2555.2400 2434.1200 2556.3200 ;
      RECT 2386.3400 2555.2400 2396.7000 2556.3200 ;
      RECT 2376.2800 2555.2400 2384.1400 2556.3200 ;
      RECT 2178.5800 2555.2400 2374.0800 2556.3200 ;
      RECT 2166.1200 2555.2400 2176.3800 2556.3200 ;
      RECT 2156.0600 2555.2400 2163.9200 2556.3200 ;
      RECT 1958.3600 2555.2400 2153.8600 2556.3200 ;
      RECT 1945.9000 2555.2400 1956.1600 2556.3200 ;
      RECT 1935.8400 2555.2400 1943.7000 2556.3200 ;
      RECT 1738.1400 2555.2400 1933.6400 2556.3200 ;
      RECT 1725.6800 2555.2400 1735.9400 2556.3200 ;
      RECT 1715.6200 2555.2400 1723.4800 2556.3200 ;
      RECT 1517.9200 2555.2400 1713.4200 2556.3200 ;
      RECT 1505.4600 2555.2400 1515.7200 2556.3200 ;
      RECT 1495.4000 2555.2400 1503.2600 2556.3200 ;
      RECT 1297.7000 2555.2400 1493.2000 2556.3200 ;
      RECT 1285.3800 2555.2400 1295.5000 2556.3200 ;
      RECT 1275.1800 2555.2400 1283.0400 2556.3200 ;
      RECT 1077.4800 2555.2400 1272.9800 2556.3200 ;
      RECT 1065.1600 2555.2400 1075.2800 2556.3200 ;
      RECT 1055.1000 2555.2400 1062.9600 2556.3200 ;
      RECT 1017.4800 2555.2400 1052.9000 2556.3200 ;
      RECT 1007.4200 2555.2400 1015.2800 2556.3200 ;
      RECT 5.3000 2555.2400 1005.2200 2556.3200 ;
      RECT 0.0000 2555.2400 1.7000 2556.3200 ;
      RECT 0.0000 2553.6000 3370.4200 2555.2400 ;
      RECT 3364.7200 2552.5200 3370.4200 2553.6000 ;
      RECT 3307.6200 2552.5200 3361.1200 2553.6000 ;
      RECT 2494.8200 2552.5200 3305.4200 2553.6000 ;
      RECT 2449.0800 2552.5200 2492.6200 2553.6000 ;
      RECT 2438.9200 2552.5200 2446.8800 2553.6000 ;
      RECT 2388.9400 2552.5200 2436.7200 2553.6000 ;
      RECT 2378.6800 2552.5200 2386.7400 2553.6000 ;
      RECT 2176.1800 2552.5200 2376.4800 2553.6000 ;
      RECT 2168.7200 2552.5200 2173.9800 2553.6000 ;
      RECT 2158.4600 2552.5200 2166.5200 2553.6000 ;
      RECT 1955.9600 2552.5200 2156.2600 2553.6000 ;
      RECT 1948.5000 2552.5200 1953.7600 2553.6000 ;
      RECT 1938.2400 2552.5200 1946.3000 2553.6000 ;
      RECT 1735.7400 2552.5200 1936.0400 2553.6000 ;
      RECT 1728.2800 2552.5200 1733.5400 2553.6000 ;
      RECT 1718.0200 2552.5200 1726.0800 2553.6000 ;
      RECT 1515.5200 2552.5200 1715.8200 2553.6000 ;
      RECT 1508.0600 2552.5200 1513.3200 2553.6000 ;
      RECT 1497.8000 2552.5200 1505.8600 2553.6000 ;
      RECT 1295.3000 2552.5200 1495.6000 2553.6000 ;
      RECT 1287.9800 2552.5200 1293.1000 2553.6000 ;
      RECT 1277.5800 2552.5200 1285.6400 2553.6000 ;
      RECT 1075.0800 2552.5200 1275.3800 2553.6000 ;
      RECT 1067.7600 2552.5200 1072.8800 2553.6000 ;
      RECT 1057.5000 2552.5200 1065.5600 2553.6000 ;
      RECT 1015.0800 2552.5200 1055.3000 2553.6000 ;
      RECT 1004.8200 2552.5200 1012.8800 2553.6000 ;
      RECT 9.3000 2552.5200 1002.6200 2553.6000 ;
      RECT 0.0000 2552.5200 5.7000 2553.6000 ;
      RECT 0.0000 2550.8800 3370.4200 2552.5200 ;
      RECT 3368.7200 2549.8000 3370.4200 2550.8800 ;
      RECT 3305.0200 2549.8000 3365.1200 2550.8800 ;
      RECT 2497.4200 2549.8000 3302.8200 2550.8800 ;
      RECT 2446.4800 2549.8000 2495.2200 2550.8800 ;
      RECT 2436.3200 2549.8000 2444.2800 2550.8800 ;
      RECT 2398.9000 2549.8000 2434.1200 2550.8800 ;
      RECT 2386.3400 2549.8000 2396.7000 2550.8800 ;
      RECT 2376.2800 2549.8000 2384.1400 2550.8800 ;
      RECT 2178.5800 2549.8000 2374.0800 2550.8800 ;
      RECT 2166.1200 2549.8000 2176.3800 2550.8800 ;
      RECT 2156.0600 2549.8000 2163.9200 2550.8800 ;
      RECT 1958.3600 2549.8000 2153.8600 2550.8800 ;
      RECT 1945.9000 2549.8000 1956.1600 2550.8800 ;
      RECT 1935.8400 2549.8000 1943.7000 2550.8800 ;
      RECT 1738.1400 2549.8000 1933.6400 2550.8800 ;
      RECT 1725.6800 2549.8000 1735.9400 2550.8800 ;
      RECT 1715.6200 2549.8000 1723.4800 2550.8800 ;
      RECT 1517.9200 2549.8000 1713.4200 2550.8800 ;
      RECT 1505.4600 2549.8000 1515.7200 2550.8800 ;
      RECT 1495.4000 2549.8000 1503.2600 2550.8800 ;
      RECT 1297.7000 2549.8000 1493.2000 2550.8800 ;
      RECT 1285.3800 2549.8000 1295.5000 2550.8800 ;
      RECT 1275.1800 2549.8000 1283.0400 2550.8800 ;
      RECT 1077.4800 2549.8000 1272.9800 2550.8800 ;
      RECT 1065.1600 2549.8000 1075.2800 2550.8800 ;
      RECT 1055.1000 2549.8000 1062.9600 2550.8800 ;
      RECT 1017.4800 2549.8000 1052.9000 2550.8800 ;
      RECT 1007.4200 2549.8000 1015.2800 2550.8800 ;
      RECT 5.3000 2549.8000 1005.2200 2550.8800 ;
      RECT 0.0000 2549.8000 1.7000 2550.8800 ;
      RECT 0.0000 2548.1600 3370.4200 2549.8000 ;
      RECT 3364.7200 2547.0800 3370.4200 2548.1600 ;
      RECT 3307.6200 2547.0800 3361.1200 2548.1600 ;
      RECT 2494.8200 2547.0800 3305.4200 2548.1600 ;
      RECT 2449.0800 2547.0800 2492.6200 2548.1600 ;
      RECT 2438.9200 2547.0800 2446.8800 2548.1600 ;
      RECT 2388.9400 2547.0800 2436.7200 2548.1600 ;
      RECT 2378.6800 2547.0800 2386.7400 2548.1600 ;
      RECT 2176.1800 2547.0800 2376.4800 2548.1600 ;
      RECT 2168.7200 2547.0800 2173.9800 2548.1600 ;
      RECT 2158.4600 2547.0800 2166.5200 2548.1600 ;
      RECT 1955.9600 2547.0800 2156.2600 2548.1600 ;
      RECT 1948.5000 2547.0800 1953.7600 2548.1600 ;
      RECT 1938.2400 2547.0800 1946.3000 2548.1600 ;
      RECT 1735.7400 2547.0800 1936.0400 2548.1600 ;
      RECT 1728.2800 2547.0800 1733.5400 2548.1600 ;
      RECT 1718.0200 2547.0800 1726.0800 2548.1600 ;
      RECT 1515.5200 2547.0800 1715.8200 2548.1600 ;
      RECT 1508.0600 2547.0800 1513.3200 2548.1600 ;
      RECT 1497.8000 2547.0800 1505.8600 2548.1600 ;
      RECT 1295.3000 2547.0800 1495.6000 2548.1600 ;
      RECT 1287.9800 2547.0800 1293.1000 2548.1600 ;
      RECT 1277.5800 2547.0800 1285.6400 2548.1600 ;
      RECT 1075.0800 2547.0800 1275.3800 2548.1600 ;
      RECT 1067.7600 2547.0800 1072.8800 2548.1600 ;
      RECT 1057.5000 2547.0800 1065.5600 2548.1600 ;
      RECT 1015.0800 2547.0800 1055.3000 2548.1600 ;
      RECT 1004.8200 2547.0800 1012.8800 2548.1600 ;
      RECT 9.3000 2547.0800 1002.6200 2548.1600 ;
      RECT 0.0000 2547.0800 5.7000 2548.1600 ;
      RECT 0.0000 2545.4400 3370.4200 2547.0800 ;
      RECT 3368.7200 2544.3600 3370.4200 2545.4400 ;
      RECT 3305.0200 2544.3600 3365.1200 2545.4400 ;
      RECT 2497.4200 2544.3600 3302.8200 2545.4400 ;
      RECT 2446.4800 2544.3600 2495.2200 2545.4400 ;
      RECT 2436.3200 2544.3600 2444.2800 2545.4400 ;
      RECT 2398.9000 2544.3600 2434.1200 2545.4400 ;
      RECT 2386.3400 2544.3600 2396.7000 2545.4400 ;
      RECT 2376.2800 2544.3600 2384.1400 2545.4400 ;
      RECT 2178.5800 2544.3600 2374.0800 2545.4400 ;
      RECT 2166.1200 2544.3600 2176.3800 2545.4400 ;
      RECT 2156.0600 2544.3600 2163.9200 2545.4400 ;
      RECT 1958.3600 2544.3600 2153.8600 2545.4400 ;
      RECT 1945.9000 2544.3600 1956.1600 2545.4400 ;
      RECT 1935.8400 2544.3600 1943.7000 2545.4400 ;
      RECT 1738.1400 2544.3600 1933.6400 2545.4400 ;
      RECT 1725.6800 2544.3600 1735.9400 2545.4400 ;
      RECT 1715.6200 2544.3600 1723.4800 2545.4400 ;
      RECT 1517.9200 2544.3600 1713.4200 2545.4400 ;
      RECT 1505.4600 2544.3600 1515.7200 2545.4400 ;
      RECT 1495.4000 2544.3600 1503.2600 2545.4400 ;
      RECT 1297.7000 2544.3600 1493.2000 2545.4400 ;
      RECT 1285.3800 2544.3600 1295.5000 2545.4400 ;
      RECT 1275.1800 2544.3600 1283.0400 2545.4400 ;
      RECT 1077.4800 2544.3600 1272.9800 2545.4400 ;
      RECT 1065.1600 2544.3600 1075.2800 2545.4400 ;
      RECT 1055.1000 2544.3600 1062.9600 2545.4400 ;
      RECT 1017.4800 2544.3600 1052.9000 2545.4400 ;
      RECT 1007.4200 2544.3600 1015.2800 2545.4400 ;
      RECT 5.3000 2544.3600 1005.2200 2545.4400 ;
      RECT 0.0000 2544.3600 1.7000 2545.4400 ;
      RECT 0.0000 2542.7200 3370.4200 2544.3600 ;
      RECT 3364.7200 2541.6400 3370.4200 2542.7200 ;
      RECT 3307.6200 2541.6400 3361.1200 2542.7200 ;
      RECT 2494.8200 2541.6400 3305.4200 2542.7200 ;
      RECT 2449.0800 2541.6400 2492.6200 2542.7200 ;
      RECT 2438.9200 2541.6400 2446.8800 2542.7200 ;
      RECT 2388.9400 2541.6400 2436.7200 2542.7200 ;
      RECT 2378.6800 2541.6400 2386.7400 2542.7200 ;
      RECT 2176.1800 2541.6400 2376.4800 2542.7200 ;
      RECT 2168.7200 2541.6400 2173.9800 2542.7200 ;
      RECT 2158.4600 2541.6400 2166.5200 2542.7200 ;
      RECT 1955.9600 2541.6400 2156.2600 2542.7200 ;
      RECT 1948.5000 2541.6400 1953.7600 2542.7200 ;
      RECT 1938.2400 2541.6400 1946.3000 2542.7200 ;
      RECT 1735.7400 2541.6400 1936.0400 2542.7200 ;
      RECT 1728.2800 2541.6400 1733.5400 2542.7200 ;
      RECT 1718.0200 2541.6400 1726.0800 2542.7200 ;
      RECT 1515.5200 2541.6400 1715.8200 2542.7200 ;
      RECT 1508.0600 2541.6400 1513.3200 2542.7200 ;
      RECT 1497.8000 2541.6400 1505.8600 2542.7200 ;
      RECT 1295.3000 2541.6400 1495.6000 2542.7200 ;
      RECT 1287.9800 2541.6400 1293.1000 2542.7200 ;
      RECT 1277.5800 2541.6400 1285.6400 2542.7200 ;
      RECT 1075.0800 2541.6400 1275.3800 2542.7200 ;
      RECT 1067.7600 2541.6400 1072.8800 2542.7200 ;
      RECT 1057.5000 2541.6400 1065.5600 2542.7200 ;
      RECT 1015.0800 2541.6400 1055.3000 2542.7200 ;
      RECT 1004.8200 2541.6400 1012.8800 2542.7200 ;
      RECT 9.3000 2541.6400 1002.6200 2542.7200 ;
      RECT 0.0000 2541.6400 5.7000 2542.7200 ;
      RECT 0.0000 2540.1500 3370.4200 2541.6400 ;
      RECT 1.1000 2540.0000 3370.4200 2540.1500 ;
      RECT 1.1000 2539.2500 1.7000 2540.0000 ;
      RECT 3368.7200 2538.9200 3370.4200 2540.0000 ;
      RECT 3305.0200 2538.9200 3365.1200 2540.0000 ;
      RECT 2497.4200 2538.9200 3302.8200 2540.0000 ;
      RECT 2446.4800 2538.9200 2495.2200 2540.0000 ;
      RECT 2436.3200 2538.9200 2444.2800 2540.0000 ;
      RECT 2398.9000 2538.9200 2434.1200 2540.0000 ;
      RECT 2386.3400 2538.9200 2396.7000 2540.0000 ;
      RECT 2376.2800 2538.9200 2384.1400 2540.0000 ;
      RECT 2178.5800 2538.9200 2374.0800 2540.0000 ;
      RECT 2166.1200 2538.9200 2176.3800 2540.0000 ;
      RECT 2156.0600 2538.9200 2163.9200 2540.0000 ;
      RECT 1958.3600 2538.9200 2153.8600 2540.0000 ;
      RECT 1945.9000 2538.9200 1956.1600 2540.0000 ;
      RECT 1935.8400 2538.9200 1943.7000 2540.0000 ;
      RECT 1738.1400 2538.9200 1933.6400 2540.0000 ;
      RECT 1725.6800 2538.9200 1735.9400 2540.0000 ;
      RECT 1715.6200 2538.9200 1723.4800 2540.0000 ;
      RECT 1517.9200 2538.9200 1713.4200 2540.0000 ;
      RECT 1505.4600 2538.9200 1515.7200 2540.0000 ;
      RECT 1495.4000 2538.9200 1503.2600 2540.0000 ;
      RECT 1297.7000 2538.9200 1493.2000 2540.0000 ;
      RECT 1285.3800 2538.9200 1295.5000 2540.0000 ;
      RECT 1275.1800 2538.9200 1283.0400 2540.0000 ;
      RECT 1077.4800 2538.9200 1272.9800 2540.0000 ;
      RECT 1065.1600 2538.9200 1075.2800 2540.0000 ;
      RECT 1055.1000 2538.9200 1062.9600 2540.0000 ;
      RECT 1017.4800 2538.9200 1052.9000 2540.0000 ;
      RECT 1007.4200 2538.9200 1015.2800 2540.0000 ;
      RECT 5.3000 2538.9200 1005.2200 2540.0000 ;
      RECT 0.0000 2538.9200 1.7000 2539.2500 ;
      RECT 0.0000 2537.2800 3370.4200 2538.9200 ;
      RECT 3364.7200 2536.2000 3370.4200 2537.2800 ;
      RECT 3307.6200 2536.2000 3361.1200 2537.2800 ;
      RECT 2494.8200 2536.2000 3305.4200 2537.2800 ;
      RECT 2449.0800 2536.2000 2492.6200 2537.2800 ;
      RECT 2438.9200 2536.2000 2446.8800 2537.2800 ;
      RECT 2388.9400 2536.2000 2436.7200 2537.2800 ;
      RECT 2378.6800 2536.2000 2386.7400 2537.2800 ;
      RECT 2176.1800 2536.2000 2376.4800 2537.2800 ;
      RECT 2168.7200 2536.2000 2173.9800 2537.2800 ;
      RECT 2158.4600 2536.2000 2166.5200 2537.2800 ;
      RECT 1955.9600 2536.2000 2156.2600 2537.2800 ;
      RECT 1948.5000 2536.2000 1953.7600 2537.2800 ;
      RECT 1938.2400 2536.2000 1946.3000 2537.2800 ;
      RECT 1735.7400 2536.2000 1936.0400 2537.2800 ;
      RECT 1728.2800 2536.2000 1733.5400 2537.2800 ;
      RECT 1718.0200 2536.2000 1726.0800 2537.2800 ;
      RECT 1515.5200 2536.2000 1715.8200 2537.2800 ;
      RECT 1508.0600 2536.2000 1513.3200 2537.2800 ;
      RECT 1497.8000 2536.2000 1505.8600 2537.2800 ;
      RECT 1295.3000 2536.2000 1495.6000 2537.2800 ;
      RECT 1287.9800 2536.2000 1293.1000 2537.2800 ;
      RECT 1277.5800 2536.2000 1285.6400 2537.2800 ;
      RECT 1075.0800 2536.2000 1275.3800 2537.2800 ;
      RECT 1067.7600 2536.2000 1072.8800 2537.2800 ;
      RECT 1057.5000 2536.2000 1065.5600 2537.2800 ;
      RECT 1015.0800 2536.2000 1055.3000 2537.2800 ;
      RECT 1004.8200 2536.2000 1012.8800 2537.2800 ;
      RECT 9.3000 2536.2000 1002.6200 2537.2800 ;
      RECT 0.0000 2536.2000 5.7000 2537.2800 ;
      RECT 0.0000 2534.5600 3370.4200 2536.2000 ;
      RECT 3368.7200 2533.4800 3370.4200 2534.5600 ;
      RECT 3305.0200 2533.4800 3365.1200 2534.5600 ;
      RECT 2497.4200 2533.4800 3302.8200 2534.5600 ;
      RECT 2446.4800 2533.4800 2495.2200 2534.5600 ;
      RECT 2436.3200 2533.4800 2444.2800 2534.5600 ;
      RECT 2398.9000 2533.4800 2434.1200 2534.5600 ;
      RECT 2386.3400 2533.4800 2396.7000 2534.5600 ;
      RECT 2376.2800 2533.4800 2384.1400 2534.5600 ;
      RECT 2178.5800 2533.4800 2374.0800 2534.5600 ;
      RECT 2166.1200 2533.4800 2176.3800 2534.5600 ;
      RECT 2156.0600 2533.4800 2163.9200 2534.5600 ;
      RECT 1958.3600 2533.4800 2153.8600 2534.5600 ;
      RECT 1945.9000 2533.4800 1956.1600 2534.5600 ;
      RECT 1935.8400 2533.4800 1943.7000 2534.5600 ;
      RECT 1738.1400 2533.4800 1933.6400 2534.5600 ;
      RECT 1725.6800 2533.4800 1735.9400 2534.5600 ;
      RECT 1715.6200 2533.4800 1723.4800 2534.5600 ;
      RECT 1517.9200 2533.4800 1713.4200 2534.5600 ;
      RECT 1505.4600 2533.4800 1515.7200 2534.5600 ;
      RECT 1495.4000 2533.4800 1503.2600 2534.5600 ;
      RECT 1297.7000 2533.4800 1493.2000 2534.5600 ;
      RECT 1285.3800 2533.4800 1295.5000 2534.5600 ;
      RECT 1275.1800 2533.4800 1283.0400 2534.5600 ;
      RECT 1077.4800 2533.4800 1272.9800 2534.5600 ;
      RECT 1065.1600 2533.4800 1075.2800 2534.5600 ;
      RECT 1055.1000 2533.4800 1062.9600 2534.5600 ;
      RECT 1017.4800 2533.4800 1052.9000 2534.5600 ;
      RECT 1007.4200 2533.4800 1015.2800 2534.5600 ;
      RECT 5.3000 2533.4800 1005.2200 2534.5600 ;
      RECT 0.0000 2533.4800 1.7000 2534.5600 ;
      RECT 0.0000 2531.8400 3370.4200 2533.4800 ;
      RECT 3364.7200 2530.7600 3370.4200 2531.8400 ;
      RECT 3307.6200 2530.7600 3361.1200 2531.8400 ;
      RECT 2494.8200 2530.7600 3305.4200 2531.8400 ;
      RECT 2449.0800 2530.7600 2492.6200 2531.8400 ;
      RECT 2438.9200 2530.7600 2446.8800 2531.8400 ;
      RECT 2388.9400 2530.7600 2436.7200 2531.8400 ;
      RECT 2378.6800 2530.7600 2386.7400 2531.8400 ;
      RECT 2176.1800 2530.7600 2376.4800 2531.8400 ;
      RECT 2168.7200 2530.7600 2173.9800 2531.8400 ;
      RECT 2158.4600 2530.7600 2166.5200 2531.8400 ;
      RECT 1955.9600 2530.7600 2156.2600 2531.8400 ;
      RECT 1948.5000 2530.7600 1953.7600 2531.8400 ;
      RECT 1938.2400 2530.7600 1946.3000 2531.8400 ;
      RECT 1735.7400 2530.7600 1936.0400 2531.8400 ;
      RECT 1728.2800 2530.7600 1733.5400 2531.8400 ;
      RECT 1718.0200 2530.7600 1726.0800 2531.8400 ;
      RECT 1515.5200 2530.7600 1715.8200 2531.8400 ;
      RECT 1508.0600 2530.7600 1513.3200 2531.8400 ;
      RECT 1497.8000 2530.7600 1505.8600 2531.8400 ;
      RECT 1295.3000 2530.7600 1495.6000 2531.8400 ;
      RECT 1287.9800 2530.7600 1293.1000 2531.8400 ;
      RECT 1277.5800 2530.7600 1285.6400 2531.8400 ;
      RECT 1075.0800 2530.7600 1275.3800 2531.8400 ;
      RECT 1067.7600 2530.7600 1072.8800 2531.8400 ;
      RECT 1057.5000 2530.7600 1065.5600 2531.8400 ;
      RECT 1015.0800 2530.7600 1055.3000 2531.8400 ;
      RECT 1004.8200 2530.7600 1012.8800 2531.8400 ;
      RECT 9.3000 2530.7600 1002.6200 2531.8400 ;
      RECT 0.0000 2530.7600 5.7000 2531.8400 ;
      RECT 0.0000 2529.7800 3370.4200 2530.7600 ;
      RECT 1.1000 2529.1200 3370.4200 2529.7800 ;
      RECT 1.1000 2528.8800 1.7000 2529.1200 ;
      RECT 3368.7200 2528.0400 3370.4200 2529.1200 ;
      RECT 3305.0200 2528.0400 3365.1200 2529.1200 ;
      RECT 2497.4200 2528.0400 3302.8200 2529.1200 ;
      RECT 2446.4800 2528.0400 2495.2200 2529.1200 ;
      RECT 2436.3200 2528.0400 2444.2800 2529.1200 ;
      RECT 2398.9000 2528.0400 2434.1200 2529.1200 ;
      RECT 2386.3400 2528.0400 2396.7000 2529.1200 ;
      RECT 2376.2800 2528.0400 2384.1400 2529.1200 ;
      RECT 2178.5800 2528.0400 2374.0800 2529.1200 ;
      RECT 2166.1200 2528.0400 2176.3800 2529.1200 ;
      RECT 2156.0600 2528.0400 2163.9200 2529.1200 ;
      RECT 1958.3600 2528.0400 2153.8600 2529.1200 ;
      RECT 1945.9000 2528.0400 1956.1600 2529.1200 ;
      RECT 1935.8400 2528.0400 1943.7000 2529.1200 ;
      RECT 1738.1400 2528.0400 1933.6400 2529.1200 ;
      RECT 1725.6800 2528.0400 1735.9400 2529.1200 ;
      RECT 1715.6200 2528.0400 1723.4800 2529.1200 ;
      RECT 1517.9200 2528.0400 1713.4200 2529.1200 ;
      RECT 1505.4600 2528.0400 1515.7200 2529.1200 ;
      RECT 1495.4000 2528.0400 1503.2600 2529.1200 ;
      RECT 1297.7000 2528.0400 1493.2000 2529.1200 ;
      RECT 1285.3800 2528.0400 1295.5000 2529.1200 ;
      RECT 1275.1800 2528.0400 1283.0400 2529.1200 ;
      RECT 1077.4800 2528.0400 1272.9800 2529.1200 ;
      RECT 1065.1600 2528.0400 1075.2800 2529.1200 ;
      RECT 1055.1000 2528.0400 1062.9600 2529.1200 ;
      RECT 1017.4800 2528.0400 1052.9000 2529.1200 ;
      RECT 1007.4200 2528.0400 1015.2800 2529.1200 ;
      RECT 5.3000 2528.0400 1005.2200 2529.1200 ;
      RECT 0.0000 2528.0400 1.7000 2528.8800 ;
      RECT 0.0000 2526.4000 3370.4200 2528.0400 ;
      RECT 3364.7200 2525.3200 3370.4200 2526.4000 ;
      RECT 3307.6200 2525.3200 3361.1200 2526.4000 ;
      RECT 2494.8200 2525.3200 3305.4200 2526.4000 ;
      RECT 2449.0800 2525.3200 2492.6200 2526.4000 ;
      RECT 2438.9200 2525.3200 2446.8800 2526.4000 ;
      RECT 2388.9400 2525.3200 2436.7200 2526.4000 ;
      RECT 2378.6800 2525.3200 2386.7400 2526.4000 ;
      RECT 2176.1800 2525.3200 2376.4800 2526.4000 ;
      RECT 2168.7200 2525.3200 2173.9800 2526.4000 ;
      RECT 2158.4600 2525.3200 2166.5200 2526.4000 ;
      RECT 1955.9600 2525.3200 2156.2600 2526.4000 ;
      RECT 1948.5000 2525.3200 1953.7600 2526.4000 ;
      RECT 1938.2400 2525.3200 1946.3000 2526.4000 ;
      RECT 1735.7400 2525.3200 1936.0400 2526.4000 ;
      RECT 1728.2800 2525.3200 1733.5400 2526.4000 ;
      RECT 1718.0200 2525.3200 1726.0800 2526.4000 ;
      RECT 1515.5200 2525.3200 1715.8200 2526.4000 ;
      RECT 1508.0600 2525.3200 1513.3200 2526.4000 ;
      RECT 1497.8000 2525.3200 1505.8600 2526.4000 ;
      RECT 1295.3000 2525.3200 1495.6000 2526.4000 ;
      RECT 1287.9800 2525.3200 1293.1000 2526.4000 ;
      RECT 1277.5800 2525.3200 1285.6400 2526.4000 ;
      RECT 1075.0800 2525.3200 1275.3800 2526.4000 ;
      RECT 1067.7600 2525.3200 1072.8800 2526.4000 ;
      RECT 1057.5000 2525.3200 1065.5600 2526.4000 ;
      RECT 1015.0800 2525.3200 1055.3000 2526.4000 ;
      RECT 1004.8200 2525.3200 1012.8800 2526.4000 ;
      RECT 9.3000 2525.3200 1002.6200 2526.4000 ;
      RECT 0.0000 2525.3200 5.7000 2526.4000 ;
      RECT 0.0000 2523.6800 3370.4200 2525.3200 ;
      RECT 3368.7200 2522.6000 3370.4200 2523.6800 ;
      RECT 3305.0200 2522.6000 3365.1200 2523.6800 ;
      RECT 2497.4200 2522.6000 3302.8200 2523.6800 ;
      RECT 2446.4800 2522.6000 2495.2200 2523.6800 ;
      RECT 2436.3200 2522.6000 2444.2800 2523.6800 ;
      RECT 2398.9000 2522.6000 2434.1200 2523.6800 ;
      RECT 2386.3400 2522.6000 2396.7000 2523.6800 ;
      RECT 2376.2800 2522.6000 2384.1400 2523.6800 ;
      RECT 2178.5800 2522.6000 2374.0800 2523.6800 ;
      RECT 2166.1200 2522.6000 2176.3800 2523.6800 ;
      RECT 2156.0600 2522.6000 2163.9200 2523.6800 ;
      RECT 1958.3600 2522.6000 2153.8600 2523.6800 ;
      RECT 1945.9000 2522.6000 1956.1600 2523.6800 ;
      RECT 1935.8400 2522.6000 1943.7000 2523.6800 ;
      RECT 1738.1400 2522.6000 1933.6400 2523.6800 ;
      RECT 1725.6800 2522.6000 1735.9400 2523.6800 ;
      RECT 1715.6200 2522.6000 1723.4800 2523.6800 ;
      RECT 1517.9200 2522.6000 1713.4200 2523.6800 ;
      RECT 1505.4600 2522.6000 1515.7200 2523.6800 ;
      RECT 1495.4000 2522.6000 1503.2600 2523.6800 ;
      RECT 1297.7000 2522.6000 1493.2000 2523.6800 ;
      RECT 1285.3800 2522.6000 1295.5000 2523.6800 ;
      RECT 1275.1800 2522.6000 1283.0400 2523.6800 ;
      RECT 1077.4800 2522.6000 1272.9800 2523.6800 ;
      RECT 1065.1600 2522.6000 1075.2800 2523.6800 ;
      RECT 1055.1000 2522.6000 1062.9600 2523.6800 ;
      RECT 1017.4800 2522.6000 1052.9000 2523.6800 ;
      RECT 1007.4200 2522.6000 1015.2800 2523.6800 ;
      RECT 5.3000 2522.6000 1005.2200 2523.6800 ;
      RECT 0.0000 2522.6000 1.7000 2523.6800 ;
      RECT 0.0000 2520.9600 3370.4200 2522.6000 ;
      RECT 3364.7200 2519.8800 3370.4200 2520.9600 ;
      RECT 3307.6200 2519.8800 3361.1200 2520.9600 ;
      RECT 2494.8200 2519.8800 3305.4200 2520.9600 ;
      RECT 2449.0800 2519.8800 2492.6200 2520.9600 ;
      RECT 2438.9200 2519.8800 2446.8800 2520.9600 ;
      RECT 2388.9400 2519.8800 2436.7200 2520.9600 ;
      RECT 2378.6800 2519.8800 2386.7400 2520.9600 ;
      RECT 2176.1800 2519.8800 2376.4800 2520.9600 ;
      RECT 2168.7200 2519.8800 2173.9800 2520.9600 ;
      RECT 2158.4600 2519.8800 2166.5200 2520.9600 ;
      RECT 1955.9600 2519.8800 2156.2600 2520.9600 ;
      RECT 1948.5000 2519.8800 1953.7600 2520.9600 ;
      RECT 1938.2400 2519.8800 1946.3000 2520.9600 ;
      RECT 1735.7400 2519.8800 1936.0400 2520.9600 ;
      RECT 1728.2800 2519.8800 1733.5400 2520.9600 ;
      RECT 1718.0200 2519.8800 1726.0800 2520.9600 ;
      RECT 1515.5200 2519.8800 1715.8200 2520.9600 ;
      RECT 1508.0600 2519.8800 1513.3200 2520.9600 ;
      RECT 1497.8000 2519.8800 1505.8600 2520.9600 ;
      RECT 1295.3000 2519.8800 1495.6000 2520.9600 ;
      RECT 1287.9800 2519.8800 1293.1000 2520.9600 ;
      RECT 1277.5800 2519.8800 1285.6400 2520.9600 ;
      RECT 1075.0800 2519.8800 1275.3800 2520.9600 ;
      RECT 1067.7600 2519.8800 1072.8800 2520.9600 ;
      RECT 1057.5000 2519.8800 1065.5600 2520.9600 ;
      RECT 1015.0800 2519.8800 1055.3000 2520.9600 ;
      RECT 1004.8200 2519.8800 1012.8800 2520.9600 ;
      RECT 9.3000 2519.8800 1002.6200 2520.9600 ;
      RECT 0.0000 2519.8800 5.7000 2520.9600 ;
      RECT 0.0000 2518.8000 3370.4200 2519.8800 ;
      RECT 1.1000 2518.2400 3370.4200 2518.8000 ;
      RECT 1.1000 2517.9000 1.7000 2518.2400 ;
      RECT 3368.7200 2517.1600 3370.4200 2518.2400 ;
      RECT 3305.0200 2517.1600 3365.1200 2518.2400 ;
      RECT 2497.4200 2517.1600 3302.8200 2518.2400 ;
      RECT 2446.4800 2517.1600 2495.2200 2518.2400 ;
      RECT 2436.3200 2517.1600 2444.2800 2518.2400 ;
      RECT 2398.9000 2517.1600 2434.1200 2518.2400 ;
      RECT 2386.3400 2517.1600 2396.7000 2518.2400 ;
      RECT 1065.1600 2517.1600 2384.1400 2518.2400 ;
      RECT 1055.1000 2517.1600 1062.9600 2518.2400 ;
      RECT 1017.4800 2517.1600 1052.9000 2518.2400 ;
      RECT 1007.4200 2517.1600 1015.2800 2518.2400 ;
      RECT 5.3000 2517.1600 1005.2200 2518.2400 ;
      RECT 0.0000 2517.1600 1.7000 2517.9000 ;
      RECT 0.0000 2515.5200 3370.4200 2517.1600 ;
      RECT 3364.7200 2514.4400 3370.4200 2515.5200 ;
      RECT 3307.6200 2514.4400 3361.1200 2515.5200 ;
      RECT 2494.8200 2514.4400 3305.4200 2515.5200 ;
      RECT 2449.0800 2514.4400 2492.6200 2515.5200 ;
      RECT 2438.9200 2514.4400 2446.8800 2515.5200 ;
      RECT 2388.9400 2514.4400 2436.7200 2515.5200 ;
      RECT 1067.7600 2514.4400 2386.7400 2515.5200 ;
      RECT 1057.5000 2514.4400 1065.5600 2515.5200 ;
      RECT 1015.0800 2514.4400 1055.3000 2515.5200 ;
      RECT 1004.8200 2514.4400 1012.8800 2515.5200 ;
      RECT 9.3000 2514.4400 1002.6200 2515.5200 ;
      RECT 0.0000 2514.4400 5.7000 2515.5200 ;
      RECT 0.0000 2512.8000 3370.4200 2514.4400 ;
      RECT 3368.7200 2511.7200 3370.4200 2512.8000 ;
      RECT 3305.0200 2511.7200 3365.1200 2512.8000 ;
      RECT 2497.4200 2511.7200 3302.8200 2512.8000 ;
      RECT 2446.4800 2511.7200 2495.2200 2512.8000 ;
      RECT 2436.3200 2511.7200 2444.2800 2512.8000 ;
      RECT 2398.9000 2511.7200 2434.1200 2512.8000 ;
      RECT 2386.3400 2511.7200 2396.7000 2512.8000 ;
      RECT 1065.1600 2511.7200 2384.1400 2512.8000 ;
      RECT 1055.1000 2511.7200 1062.9600 2512.8000 ;
      RECT 1017.4800 2511.7200 1052.9000 2512.8000 ;
      RECT 1007.4200 2511.7200 1015.2800 2512.8000 ;
      RECT 5.3000 2511.7200 1005.2200 2512.8000 ;
      RECT 0.0000 2511.7200 1.7000 2512.8000 ;
      RECT 0.0000 2510.0800 3370.4200 2511.7200 ;
      RECT 3364.7200 2509.0000 3370.4200 2510.0800 ;
      RECT 3307.6200 2509.0000 3361.1200 2510.0800 ;
      RECT 2494.8200 2509.0000 3305.4200 2510.0800 ;
      RECT 2449.0800 2509.0000 2492.6200 2510.0800 ;
      RECT 2438.9200 2509.0000 2446.8800 2510.0800 ;
      RECT 2388.9400 2509.0000 2436.7200 2510.0800 ;
      RECT 1067.7600 2509.0000 2386.7400 2510.0800 ;
      RECT 1057.5000 2509.0000 1065.5600 2510.0800 ;
      RECT 1015.0800 2509.0000 1055.3000 2510.0800 ;
      RECT 1004.8200 2509.0000 1012.8800 2510.0800 ;
      RECT 9.3000 2509.0000 1002.6200 2510.0800 ;
      RECT 0.0000 2509.0000 5.7000 2510.0800 ;
      RECT 0.0000 2508.2100 3370.4200 2509.0000 ;
      RECT 0.0000 2507.8200 2384.1400 2508.2100 ;
      RECT 2386.3400 2507.4000 3370.4200 2508.2100 ;
      RECT 1.1000 2507.4000 2384.1400 2507.8200 ;
      RECT 2388.9400 2507.3600 3370.4200 2507.4000 ;
      RECT 1.1000 2507.3600 1065.5600 2507.4000 ;
      RECT 1.1000 2506.9200 1.7000 2507.3600 ;
      RECT 3368.7200 2506.2800 3370.4200 2507.3600 ;
      RECT 3305.0200 2506.2800 3365.1200 2507.3600 ;
      RECT 2497.4200 2506.2800 3302.8200 2507.3600 ;
      RECT 2446.4800 2506.2800 2495.2200 2507.3600 ;
      RECT 2436.3200 2506.2800 2444.2800 2507.3600 ;
      RECT 2398.9000 2506.2800 2434.1200 2507.3600 ;
      RECT 2388.9400 2506.2800 2396.7000 2507.3600 ;
      RECT 1065.1600 2506.2800 1065.5600 2507.3600 ;
      RECT 1055.1000 2506.2800 1062.9600 2507.3600 ;
      RECT 1017.4800 2506.2800 1052.9000 2507.3600 ;
      RECT 1007.4200 2506.2800 1015.2800 2507.3600 ;
      RECT 5.3000 2506.2800 1005.2200 2507.3600 ;
      RECT 0.0000 2506.2800 1.7000 2506.9200 ;
      RECT 2388.9400 2505.2000 3370.4200 2506.2800 ;
      RECT 2172.3200 2505.2000 2380.3400 2507.4000 ;
      RECT 1952.1000 2505.2000 2160.1200 2507.4000 ;
      RECT 1731.8800 2505.2000 1939.9000 2507.4000 ;
      RECT 1511.6600 2505.2000 1719.6800 2507.4000 ;
      RECT 1291.4400 2505.2000 1499.4600 2507.4000 ;
      RECT 1071.2200 2505.2000 1279.2400 2507.4000 ;
      RECT 1067.7600 2505.0000 3370.4200 2505.2000 ;
      RECT 0.0000 2505.0000 1065.5600 2506.2800 ;
      RECT 2386.3400 2504.6400 3370.4200 2505.0000 ;
      RECT 0.0000 2504.6400 1062.9600 2505.0000 ;
      RECT 3364.7200 2503.5600 3370.4200 2504.6400 ;
      RECT 3307.6200 2503.5600 3361.1200 2504.6400 ;
      RECT 2494.8200 2503.5600 3305.4200 2504.6400 ;
      RECT 2449.0800 2503.5600 2492.6200 2504.6400 ;
      RECT 2438.9200 2503.5600 2446.8800 2504.6400 ;
      RECT 2388.9400 2503.5600 2436.7200 2504.6400 ;
      RECT 2386.3400 2503.5600 2386.7400 2504.6400 ;
      RECT 1057.5000 2503.5600 1062.9600 2504.6400 ;
      RECT 1015.0800 2503.5600 1055.3000 2504.6400 ;
      RECT 1004.8200 2503.5600 1012.8800 2504.6400 ;
      RECT 9.3000 2503.5600 1002.6200 2504.6400 ;
      RECT 0.0000 2503.5600 5.7000 2504.6400 ;
      RECT 2386.3400 2502.8000 3370.4200 2503.5600 ;
      RECT 2172.3200 2502.8000 2380.3400 2505.0000 ;
      RECT 1952.1000 2502.8000 2160.1200 2505.0000 ;
      RECT 1731.8800 2502.8000 1939.9000 2505.0000 ;
      RECT 1511.6600 2502.8000 1719.6800 2505.0000 ;
      RECT 1291.4400 2502.8000 1499.4600 2505.0000 ;
      RECT 1071.2200 2502.8000 1279.2400 2505.0000 ;
      RECT 0.0000 2502.8000 1062.9600 2503.5600 ;
      RECT 0.0000 2501.9200 3370.4200 2502.8000 ;
      RECT 3368.7200 2500.8400 3370.4200 2501.9200 ;
      RECT 3305.0200 2500.8400 3365.1200 2501.9200 ;
      RECT 2497.4200 2500.8400 3302.8200 2501.9200 ;
      RECT 2446.4800 2500.8400 2495.2200 2501.9200 ;
      RECT 2436.3200 2500.8400 2444.2800 2501.9200 ;
      RECT 2398.9000 2500.8400 2434.1200 2501.9200 ;
      RECT 2386.3400 2500.8400 2396.7000 2501.9200 ;
      RECT 1065.1600 2500.8400 2384.1400 2501.9200 ;
      RECT 1055.1000 2500.8400 1062.9600 2501.9200 ;
      RECT 1017.4800 2500.8400 1052.9000 2501.9200 ;
      RECT 1007.4200 2500.8400 1015.2800 2501.9200 ;
      RECT 5.3000 2500.8400 1005.2200 2501.9200 ;
      RECT 0.0000 2500.8400 1.7000 2501.9200 ;
      RECT 0.0000 2499.2000 3370.4200 2500.8400 ;
      RECT 3364.7200 2498.1200 3370.4200 2499.2000 ;
      RECT 3307.6200 2498.1200 3361.1200 2499.2000 ;
      RECT 2494.8200 2498.1200 3305.4200 2499.2000 ;
      RECT 2449.0800 2498.1200 2492.6200 2499.2000 ;
      RECT 2438.9200 2498.1200 2446.8800 2499.2000 ;
      RECT 2388.9400 2498.1200 2436.7200 2499.2000 ;
      RECT 1067.7600 2498.1200 2386.7400 2499.2000 ;
      RECT 1057.5000 2498.1200 1065.5600 2499.2000 ;
      RECT 1015.0800 2498.1200 1055.3000 2499.2000 ;
      RECT 1004.8200 2498.1200 1012.8800 2499.2000 ;
      RECT 9.3000 2498.1200 1002.6200 2499.2000 ;
      RECT 0.0000 2498.1200 5.7000 2499.2000 ;
      RECT 0.0000 2496.8400 3370.4200 2498.1200 ;
      RECT 1.1000 2496.4800 3370.4200 2496.8400 ;
      RECT 1.1000 2495.9400 1.7000 2496.4800 ;
      RECT 3368.7200 2495.4000 3370.4200 2496.4800 ;
      RECT 3305.0200 2495.4000 3365.1200 2496.4800 ;
      RECT 2497.4200 2495.4000 3302.8200 2496.4800 ;
      RECT 2446.4800 2495.4000 2495.2200 2496.4800 ;
      RECT 2436.3200 2495.4000 2444.2800 2496.4800 ;
      RECT 2398.9000 2495.4000 2434.1200 2496.4800 ;
      RECT 2386.3400 2495.4000 2396.7000 2496.4800 ;
      RECT 1065.1600 2495.4000 2384.1400 2496.4800 ;
      RECT 1055.1000 2495.4000 1062.9600 2496.4800 ;
      RECT 1017.4800 2495.4000 1052.9000 2496.4800 ;
      RECT 1007.4200 2495.4000 1015.2800 2496.4800 ;
      RECT 5.3000 2495.4000 1005.2200 2496.4800 ;
      RECT 0.0000 2495.4000 1.7000 2495.9400 ;
      RECT 0.0000 2493.7600 3370.4200 2495.4000 ;
      RECT 3364.7200 2492.6800 3370.4200 2493.7600 ;
      RECT 3307.6200 2492.6800 3361.1200 2493.7600 ;
      RECT 2494.8200 2492.6800 3305.4200 2493.7600 ;
      RECT 2449.0800 2492.6800 2492.6200 2493.7600 ;
      RECT 2438.9200 2492.6800 2446.8800 2493.7600 ;
      RECT 2388.9400 2492.6800 2436.7200 2493.7600 ;
      RECT 1067.7600 2492.6800 2386.7400 2493.7600 ;
      RECT 1057.5000 2492.6800 1065.5600 2493.7600 ;
      RECT 1015.0800 2492.6800 1055.3000 2493.7600 ;
      RECT 1004.8200 2492.6800 1012.8800 2493.7600 ;
      RECT 9.3000 2492.6800 1002.6200 2493.7600 ;
      RECT 0.0000 2492.6800 5.7000 2493.7600 ;
      RECT 0.0000 2491.0400 3370.4200 2492.6800 ;
      RECT 1065.1600 2490.0000 2384.1400 2491.0400 ;
      RECT 3368.7200 2489.9600 3370.4200 2491.0400 ;
      RECT 3305.0200 2489.9600 3365.1200 2491.0400 ;
      RECT 2497.4200 2489.9600 3302.8200 2491.0400 ;
      RECT 2446.4800 2489.9600 2495.2200 2491.0400 ;
      RECT 2436.3200 2489.9600 2444.2800 2491.0400 ;
      RECT 2398.9000 2489.9600 2434.1200 2491.0400 ;
      RECT 2386.3400 2489.9600 2396.7000 2491.0400 ;
      RECT 2176.1800 2489.9600 2384.1400 2490.0000 ;
      RECT 1065.1600 2489.9600 1072.8800 2490.0000 ;
      RECT 1055.1000 2489.9600 1062.9600 2491.0400 ;
      RECT 1017.4800 2489.9600 1052.9000 2491.0400 ;
      RECT 1007.4200 2489.9600 1015.2800 2491.0400 ;
      RECT 5.3000 2489.9600 1005.2200 2491.0400 ;
      RECT 0.0000 2489.9600 1.7000 2491.0400 ;
      RECT 2176.1800 2488.9200 3370.4200 2489.9600 ;
      RECT 1955.9600 2488.9200 2173.9800 2490.0000 ;
      RECT 1735.7400 2488.9200 1953.7600 2490.0000 ;
      RECT 1515.5200 2488.9200 1733.5400 2490.0000 ;
      RECT 1295.3000 2488.9200 1513.3200 2490.0000 ;
      RECT 1075.0800 2488.9200 1293.1000 2490.0000 ;
      RECT 0.0000 2488.9200 1072.8800 2489.9600 ;
      RECT 0.0000 2488.3200 3370.4200 2488.9200 ;
      RECT 1067.7600 2487.2800 2386.7400 2488.3200 ;
      RECT 3364.7200 2487.2400 3370.4200 2488.3200 ;
      RECT 3307.6200 2487.2400 3361.1200 2488.3200 ;
      RECT 2494.8200 2487.2400 3305.4200 2488.3200 ;
      RECT 2449.0800 2487.2400 2492.6200 2488.3200 ;
      RECT 2438.9200 2487.2400 2446.8800 2488.3200 ;
      RECT 2388.9400 2487.2400 2436.7200 2488.3200 ;
      RECT 2376.2800 2487.2400 2386.7400 2487.2800 ;
      RECT 1067.7600 2487.2400 1272.9800 2487.2800 ;
      RECT 1057.5000 2487.2400 1065.5600 2488.3200 ;
      RECT 1015.0800 2487.2400 1055.3000 2488.3200 ;
      RECT 1004.8200 2487.2400 1012.8800 2488.3200 ;
      RECT 9.3000 2487.2400 1002.6200 2488.3200 ;
      RECT 0.0000 2487.2400 5.7000 2488.3200 ;
      RECT 2376.2800 2486.2000 3370.4200 2487.2400 ;
      RECT 2156.0600 2486.2000 2374.0800 2487.2800 ;
      RECT 1935.8400 2486.2000 2153.8600 2487.2800 ;
      RECT 1715.6200 2486.2000 1933.6400 2487.2800 ;
      RECT 1495.4000 2486.2000 1713.4200 2487.2800 ;
      RECT 1275.1800 2486.2000 1493.2000 2487.2800 ;
      RECT 0.0000 2486.2000 1272.9800 2487.2400 ;
      RECT 0.0000 2485.8600 3370.4200 2486.2000 ;
      RECT 1.1000 2485.6000 3370.4200 2485.8600 ;
      RECT 1065.1600 2485.4700 2384.1400 2485.6000 ;
      RECT 1.1000 2484.9600 1.7000 2485.6000 ;
      RECT 3368.7200 2484.5200 3370.4200 2485.6000 ;
      RECT 3305.0200 2484.5200 3365.1200 2485.6000 ;
      RECT 2497.4200 2484.5200 3302.8200 2485.6000 ;
      RECT 2446.4800 2484.5200 2495.2200 2485.6000 ;
      RECT 2436.3200 2484.5200 2444.2800 2485.6000 ;
      RECT 2398.9000 2484.5200 2434.1200 2485.6000 ;
      RECT 2386.3400 2484.5200 2396.7000 2485.6000 ;
      RECT 1055.1000 2484.5200 1062.9600 2485.6000 ;
      RECT 1017.4800 2484.5200 1052.9000 2485.6000 ;
      RECT 1007.4200 2484.5200 1015.2800 2485.6000 ;
      RECT 5.3000 2484.5200 1005.2200 2485.6000 ;
      RECT 0.0000 2484.5200 1.7000 2484.9600 ;
      RECT 2386.3400 2483.2700 3370.4200 2484.5200 ;
      RECT 2172.3200 2483.2700 2380.3400 2485.4700 ;
      RECT 1952.1000 2483.2700 2160.1200 2485.4700 ;
      RECT 1731.8800 2483.2700 1939.9000 2485.4700 ;
      RECT 1511.6600 2483.2700 1719.6800 2485.4700 ;
      RECT 1291.4400 2483.2700 1499.4600 2485.4700 ;
      RECT 1071.2200 2483.2700 1279.2400 2485.4700 ;
      RECT 0.0000 2483.2700 1062.9600 2484.5200 ;
      RECT 0.0000 2483.0700 3370.4200 2483.2700 ;
      RECT 2172.3200 2482.8800 3370.4200 2483.0700 ;
      RECT 0.0000 2482.8800 1065.5600 2483.0700 ;
      RECT 3364.7200 2481.8000 3370.4200 2482.8800 ;
      RECT 3307.6200 2481.8000 3361.1200 2482.8800 ;
      RECT 2494.8200 2481.8000 3305.4200 2482.8800 ;
      RECT 2449.0800 2481.8000 2492.6200 2482.8800 ;
      RECT 2438.9200 2481.8000 2446.8800 2482.8800 ;
      RECT 2388.9400 2481.8000 2436.7200 2482.8800 ;
      RECT 2172.3200 2481.8000 2386.7400 2482.8800 ;
      RECT 1057.5000 2481.8000 1065.5600 2482.8800 ;
      RECT 1015.0800 2481.8000 1055.3000 2482.8800 ;
      RECT 1004.8200 2481.8000 1012.8800 2482.8800 ;
      RECT 9.3000 2481.8000 1002.6200 2482.8800 ;
      RECT 0.0000 2481.8000 5.7000 2482.8800 ;
      RECT 2172.3200 2480.8700 3370.4200 2481.8000 ;
      RECT 1952.1000 2480.8700 2166.5200 2483.0700 ;
      RECT 1731.8800 2480.8700 1946.3000 2483.0700 ;
      RECT 1511.6600 2480.8700 1726.0800 2483.0700 ;
      RECT 1291.4400 2480.8700 1499.4600 2483.0700 ;
      RECT 1071.2200 2480.8700 1279.2400 2483.0700 ;
      RECT 0.0000 2480.8700 1065.5600 2481.8000 ;
      RECT 0.0000 2480.1600 3370.4200 2480.8700 ;
      RECT 3368.7200 2479.0800 3370.4200 2480.1600 ;
      RECT 3305.0200 2479.0800 3365.1200 2480.1600 ;
      RECT 2497.4200 2479.0800 3302.8200 2480.1600 ;
      RECT 2446.4800 2479.0800 2495.2200 2480.1600 ;
      RECT 2436.3200 2479.0800 2444.2800 2480.1600 ;
      RECT 2398.9000 2479.0800 2434.1200 2480.1600 ;
      RECT 2386.3400 2479.0800 2396.7000 2480.1600 ;
      RECT 1007.4200 2479.0800 2384.1400 2480.1600 ;
      RECT 5.3000 2479.0800 1005.2200 2480.1600 ;
      RECT 0.0000 2479.0800 1.7000 2480.1600 ;
      RECT 0.0000 2477.4400 3370.4200 2479.0800 ;
      RECT 1004.8200 2476.9000 2446.8800 2477.4400 ;
      RECT 3364.7200 2476.3600 3370.4200 2477.4400 ;
      RECT 3307.6200 2476.3600 3361.1200 2477.4400 ;
      RECT 2494.8200 2476.3600 3305.4200 2477.4400 ;
      RECT 2449.0800 2476.3600 2492.6200 2477.4400 ;
      RECT 2386.3400 2476.3600 2446.8800 2476.9000 ;
      RECT 1004.8200 2476.3600 1062.9600 2476.9000 ;
      RECT 9.3000 2476.3600 1002.6200 2477.4400 ;
      RECT 0.0000 2476.3600 5.7000 2477.4400 ;
      RECT 0.0000 2475.4900 1062.9600 2476.3600 ;
      RECT 2386.3400 2474.7200 3370.4200 2476.3600 ;
      RECT 1.1000 2474.7200 1062.9600 2475.4900 ;
      RECT 2386.3400 2474.7000 2444.2800 2474.7200 ;
      RECT 1007.4200 2474.7000 1062.9600 2474.7200 ;
      RECT 1.1000 2474.5900 1.7000 2474.7200 ;
      RECT 1007.4200 2474.4000 2444.2800 2474.7000 ;
      RECT 1945.8000 2474.3000 2444.2800 2474.4000 ;
      RECT 1007.4200 2474.3000 1943.4000 2474.4000 ;
      RECT 3368.7200 2473.6400 3370.4200 2474.7200 ;
      RECT 3305.0200 2473.6400 3365.1200 2474.7200 ;
      RECT 2497.4200 2473.6400 3302.8200 2474.7200 ;
      RECT 2446.4800 2473.6400 2495.2200 2474.7200 ;
      RECT 2388.9400 2473.6400 2444.2800 2474.3000 ;
      RECT 1007.4200 2473.6400 1065.5600 2474.3000 ;
      RECT 5.3000 2473.6400 1005.2200 2474.7200 ;
      RECT 0.0000 2473.6400 1.7000 2474.5900 ;
      RECT 2388.9400 2472.1000 3370.4200 2473.6400 ;
      RECT 0.0000 2472.1000 1065.5600 2473.6400 ;
      RECT 1945.8000 2472.0000 3370.4200 2472.1000 ;
      RECT 0.0000 2472.0000 1943.4000 2472.1000 ;
      RECT 3364.7200 2470.9200 3370.4200 2472.0000 ;
      RECT 3307.6200 2470.9200 3361.1200 2472.0000 ;
      RECT 2494.8200 2470.9200 3305.4200 2472.0000 ;
      RECT 2449.0800 2470.9200 2492.6200 2472.0000 ;
      RECT 1945.8000 2470.9200 2446.8800 2472.0000 ;
      RECT 1004.8200 2470.9200 1943.4000 2472.0000 ;
      RECT 9.3000 2470.9200 1002.6200 2472.0000 ;
      RECT 0.0000 2470.9200 5.7000 2472.0000 ;
      RECT 1945.8000 2470.4000 3370.4200 2470.9200 ;
      RECT 0.0000 2470.4000 1943.4000 2470.9200 ;
      RECT 0.0000 2469.2800 3370.4200 2470.4000 ;
      RECT 3368.7200 2468.2000 3370.4200 2469.2800 ;
      RECT 3305.0200 2468.2000 3365.1200 2469.2800 ;
      RECT 2497.4200 2468.2000 3302.8200 2469.2800 ;
      RECT 2446.4800 2468.2000 2495.2200 2469.2800 ;
      RECT 1007.4200 2468.2000 2444.2800 2469.2800 ;
      RECT 5.3000 2468.2000 1005.2200 2469.2800 ;
      RECT 0.0000 2468.2000 1.7000 2469.2800 ;
      RECT 0.0000 2467.7000 3370.4200 2468.2000 ;
      RECT 1287.9800 2467.4400 3370.4200 2467.7000 ;
      RECT 2168.7200 2466.5600 3370.4200 2467.4400 ;
      RECT 0.0000 2466.5600 1065.5600 2467.7000 ;
      RECT 1004.8200 2466.5500 1065.5600 2466.5600 ;
      RECT 2168.7200 2466.3900 2446.8800 2466.5600 ;
      RECT 1287.9800 2466.3900 1946.3000 2467.4400 ;
      RECT 1071.3600 2465.5000 1279.3800 2467.7000 ;
      RECT 1062.4600 2465.5000 1065.5600 2466.5500 ;
      RECT 3364.7200 2465.4800 3370.4200 2466.5600 ;
      RECT 3307.6200 2465.4800 3361.1200 2466.5600 ;
      RECT 2494.8200 2465.4800 3305.4200 2466.5600 ;
      RECT 2449.0800 2465.4800 2492.6200 2466.5600 ;
      RECT 9.3000 2465.4800 1002.6200 2466.5600 ;
      RECT 0.0000 2465.4800 5.7000 2466.5600 ;
      RECT 1952.1000 2465.2400 2160.1200 2467.4400 ;
      RECT 1943.2000 2465.2400 1946.3000 2466.3900 ;
      RECT 1062.4600 2465.1000 1285.6400 2465.5000 ;
      RECT 1943.2000 2464.8400 2166.5200 2465.2400 ;
      RECT 0.0000 2464.5100 1002.6200 2465.4800 ;
      RECT 1062.4600 2464.3500 1062.9600 2465.1000 ;
      RECT 1011.2200 2464.3500 1059.1600 2466.5500 ;
      RECT 1.1000 2464.3500 1002.6200 2464.5100 ;
      RECT 2449.0800 2464.1900 3370.4200 2465.4800 ;
      RECT 2392.5400 2464.1900 2440.4800 2466.3900 ;
      RECT 2172.3200 2464.1900 2380.3400 2466.3900 ;
      RECT 2166.1200 2464.1900 2166.5200 2464.8400 ;
      RECT 1943.2000 2464.1900 1943.7000 2464.8400 ;
      RECT 1731.8800 2464.1900 1939.9000 2466.3900 ;
      RECT 1511.6600 2464.1900 1719.6800 2466.3900 ;
      RECT 1291.4400 2464.1900 1499.4600 2466.3900 ;
      RECT 1285.3800 2464.1900 1285.6400 2465.1000 ;
      RECT 1.1000 2464.1500 1062.9600 2464.3500 ;
      RECT 2166.1200 2463.8400 3370.4200 2464.1900 ;
      RECT 1.1000 2463.8400 1005.2200 2464.1500 ;
      RECT 2166.1200 2463.7900 2444.2800 2463.8400 ;
      RECT 1285.3800 2463.7900 1943.7000 2464.1900 ;
      RECT 1.1000 2463.6100 1.7000 2463.8400 ;
      RECT 1071.3600 2462.9000 1279.3800 2465.1000 ;
      RECT 3368.7200 2462.7600 3370.4200 2463.8400 ;
      RECT 3305.0200 2462.7600 3365.1200 2463.8400 ;
      RECT 2497.4200 2462.7600 3302.8200 2463.8400 ;
      RECT 2446.4800 2462.7600 2495.2200 2463.8400 ;
      RECT 5.3000 2462.7600 1005.2200 2463.8400 ;
      RECT 0.0000 2462.7600 1.7000 2463.6100 ;
      RECT 1952.1000 2462.6400 2160.1200 2464.8400 ;
      RECT 1065.1600 2461.9500 1283.0400 2462.9000 ;
      RECT 1011.2200 2461.9500 1059.1600 2464.1500 ;
      RECT 0.0000 2461.9500 1005.2200 2462.7600 ;
      RECT 2446.4800 2461.5900 3370.4200 2462.7600 ;
      RECT 2392.5400 2461.5900 2440.4800 2463.7900 ;
      RECT 2172.3200 2461.5900 2380.3400 2463.7900 ;
      RECT 1945.9000 2461.5900 2163.9200 2462.6400 ;
      RECT 1731.8800 2461.5900 1939.9000 2463.7900 ;
      RECT 1511.6600 2461.5900 1719.6800 2463.7900 ;
      RECT 1291.4400 2461.5900 1499.4600 2463.7900 ;
      RECT 0.0000 2461.5900 1283.0400 2461.9500 ;
      RECT 0.0000 2461.1200 3370.4200 2461.5900 ;
      RECT 3364.7200 2460.0400 3370.4200 2461.1200 ;
      RECT 3307.6200 2460.0400 3361.1200 2461.1200 ;
      RECT 2494.8200 2460.0400 3305.4200 2461.1200 ;
      RECT 2449.0800 2460.0400 2492.6200 2461.1200 ;
      RECT 1004.8200 2460.0400 2446.8800 2461.1200 ;
      RECT 9.3000 2460.0400 1002.6200 2461.1200 ;
      RECT 0.0000 2460.0400 5.7000 2461.1200 ;
      RECT 0.0000 2458.9200 3370.4200 2460.0400 ;
      RECT 2183.2400 2458.4000 3370.4200 2458.9200 ;
      RECT 0.0000 2458.4000 1300.1600 2458.9200 ;
      RECT 1007.4200 2458.0200 1300.1600 2458.4000 ;
      RECT 2183.2400 2457.8400 2444.2800 2458.4000 ;
      RECT 1742.8000 2457.8400 2181.0400 2458.9200 ;
      RECT 1522.5800 2457.8400 1740.6000 2458.9200 ;
      RECT 1302.3600 2457.8400 1520.3800 2458.9200 ;
      RECT 1075.1200 2457.8400 1300.1600 2458.0200 ;
      RECT 1075.1200 2457.7600 2444.2800 2457.8400 ;
      RECT 3368.7200 2457.3200 3370.4200 2458.4000 ;
      RECT 3305.0200 2457.3200 3365.1200 2458.4000 ;
      RECT 2497.4200 2457.3200 3302.8200 2458.4000 ;
      RECT 2446.4800 2457.3200 2495.2200 2458.4000 ;
      RECT 1955.8600 2457.3200 2444.2800 2457.7600 ;
      RECT 1007.4200 2457.3200 1072.9200 2458.0200 ;
      RECT 5.3000 2457.3200 1005.2200 2458.4000 ;
      RECT 0.0000 2457.3200 1.7000 2458.4000 ;
      RECT 1075.1200 2456.9400 1953.6600 2457.7600 ;
      RECT 0.0000 2456.9400 1072.9200 2457.3200 ;
      RECT 1955.8600 2456.6800 3370.4200 2457.3200 ;
      RECT 0.0000 2456.6800 1953.6600 2456.9400 ;
      RECT 0.0000 2455.6800 3370.4200 2456.6800 ;
      RECT 3364.7200 2454.6000 3370.4200 2455.6800 ;
      RECT 3307.6200 2454.6000 3361.1200 2455.6800 ;
      RECT 2494.8200 2454.6000 3305.4200 2455.6800 ;
      RECT 2449.0800 2454.6000 2492.6200 2455.6800 ;
      RECT 1004.8200 2454.6000 2446.8800 2455.6800 ;
      RECT 9.3000 2454.6000 1002.6200 2455.6800 ;
      RECT 0.0000 2454.6000 5.7000 2455.6800 ;
      RECT 0.0000 2453.5300 3370.4200 2454.6000 ;
      RECT 1.1000 2452.9600 3370.4200 2453.5300 ;
      RECT 1.1000 2452.6300 1.7000 2452.9600 ;
      RECT 3368.7200 2451.8800 3370.4200 2452.9600 ;
      RECT 3305.0200 2451.8800 3365.1200 2452.9600 ;
      RECT 2497.4200 2451.8800 3302.8200 2452.9600 ;
      RECT 2446.4800 2451.8800 2495.2200 2452.9600 ;
      RECT 1007.4200 2451.8800 2444.2800 2452.9600 ;
      RECT 5.3000 2451.8800 1005.2200 2452.9600 ;
      RECT 0.0000 2451.8800 1.7000 2452.6300 ;
      RECT 0.0000 2450.2400 3370.4200 2451.8800 ;
      RECT 3364.7200 2449.1600 3370.4200 2450.2400 ;
      RECT 3307.6200 2449.1600 3361.1200 2450.2400 ;
      RECT 2494.8200 2449.1600 3305.4200 2450.2400 ;
      RECT 2449.0800 2449.1600 2492.6200 2450.2400 ;
      RECT 1004.8200 2449.1600 2446.8800 2450.2400 ;
      RECT 9.3000 2449.1600 1002.6200 2450.2400 ;
      RECT 0.0000 2449.1600 5.7000 2450.2400 ;
      RECT 0.0000 2447.5200 3370.4200 2449.1600 ;
      RECT 3368.7200 2446.4400 3370.4200 2447.5200 ;
      RECT 3305.0200 2446.4400 3365.1200 2447.5200 ;
      RECT 2497.4200 2446.4400 3302.8200 2447.5200 ;
      RECT 2446.4800 2446.4400 2495.2200 2447.5200 ;
      RECT 1007.4200 2446.4400 2444.2800 2447.5200 ;
      RECT 5.3000 2446.4400 1005.2200 2447.5200 ;
      RECT 0.0000 2446.4400 1.7000 2447.5200 ;
      RECT 0.0000 2444.8000 3370.4200 2446.4400 ;
      RECT 3364.7200 2443.7200 3370.4200 2444.8000 ;
      RECT 3307.6200 2443.7200 3361.1200 2444.8000 ;
      RECT 2494.8200 2443.7200 3305.4200 2444.8000 ;
      RECT 2449.0800 2443.7200 2492.6200 2444.8000 ;
      RECT 1004.8200 2443.7200 2446.8800 2444.8000 ;
      RECT 9.3000 2443.7200 1002.6200 2444.8000 ;
      RECT 0.0000 2443.7200 5.7000 2444.8000 ;
      RECT 0.0000 2442.5500 3370.4200 2443.7200 ;
      RECT 1.1000 2442.0800 3370.4200 2442.5500 ;
      RECT 1.1000 2441.6500 1.7000 2442.0800 ;
      RECT 3368.7200 2441.0000 3370.4200 2442.0800 ;
      RECT 3305.0200 2441.0000 3365.1200 2442.0800 ;
      RECT 2497.4200 2441.0000 3302.8200 2442.0800 ;
      RECT 2446.4800 2441.0000 2495.2200 2442.0800 ;
      RECT 1007.4200 2441.0000 2444.2800 2442.0800 ;
      RECT 5.3000 2441.0000 1005.2200 2442.0800 ;
      RECT 0.0000 2441.0000 1.7000 2441.6500 ;
      RECT 0.0000 2439.3600 3370.4200 2441.0000 ;
      RECT 3364.7200 2438.2800 3370.4200 2439.3600 ;
      RECT 3307.6200 2438.2800 3361.1200 2439.3600 ;
      RECT 2494.8200 2438.2800 3305.4200 2439.3600 ;
      RECT 2449.0800 2438.2800 2492.6200 2439.3600 ;
      RECT 1004.8200 2438.2800 2446.8800 2439.3600 ;
      RECT 9.3000 2438.2800 1002.6200 2439.3600 ;
      RECT 0.0000 2438.2800 5.7000 2439.3600 ;
      RECT 0.0000 2436.6400 3370.4200 2438.2800 ;
      RECT 3368.7200 2435.5600 3370.4200 2436.6400 ;
      RECT 3305.0200 2435.5600 3365.1200 2436.6400 ;
      RECT 2497.4200 2435.5600 3302.8200 2436.6400 ;
      RECT 2446.4800 2435.5600 2495.2200 2436.6400 ;
      RECT 1007.4200 2435.5600 2444.2800 2436.6400 ;
      RECT 5.3000 2435.5600 1005.2200 2436.6400 ;
      RECT 0.0000 2435.5600 1.7000 2436.6400 ;
      RECT 0.0000 2433.9200 3370.4200 2435.5600 ;
      RECT 3364.7200 2432.8400 3370.4200 2433.9200 ;
      RECT 3307.6200 2432.8400 3361.1200 2433.9200 ;
      RECT 2494.8200 2432.8400 3305.4200 2433.9200 ;
      RECT 2449.0800 2432.8400 2492.6200 2433.9200 ;
      RECT 1004.8200 2432.8400 2446.8800 2433.9200 ;
      RECT 9.3000 2432.8400 1002.6200 2433.9200 ;
      RECT 0.0000 2432.8400 5.7000 2433.9200 ;
      RECT 0.0000 2431.5700 3370.4200 2432.8400 ;
      RECT 1.1000 2431.2000 3370.4200 2431.5700 ;
      RECT 1.1000 2430.6700 1.7000 2431.2000 ;
      RECT 3368.7200 2430.1200 3370.4200 2431.2000 ;
      RECT 3305.0200 2430.1200 3365.1200 2431.2000 ;
      RECT 2497.4200 2430.1200 3302.8200 2431.2000 ;
      RECT 2446.4800 2430.1200 2495.2200 2431.2000 ;
      RECT 1007.4200 2430.1200 2444.2800 2431.2000 ;
      RECT 5.3000 2430.1200 1005.2200 2431.2000 ;
      RECT 0.0000 2430.1200 1.7000 2430.6700 ;
      RECT 0.0000 2428.4800 3370.4200 2430.1200 ;
      RECT 3364.7200 2427.4000 3370.4200 2428.4800 ;
      RECT 3307.6200 2427.4000 3361.1200 2428.4800 ;
      RECT 2494.8200 2427.4000 3305.4200 2428.4800 ;
      RECT 2449.0800 2427.4000 2492.6200 2428.4800 ;
      RECT 1004.8200 2427.4000 2446.8800 2428.4800 ;
      RECT 9.3000 2427.4000 1002.6200 2428.4800 ;
      RECT 0.0000 2427.4000 5.7000 2428.4800 ;
      RECT 0.0000 2425.7600 3370.4200 2427.4000 ;
      RECT 3368.7200 2424.6800 3370.4200 2425.7600 ;
      RECT 3305.0200 2424.6800 3365.1200 2425.7600 ;
      RECT 2497.4200 2424.6800 3302.8200 2425.7600 ;
      RECT 2446.4800 2424.6800 2495.2200 2425.7600 ;
      RECT 1007.4200 2424.6800 2444.2800 2425.7600 ;
      RECT 5.3000 2424.6800 1005.2200 2425.7600 ;
      RECT 0.0000 2424.6800 1.7000 2425.7600 ;
      RECT 0.0000 2423.0400 3370.4200 2424.6800 ;
      RECT 3364.7200 2421.9600 3370.4200 2423.0400 ;
      RECT 3307.6200 2421.9600 3361.1200 2423.0400 ;
      RECT 2494.8200 2421.9600 3305.4200 2423.0400 ;
      RECT 2449.0800 2421.9600 2492.6200 2423.0400 ;
      RECT 1004.8200 2421.9600 2446.8800 2423.0400 ;
      RECT 9.3000 2421.9600 1002.6200 2423.0400 ;
      RECT 0.0000 2421.9600 5.7000 2423.0400 ;
      RECT 0.0000 2421.2000 3370.4200 2421.9600 ;
      RECT 1.1000 2420.3200 3370.4200 2421.2000 ;
      RECT 1.1000 2420.3000 1.7000 2420.3200 ;
      RECT 3368.7200 2419.2400 3370.4200 2420.3200 ;
      RECT 3305.0200 2419.2400 3365.1200 2420.3200 ;
      RECT 2497.4200 2419.2400 3302.8200 2420.3200 ;
      RECT 2446.4800 2419.2400 2495.2200 2420.3200 ;
      RECT 1007.4200 2419.2400 2444.2800 2420.3200 ;
      RECT 5.3000 2419.2400 1005.2200 2420.3200 ;
      RECT 0.0000 2419.2400 1.7000 2420.3000 ;
      RECT 0.0000 2417.6000 3370.4200 2419.2400 ;
      RECT 3364.7200 2416.5200 3370.4200 2417.6000 ;
      RECT 3307.6200 2416.5200 3361.1200 2417.6000 ;
      RECT 2494.8200 2416.5200 3305.4200 2417.6000 ;
      RECT 2449.0800 2416.5200 2492.6200 2417.6000 ;
      RECT 1004.8200 2416.5200 2446.8800 2417.6000 ;
      RECT 9.3000 2416.5200 1002.6200 2417.6000 ;
      RECT 0.0000 2416.5200 5.7000 2417.6000 ;
      RECT 0.0000 2414.8800 3370.4200 2416.5200 ;
      RECT 3368.7200 2413.8000 3370.4200 2414.8800 ;
      RECT 3305.0200 2413.8000 3365.1200 2414.8800 ;
      RECT 2497.4200 2413.8000 3302.8200 2414.8800 ;
      RECT 2446.4800 2413.8000 2495.2200 2414.8800 ;
      RECT 1007.4200 2413.8000 2444.2800 2414.8800 ;
      RECT 5.3000 2413.8000 1005.2200 2414.8800 ;
      RECT 0.0000 2413.8000 1.7000 2414.8800 ;
      RECT 0.0000 2412.1600 3370.4200 2413.8000 ;
      RECT 3364.7200 2411.0800 3370.4200 2412.1600 ;
      RECT 3307.6200 2411.0800 3361.1200 2412.1600 ;
      RECT 2494.8200 2411.0800 3305.4200 2412.1600 ;
      RECT 2449.0800 2411.0800 2492.6200 2412.1600 ;
      RECT 1004.8200 2411.0800 2446.8800 2412.1600 ;
      RECT 9.3000 2411.0800 1002.6200 2412.1600 ;
      RECT 0.0000 2411.0800 5.7000 2412.1600 ;
      RECT 0.0000 2410.2200 3370.4200 2411.0800 ;
      RECT 1.1000 2409.4400 3370.4200 2410.2200 ;
      RECT 1.1000 2409.3200 1.7000 2409.4400 ;
      RECT 3368.7200 2408.3600 3370.4200 2409.4400 ;
      RECT 3305.0200 2408.3600 3365.1200 2409.4400 ;
      RECT 2497.4200 2408.3600 3302.8200 2409.4400 ;
      RECT 2446.4800 2408.3600 2495.2200 2409.4400 ;
      RECT 1007.4200 2408.3600 2444.2800 2409.4400 ;
      RECT 5.3000 2408.3600 1005.2200 2409.4400 ;
      RECT 0.0000 2408.3600 1.7000 2409.3200 ;
      RECT 0.0000 2406.7200 3370.4200 2408.3600 ;
      RECT 3364.7200 2405.6400 3370.4200 2406.7200 ;
      RECT 3307.6200 2405.6400 3361.1200 2406.7200 ;
      RECT 2494.8200 2405.6400 3305.4200 2406.7200 ;
      RECT 2449.0800 2405.6400 2492.6200 2406.7200 ;
      RECT 1004.8200 2405.6400 2446.8800 2406.7200 ;
      RECT 9.3000 2405.6400 1002.6200 2406.7200 ;
      RECT 0.0000 2405.6400 5.7000 2406.7200 ;
      RECT 0.0000 2404.0000 3370.4200 2405.6400 ;
      RECT 3368.7200 2402.9200 3370.4200 2404.0000 ;
      RECT 3305.0200 2402.9200 3365.1200 2404.0000 ;
      RECT 2497.4200 2402.9200 3302.8200 2404.0000 ;
      RECT 2446.4800 2402.9200 2495.2200 2404.0000 ;
      RECT 1007.4200 2402.9200 2444.2800 2404.0000 ;
      RECT 5.3000 2402.9200 1005.2200 2404.0000 ;
      RECT 0.0000 2402.9200 1.7000 2404.0000 ;
      RECT 0.0000 2401.2800 3370.4200 2402.9200 ;
      RECT 3364.7200 2400.2000 3370.4200 2401.2800 ;
      RECT 3307.6200 2400.2000 3361.1200 2401.2800 ;
      RECT 2494.8200 2400.2000 3305.4200 2401.2800 ;
      RECT 2449.0800 2400.2000 2492.6200 2401.2800 ;
      RECT 1004.8200 2400.2000 2446.8800 2401.2800 ;
      RECT 9.3000 2400.2000 1002.6200 2401.2800 ;
      RECT 0.0000 2400.2000 5.7000 2401.2800 ;
      RECT 0.0000 2399.2400 3370.4200 2400.2000 ;
      RECT 1.1000 2398.5600 3370.4200 2399.2400 ;
      RECT 1.1000 2398.3400 1.7000 2398.5600 ;
      RECT 3368.7200 2397.4800 3370.4200 2398.5600 ;
      RECT 3305.0200 2397.4800 3365.1200 2398.5600 ;
      RECT 2497.4200 2397.4800 3302.8200 2398.5600 ;
      RECT 2446.4800 2397.4800 2495.2200 2398.5600 ;
      RECT 1007.4200 2397.4800 2444.2800 2398.5600 ;
      RECT 5.3000 2397.4800 1005.2200 2398.5600 ;
      RECT 0.0000 2397.4800 1.7000 2398.3400 ;
      RECT 0.0000 2395.8400 3370.4200 2397.4800 ;
      RECT 3364.7200 2394.7600 3370.4200 2395.8400 ;
      RECT 3307.6200 2394.7600 3361.1200 2395.8400 ;
      RECT 2494.8200 2394.7600 3305.4200 2395.8400 ;
      RECT 2449.0800 2394.7600 2492.6200 2395.8400 ;
      RECT 1004.8200 2394.7600 2446.8800 2395.8400 ;
      RECT 9.3000 2394.7600 1002.6200 2395.8400 ;
      RECT 0.0000 2394.7600 5.7000 2395.8400 ;
      RECT 0.0000 2393.1200 3370.4200 2394.7600 ;
      RECT 3368.7200 2392.0400 3370.4200 2393.1200 ;
      RECT 3305.0200 2392.0400 3365.1200 2393.1200 ;
      RECT 2497.4200 2392.0400 3302.8200 2393.1200 ;
      RECT 2446.4800 2392.0400 2495.2200 2393.1200 ;
      RECT 1007.4200 2392.0400 2444.2800 2393.1200 ;
      RECT 5.3000 2392.0400 1005.2200 2393.1200 ;
      RECT 0.0000 2392.0400 1.7000 2393.1200 ;
      RECT 0.0000 2390.4000 3370.4200 2392.0400 ;
      RECT 3364.7200 2389.3200 3370.4200 2390.4000 ;
      RECT 3307.6200 2389.3200 3361.1200 2390.4000 ;
      RECT 2494.8200 2389.3200 3305.4200 2390.4000 ;
      RECT 2449.0800 2389.3200 2492.6200 2390.4000 ;
      RECT 1004.8200 2389.3200 2446.8800 2390.4000 ;
      RECT 9.3000 2389.3200 1002.6200 2390.4000 ;
      RECT 0.0000 2389.3200 5.7000 2390.4000 ;
      RECT 0.0000 2388.2600 3370.4200 2389.3200 ;
      RECT 1.1000 2387.6800 3370.4200 2388.2600 ;
      RECT 1.1000 2387.3600 1.7000 2387.6800 ;
      RECT 3368.7200 2386.6000 3370.4200 2387.6800 ;
      RECT 3305.0200 2386.6000 3365.1200 2387.6800 ;
      RECT 2497.4200 2386.6000 3302.8200 2387.6800 ;
      RECT 2446.4800 2386.6000 2495.2200 2387.6800 ;
      RECT 1007.4200 2386.6000 2444.2800 2387.6800 ;
      RECT 5.3000 2386.6000 1005.2200 2387.6800 ;
      RECT 0.0000 2386.6000 1.7000 2387.3600 ;
      RECT 0.0000 2384.9600 3370.4200 2386.6000 ;
      RECT 3364.7200 2383.8800 3370.4200 2384.9600 ;
      RECT 3307.6200 2383.8800 3361.1200 2384.9600 ;
      RECT 2494.8200 2383.8800 3305.4200 2384.9600 ;
      RECT 2449.0800 2383.8800 2492.6200 2384.9600 ;
      RECT 1004.8200 2383.8800 2446.8800 2384.9600 ;
      RECT 9.3000 2383.8800 1002.6200 2384.9600 ;
      RECT 0.0000 2383.8800 5.7000 2384.9600 ;
      RECT 0.0000 2382.2400 3370.4200 2383.8800 ;
      RECT 3368.7200 2381.1600 3370.4200 2382.2400 ;
      RECT 3305.0200 2381.1600 3365.1200 2382.2400 ;
      RECT 2497.4200 2381.1600 3302.8200 2382.2400 ;
      RECT 2446.4800 2381.1600 2495.2200 2382.2400 ;
      RECT 1007.4200 2381.1600 2444.2800 2382.2400 ;
      RECT 5.3000 2381.1600 1005.2200 2382.2400 ;
      RECT 0.0000 2381.1600 1.7000 2382.2400 ;
      RECT 0.0000 2379.5200 3370.4200 2381.1600 ;
      RECT 3364.7200 2378.4400 3370.4200 2379.5200 ;
      RECT 3307.6200 2378.4400 3361.1200 2379.5200 ;
      RECT 2494.8200 2378.4400 3305.4200 2379.5200 ;
      RECT 2449.0800 2378.4400 2492.6200 2379.5200 ;
      RECT 1004.8200 2378.4400 2446.8800 2379.5200 ;
      RECT 9.3000 2378.4400 1002.6200 2379.5200 ;
      RECT 0.0000 2378.4400 5.7000 2379.5200 ;
      RECT 0.0000 2377.2800 3370.4200 2378.4400 ;
      RECT 1.1000 2376.8000 3370.4200 2377.2800 ;
      RECT 1.1000 2376.3800 1.7000 2376.8000 ;
      RECT 3368.7200 2375.7200 3370.4200 2376.8000 ;
      RECT 3305.0200 2375.7200 3365.1200 2376.8000 ;
      RECT 2497.4200 2375.7200 3302.8200 2376.8000 ;
      RECT 2446.4800 2375.7200 2495.2200 2376.8000 ;
      RECT 1007.4200 2375.7200 2444.2800 2376.8000 ;
      RECT 5.3000 2375.7200 1005.2200 2376.8000 ;
      RECT 0.0000 2375.7200 1.7000 2376.3800 ;
      RECT 0.0000 2374.0800 3370.4200 2375.7200 ;
      RECT 3364.7200 2373.0000 3370.4200 2374.0800 ;
      RECT 3307.6200 2373.0000 3361.1200 2374.0800 ;
      RECT 2494.8200 2373.0000 3305.4200 2374.0800 ;
      RECT 2449.0800 2373.0000 2492.6200 2374.0800 ;
      RECT 1004.8200 2373.0000 2446.8800 2374.0800 ;
      RECT 9.3000 2373.0000 1002.6200 2374.0800 ;
      RECT 0.0000 2373.0000 5.7000 2374.0800 ;
      RECT 0.0000 2371.3600 3370.4200 2373.0000 ;
      RECT 3368.7200 2370.2800 3370.4200 2371.3600 ;
      RECT 3305.0200 2370.2800 3365.1200 2371.3600 ;
      RECT 2497.4200 2370.2800 3302.8200 2371.3600 ;
      RECT 2446.4800 2370.2800 2495.2200 2371.3600 ;
      RECT 1007.4200 2370.2800 2444.2800 2371.3600 ;
      RECT 5.3000 2370.2800 1005.2200 2371.3600 ;
      RECT 0.0000 2370.2800 1.7000 2371.3600 ;
      RECT 0.0000 2368.6400 3370.4200 2370.2800 ;
      RECT 3364.7200 2367.5600 3370.4200 2368.6400 ;
      RECT 3307.6200 2367.5600 3361.1200 2368.6400 ;
      RECT 2494.8200 2367.5600 3305.4200 2368.6400 ;
      RECT 2449.0800 2367.5600 2492.6200 2368.6400 ;
      RECT 1004.8200 2367.5600 2446.8800 2368.6400 ;
      RECT 9.3000 2367.5600 1002.6200 2368.6400 ;
      RECT 0.0000 2367.5600 5.7000 2368.6400 ;
      RECT 0.0000 2366.9100 3370.4200 2367.5600 ;
      RECT 1.1000 2366.0100 3370.4200 2366.9100 ;
      RECT 0.0000 2365.9200 3370.4200 2366.0100 ;
      RECT 3368.7200 2364.8400 3370.4200 2365.9200 ;
      RECT 3305.0200 2364.8400 3365.1200 2365.9200 ;
      RECT 2497.4200 2364.8400 3302.8200 2365.9200 ;
      RECT 2446.4800 2364.8400 2495.2200 2365.9200 ;
      RECT 1007.4200 2364.8400 2444.2800 2365.9200 ;
      RECT 5.3000 2364.8400 1005.2200 2365.9200 ;
      RECT 0.0000 2364.8400 1.7000 2365.9200 ;
      RECT 0.0000 2363.2000 3370.4200 2364.8400 ;
      RECT 3364.7200 2362.1200 3370.4200 2363.2000 ;
      RECT 3307.6200 2362.1200 3361.1200 2363.2000 ;
      RECT 2494.8200 2362.1200 3305.4200 2363.2000 ;
      RECT 2449.0800 2362.1200 2492.6200 2363.2000 ;
      RECT 1004.8200 2362.1200 2446.8800 2363.2000 ;
      RECT 9.3000 2362.1200 1002.6200 2363.2000 ;
      RECT 0.0000 2362.1200 5.7000 2363.2000 ;
      RECT 0.0000 2360.4800 3370.4200 2362.1200 ;
      RECT 3368.7200 2359.4000 3370.4200 2360.4800 ;
      RECT 3305.0200 2359.4000 3365.1200 2360.4800 ;
      RECT 2497.4200 2359.4000 3302.8200 2360.4800 ;
      RECT 2446.4800 2359.4000 2495.2200 2360.4800 ;
      RECT 1007.4200 2359.4000 2444.2800 2360.4800 ;
      RECT 5.3000 2359.4000 1005.2200 2360.4800 ;
      RECT 0.0000 2359.4000 1.7000 2360.4800 ;
      RECT 0.0000 2357.7600 3370.4200 2359.4000 ;
      RECT 3364.7200 2356.6800 3370.4200 2357.7600 ;
      RECT 3307.6200 2356.6800 3361.1200 2357.7600 ;
      RECT 2494.8200 2356.6800 3305.4200 2357.7600 ;
      RECT 2449.0800 2356.6800 2492.6200 2357.7600 ;
      RECT 1004.8200 2356.6800 2446.8800 2357.7600 ;
      RECT 9.3000 2356.6800 1002.6200 2357.7600 ;
      RECT 0.0000 2356.6800 5.7000 2357.7600 ;
      RECT 0.0000 2355.9300 3370.4200 2356.6800 ;
      RECT 1.1000 2355.0400 3370.4200 2355.9300 ;
      RECT 1.1000 2355.0300 1.7000 2355.0400 ;
      RECT 3368.7200 2353.9600 3370.4200 2355.0400 ;
      RECT 3305.0200 2353.9600 3365.1200 2355.0400 ;
      RECT 2497.4200 2353.9600 3302.8200 2355.0400 ;
      RECT 2446.4800 2353.9600 2495.2200 2355.0400 ;
      RECT 1007.4200 2353.9600 2444.2800 2355.0400 ;
      RECT 5.3000 2353.9600 1005.2200 2355.0400 ;
      RECT 0.0000 2353.9600 1.7000 2355.0300 ;
      RECT 0.0000 2352.3200 3370.4200 2353.9600 ;
      RECT 3364.7200 2351.2400 3370.4200 2352.3200 ;
      RECT 3307.6200 2351.2400 3361.1200 2352.3200 ;
      RECT 2494.8200 2351.2400 3305.4200 2352.3200 ;
      RECT 2449.0800 2351.2400 2492.6200 2352.3200 ;
      RECT 1004.8200 2351.2400 2446.8800 2352.3200 ;
      RECT 9.3000 2351.2400 1002.6200 2352.3200 ;
      RECT 0.0000 2351.2400 5.7000 2352.3200 ;
      RECT 0.0000 2349.6000 3370.4200 2351.2400 ;
      RECT 3368.7200 2348.5200 3370.4200 2349.6000 ;
      RECT 3305.0200 2348.5200 3365.1200 2349.6000 ;
      RECT 2497.4200 2348.5200 3302.8200 2349.6000 ;
      RECT 2446.4800 2348.5200 2495.2200 2349.6000 ;
      RECT 1007.4200 2348.5200 2444.2800 2349.6000 ;
      RECT 5.3000 2348.5200 1005.2200 2349.6000 ;
      RECT 0.0000 2348.5200 1.7000 2349.6000 ;
      RECT 0.0000 2346.8800 3370.4200 2348.5200 ;
      RECT 3364.7200 2345.8000 3370.4200 2346.8800 ;
      RECT 3307.6200 2345.8000 3361.1200 2346.8800 ;
      RECT 2494.8200 2345.8000 3305.4200 2346.8800 ;
      RECT 2449.0800 2345.8000 2492.6200 2346.8800 ;
      RECT 1004.8200 2345.8000 2446.8800 2346.8800 ;
      RECT 9.3000 2345.8000 1002.6200 2346.8800 ;
      RECT 0.0000 2345.8000 5.7000 2346.8800 ;
      RECT 0.0000 2344.9500 3370.4200 2345.8000 ;
      RECT 1.1000 2344.1600 3370.4200 2344.9500 ;
      RECT 1.1000 2344.0500 1.7000 2344.1600 ;
      RECT 3368.7200 2343.0800 3370.4200 2344.1600 ;
      RECT 3305.0200 2343.0800 3365.1200 2344.1600 ;
      RECT 2497.4200 2343.0800 3302.8200 2344.1600 ;
      RECT 2446.4800 2343.0800 2495.2200 2344.1600 ;
      RECT 1007.4200 2343.0800 2444.2800 2344.1600 ;
      RECT 5.3000 2343.0800 1005.2200 2344.1600 ;
      RECT 0.0000 2343.0800 1.7000 2344.0500 ;
      RECT 0.0000 2341.4400 3370.4200 2343.0800 ;
      RECT 3364.7200 2340.3600 3370.4200 2341.4400 ;
      RECT 3307.6200 2340.3600 3361.1200 2341.4400 ;
      RECT 2494.8200 2340.3600 3305.4200 2341.4400 ;
      RECT 2449.0800 2340.3600 2492.6200 2341.4400 ;
      RECT 1004.8200 2340.3600 2446.8800 2341.4400 ;
      RECT 9.3000 2340.3600 1002.6200 2341.4400 ;
      RECT 0.0000 2340.3600 5.7000 2341.4400 ;
      RECT 0.0000 2338.7200 3370.4200 2340.3600 ;
      RECT 3368.7200 2337.6400 3370.4200 2338.7200 ;
      RECT 3305.0200 2337.6400 3365.1200 2338.7200 ;
      RECT 2497.4200 2337.6400 3302.8200 2338.7200 ;
      RECT 2446.4800 2337.6400 2495.2200 2338.7200 ;
      RECT 1007.4200 2337.6400 2444.2800 2338.7200 ;
      RECT 5.3000 2337.6400 1005.2200 2338.7200 ;
      RECT 0.0000 2337.6400 1.7000 2338.7200 ;
      RECT 0.0000 2336.0000 3370.4200 2337.6400 ;
      RECT 3364.7200 2334.9200 3370.4200 2336.0000 ;
      RECT 3307.6200 2334.9200 3361.1200 2336.0000 ;
      RECT 2494.8200 2334.9200 3305.4200 2336.0000 ;
      RECT 2449.0800 2334.9200 2492.6200 2336.0000 ;
      RECT 1004.8200 2334.9200 2446.8800 2336.0000 ;
      RECT 9.3000 2334.9200 1002.6200 2336.0000 ;
      RECT 0.0000 2334.9200 5.7000 2336.0000 ;
      RECT 0.0000 2333.9700 3370.4200 2334.9200 ;
      RECT 1.1000 2333.2800 3370.4200 2333.9700 ;
      RECT 1.1000 2333.0700 1.7000 2333.2800 ;
      RECT 3368.7200 2332.2000 3370.4200 2333.2800 ;
      RECT 3305.0200 2332.2000 3365.1200 2333.2800 ;
      RECT 2497.4200 2332.2000 3302.8200 2333.2800 ;
      RECT 2446.4800 2332.2000 2495.2200 2333.2800 ;
      RECT 1007.4200 2332.2000 2444.2800 2333.2800 ;
      RECT 5.3000 2332.2000 1005.2200 2333.2800 ;
      RECT 0.0000 2332.2000 1.7000 2333.0700 ;
      RECT 0.0000 2330.5600 3370.4200 2332.2000 ;
      RECT 3364.7200 2329.4800 3370.4200 2330.5600 ;
      RECT 3307.6200 2329.4800 3361.1200 2330.5600 ;
      RECT 2494.8200 2329.4800 3305.4200 2330.5600 ;
      RECT 2449.0800 2329.4800 2492.6200 2330.5600 ;
      RECT 1004.8200 2329.4800 2446.8800 2330.5600 ;
      RECT 9.3000 2329.4800 1002.6200 2330.5600 ;
      RECT 0.0000 2329.4800 5.7000 2330.5600 ;
      RECT 0.0000 2327.8400 3370.4200 2329.4800 ;
      RECT 3368.7200 2326.7600 3370.4200 2327.8400 ;
      RECT 3305.0200 2326.7600 3365.1200 2327.8400 ;
      RECT 2497.4200 2326.7600 3302.8200 2327.8400 ;
      RECT 2446.4800 2326.7600 2495.2200 2327.8400 ;
      RECT 1007.4200 2326.7600 2444.2800 2327.8400 ;
      RECT 5.3000 2326.7600 1005.2200 2327.8400 ;
      RECT 0.0000 2326.7600 1.7000 2327.8400 ;
      RECT 0.0000 2325.1200 3370.4200 2326.7600 ;
      RECT 3364.7200 2324.0400 3370.4200 2325.1200 ;
      RECT 3307.6200 2324.0400 3361.1200 2325.1200 ;
      RECT 2494.8200 2324.0400 3305.4200 2325.1200 ;
      RECT 2449.0800 2324.0400 2492.6200 2325.1200 ;
      RECT 1004.8200 2324.0400 2446.8800 2325.1200 ;
      RECT 9.3000 2324.0400 1002.6200 2325.1200 ;
      RECT 0.0000 2324.0400 5.7000 2325.1200 ;
      RECT 0.0000 2322.9900 3370.4200 2324.0400 ;
      RECT 1.1000 2322.4000 3370.4200 2322.9900 ;
      RECT 1.1000 2322.0900 1.7000 2322.4000 ;
      RECT 3368.7200 2321.3200 3370.4200 2322.4000 ;
      RECT 3305.0200 2321.3200 3365.1200 2322.4000 ;
      RECT 2497.4200 2321.3200 3302.8200 2322.4000 ;
      RECT 2446.4800 2321.3200 2495.2200 2322.4000 ;
      RECT 1007.4200 2321.3200 2444.2800 2322.4000 ;
      RECT 5.3000 2321.3200 1005.2200 2322.4000 ;
      RECT 0.0000 2321.3200 1.7000 2322.0900 ;
      RECT 0.0000 2319.6800 3370.4200 2321.3200 ;
      RECT 3364.7200 2318.6000 3370.4200 2319.6800 ;
      RECT 3307.6200 2318.6000 3361.1200 2319.6800 ;
      RECT 2494.8200 2318.6000 3305.4200 2319.6800 ;
      RECT 2449.0800 2318.6000 2492.6200 2319.6800 ;
      RECT 1004.8200 2318.6000 2446.8800 2319.6800 ;
      RECT 9.3000 2318.6000 1002.6200 2319.6800 ;
      RECT 0.0000 2318.6000 5.7000 2319.6800 ;
      RECT 0.0000 2316.9600 3370.4200 2318.6000 ;
      RECT 3368.7200 2315.8800 3370.4200 2316.9600 ;
      RECT 3305.0200 2315.8800 3365.1200 2316.9600 ;
      RECT 2497.4200 2315.8800 3302.8200 2316.9600 ;
      RECT 2446.4800 2315.8800 2495.2200 2316.9600 ;
      RECT 1007.4200 2315.8800 2444.2800 2316.9600 ;
      RECT 5.3000 2315.8800 1005.2200 2316.9600 ;
      RECT 0.0000 2315.8800 1.7000 2316.9600 ;
      RECT 0.0000 2314.2400 3370.4200 2315.8800 ;
      RECT 3364.7200 2313.1600 3370.4200 2314.2400 ;
      RECT 3307.6200 2313.1600 3361.1200 2314.2400 ;
      RECT 2494.8200 2313.1600 3305.4200 2314.2400 ;
      RECT 2449.0800 2313.1600 2492.6200 2314.2400 ;
      RECT 1004.8200 2313.1600 2446.8800 2314.2400 ;
      RECT 9.3000 2313.1600 1002.6200 2314.2400 ;
      RECT 0.0000 2313.1600 5.7000 2314.2400 ;
      RECT 0.0000 2312.6200 3370.4200 2313.1600 ;
      RECT 1.1000 2311.7200 3370.4200 2312.6200 ;
      RECT 0.0000 2311.5200 3370.4200 2311.7200 ;
      RECT 3368.7200 2310.4400 3370.4200 2311.5200 ;
      RECT 3305.0200 2310.4400 3365.1200 2311.5200 ;
      RECT 2497.4200 2310.4400 3302.8200 2311.5200 ;
      RECT 2446.4800 2310.4400 2495.2200 2311.5200 ;
      RECT 1007.4200 2310.4400 2444.2800 2311.5200 ;
      RECT 5.3000 2310.4400 1005.2200 2311.5200 ;
      RECT 0.0000 2310.4400 1.7000 2311.5200 ;
      RECT 0.0000 2308.8000 3370.4200 2310.4400 ;
      RECT 3364.7200 2307.7200 3370.4200 2308.8000 ;
      RECT 3307.6200 2307.7200 3361.1200 2308.8000 ;
      RECT 2494.8200 2307.7200 3305.4200 2308.8000 ;
      RECT 2449.0800 2307.7200 2492.6200 2308.8000 ;
      RECT 1004.8200 2307.7200 2446.8800 2308.8000 ;
      RECT 9.3000 2307.7200 1002.6200 2308.8000 ;
      RECT 0.0000 2307.7200 5.7000 2308.8000 ;
      RECT 0.0000 2306.0800 3370.4200 2307.7200 ;
      RECT 3368.7200 2305.0000 3370.4200 2306.0800 ;
      RECT 3305.0200 2305.0000 3365.1200 2306.0800 ;
      RECT 2497.4200 2305.0000 3302.8200 2306.0800 ;
      RECT 2446.4800 2305.0000 2495.2200 2306.0800 ;
      RECT 1007.4200 2305.0000 2444.2800 2306.0800 ;
      RECT 5.3000 2305.0000 1005.2200 2306.0800 ;
      RECT 0.0000 2305.0000 1.7000 2306.0800 ;
      RECT 0.0000 2303.3600 3370.4200 2305.0000 ;
      RECT 3364.7200 2302.2800 3370.4200 2303.3600 ;
      RECT 3307.6200 2302.2800 3361.1200 2303.3600 ;
      RECT 2494.8200 2302.2800 3305.4200 2303.3600 ;
      RECT 2449.0800 2302.2800 2492.6200 2303.3600 ;
      RECT 1004.8200 2302.2800 2446.8800 2303.3600 ;
      RECT 9.3000 2302.2800 1002.6200 2303.3600 ;
      RECT 0.0000 2302.2800 5.7000 2303.3600 ;
      RECT 0.0000 2301.6400 3370.4200 2302.2800 ;
      RECT 1.1000 2300.7400 3370.4200 2301.6400 ;
      RECT 0.0000 2300.6400 3370.4200 2300.7400 ;
      RECT 3368.7200 2299.5600 3370.4200 2300.6400 ;
      RECT 3305.0200 2299.5600 3365.1200 2300.6400 ;
      RECT 2497.4200 2299.5600 3302.8200 2300.6400 ;
      RECT 2446.4800 2299.5600 2495.2200 2300.6400 ;
      RECT 1007.4200 2299.5600 2444.2800 2300.6400 ;
      RECT 5.3000 2299.5600 1005.2200 2300.6400 ;
      RECT 0.0000 2299.5600 1.7000 2300.6400 ;
      RECT 0.0000 2297.9200 3370.4200 2299.5600 ;
      RECT 3364.7200 2296.8400 3370.4200 2297.9200 ;
      RECT 3307.6200 2296.8400 3361.1200 2297.9200 ;
      RECT 2494.8200 2296.8400 3305.4200 2297.9200 ;
      RECT 2449.0800 2296.8400 2492.6200 2297.9200 ;
      RECT 1004.8200 2296.8400 2446.8800 2297.9200 ;
      RECT 9.3000 2296.8400 1002.6200 2297.9200 ;
      RECT 0.0000 2296.8400 5.7000 2297.9200 ;
      RECT 0.0000 2295.2000 3370.4200 2296.8400 ;
      RECT 3368.7200 2294.1200 3370.4200 2295.2000 ;
      RECT 3305.0200 2294.1200 3365.1200 2295.2000 ;
      RECT 2497.4200 2294.1200 3302.8200 2295.2000 ;
      RECT 2446.4800 2294.1200 2495.2200 2295.2000 ;
      RECT 1007.4200 2294.1200 2444.2800 2295.2000 ;
      RECT 5.3000 2294.1200 1005.2200 2295.2000 ;
      RECT 0.0000 2294.1200 1.7000 2295.2000 ;
      RECT 0.0000 2292.4800 3370.4200 2294.1200 ;
      RECT 3364.7200 2291.4000 3370.4200 2292.4800 ;
      RECT 3307.6200 2291.4000 3361.1200 2292.4800 ;
      RECT 2494.8200 2291.4000 3305.4200 2292.4800 ;
      RECT 2449.0800 2291.4000 2492.6200 2292.4800 ;
      RECT 1004.8200 2291.4000 2446.8800 2292.4800 ;
      RECT 9.3000 2291.4000 1002.6200 2292.4800 ;
      RECT 0.0000 2291.4000 5.7000 2292.4800 ;
      RECT 0.0000 2290.6600 3370.4200 2291.4000 ;
      RECT 1.1000 2289.7600 3370.4200 2290.6600 ;
      RECT 3368.7200 2288.6800 3370.4200 2289.7600 ;
      RECT 3305.0200 2288.6800 3365.1200 2289.7600 ;
      RECT 2497.4200 2288.6800 3302.8200 2289.7600 ;
      RECT 2446.4800 2288.6800 2495.2200 2289.7600 ;
      RECT 1007.4200 2288.6800 2444.2800 2289.7600 ;
      RECT 5.3000 2288.6800 1005.2200 2289.7600 ;
      RECT 0.0000 2288.6800 1.7000 2289.7600 ;
      RECT 0.0000 2287.0400 3370.4200 2288.6800 ;
      RECT 3364.7200 2285.9600 3370.4200 2287.0400 ;
      RECT 3307.6200 2285.9600 3361.1200 2287.0400 ;
      RECT 2494.8200 2285.9600 3305.4200 2287.0400 ;
      RECT 2449.0800 2285.9600 2492.6200 2287.0400 ;
      RECT 1004.8200 2285.9600 2446.8800 2287.0400 ;
      RECT 9.3000 2285.9600 1002.6200 2287.0400 ;
      RECT 0.0000 2285.9600 5.7000 2287.0400 ;
      RECT 0.0000 2284.3200 3370.4200 2285.9600 ;
      RECT 3368.7200 2283.2400 3370.4200 2284.3200 ;
      RECT 3305.0200 2283.2400 3365.1200 2284.3200 ;
      RECT 2497.4200 2283.2400 3302.8200 2284.3200 ;
      RECT 2446.4800 2283.2400 2495.2200 2284.3200 ;
      RECT 1007.4200 2283.2400 2444.2800 2284.3200 ;
      RECT 5.3000 2283.2400 1005.2200 2284.3200 ;
      RECT 0.0000 2283.2400 1.7000 2284.3200 ;
      RECT 0.0000 2281.6000 3370.4200 2283.2400 ;
      RECT 3364.7200 2280.5200 3370.4200 2281.6000 ;
      RECT 3307.6200 2280.5200 3361.1200 2281.6000 ;
      RECT 2494.8200 2280.5200 3305.4200 2281.6000 ;
      RECT 2449.0800 2280.5200 2492.6200 2281.6000 ;
      RECT 1004.8200 2280.5200 2446.8800 2281.6000 ;
      RECT 9.3000 2280.5200 1002.6200 2281.6000 ;
      RECT 0.0000 2280.5200 5.7000 2281.6000 ;
      RECT 0.0000 2279.6800 3370.4200 2280.5200 ;
      RECT 1.1000 2278.8800 3370.4200 2279.6800 ;
      RECT 1.1000 2278.7800 1.7000 2278.8800 ;
      RECT 3368.7200 2277.8000 3370.4200 2278.8800 ;
      RECT 3305.0200 2277.8000 3365.1200 2278.8800 ;
      RECT 2497.4200 2277.8000 3302.8200 2278.8800 ;
      RECT 2446.4800 2277.8000 2495.2200 2278.8800 ;
      RECT 1007.4200 2277.8000 2444.2800 2278.8800 ;
      RECT 5.3000 2277.8000 1005.2200 2278.8800 ;
      RECT 0.0000 2277.8000 1.7000 2278.7800 ;
      RECT 0.0000 2276.1600 3370.4200 2277.8000 ;
      RECT 3364.7200 2275.0800 3370.4200 2276.1600 ;
      RECT 3307.6200 2275.0800 3361.1200 2276.1600 ;
      RECT 2494.8200 2275.0800 3305.4200 2276.1600 ;
      RECT 2449.0800 2275.0800 2492.6200 2276.1600 ;
      RECT 1004.8200 2275.0800 2446.8800 2276.1600 ;
      RECT 9.3000 2275.0800 1002.6200 2276.1600 ;
      RECT 0.0000 2275.0800 5.7000 2276.1600 ;
      RECT 0.0000 2273.4400 3370.4200 2275.0800 ;
      RECT 3368.7200 2272.3600 3370.4200 2273.4400 ;
      RECT 3305.0200 2272.3600 3365.1200 2273.4400 ;
      RECT 2497.4200 2272.3600 3302.8200 2273.4400 ;
      RECT 2446.4800 2272.3600 2495.2200 2273.4400 ;
      RECT 1007.4200 2272.3600 2444.2800 2273.4400 ;
      RECT 5.3000 2272.3600 1005.2200 2273.4400 ;
      RECT 0.0000 2272.3600 1.7000 2273.4400 ;
      RECT 0.0000 2270.7200 3370.4200 2272.3600 ;
      RECT 3364.7200 2269.6400 3370.4200 2270.7200 ;
      RECT 3307.6200 2269.6400 3361.1200 2270.7200 ;
      RECT 2494.8200 2269.6400 3305.4200 2270.7200 ;
      RECT 2449.0800 2269.6400 2492.6200 2270.7200 ;
      RECT 1004.8200 2269.6400 2446.8800 2270.7200 ;
      RECT 9.3000 2269.6400 1002.6200 2270.7200 ;
      RECT 0.0000 2269.6400 5.7000 2270.7200 ;
      RECT 0.0000 2268.7000 3370.4200 2269.6400 ;
      RECT 1.1000 2268.0000 3370.4200 2268.7000 ;
      RECT 1.1000 2267.8000 1.7000 2268.0000 ;
      RECT 3368.7200 2266.9200 3370.4200 2268.0000 ;
      RECT 3305.0200 2266.9200 3365.1200 2268.0000 ;
      RECT 2497.4200 2266.9200 3302.8200 2268.0000 ;
      RECT 2446.4800 2266.9200 2495.2200 2268.0000 ;
      RECT 1007.4200 2266.9200 2444.2800 2268.0000 ;
      RECT 5.3000 2266.9200 1005.2200 2268.0000 ;
      RECT 0.0000 2266.9200 1.7000 2267.8000 ;
      RECT 0.0000 2265.2800 3370.4200 2266.9200 ;
      RECT 3364.7200 2264.2000 3370.4200 2265.2800 ;
      RECT 3307.6200 2264.2000 3361.1200 2265.2800 ;
      RECT 2494.8200 2264.2000 3305.4200 2265.2800 ;
      RECT 2449.0800 2264.2000 2492.6200 2265.2800 ;
      RECT 1004.8200 2264.2000 2446.8800 2265.2800 ;
      RECT 9.3000 2264.2000 1002.6200 2265.2800 ;
      RECT 0.0000 2264.2000 5.7000 2265.2800 ;
      RECT 0.0000 2263.3400 3370.4200 2264.2000 ;
      RECT 1057.5000 2263.0800 3370.4200 2263.3400 ;
      RECT 2396.3000 2262.5600 3370.4200 2263.0800 ;
      RECT 0.0000 2262.5600 1055.3000 2263.3400 ;
      RECT 1057.5000 2262.2600 2394.1000 2263.0800 ;
      RECT 1007.4200 2262.2600 1055.3000 2262.5600 ;
      RECT 2396.3000 2262.0000 2444.2800 2262.5600 ;
      RECT 1007.4200 2262.0000 2394.1000 2262.2600 ;
      RECT 3368.7200 2261.4800 3370.4200 2262.5600 ;
      RECT 3305.0200 2261.4800 3365.1200 2262.5600 ;
      RECT 2497.4200 2261.4800 3302.8200 2262.5600 ;
      RECT 2446.4800 2261.4800 2495.2200 2262.5600 ;
      RECT 1007.4200 2261.4800 2444.2800 2262.0000 ;
      RECT 5.3000 2261.4800 1005.2200 2262.5600 ;
      RECT 0.0000 2261.4800 1.7000 2262.5600 ;
      RECT 0.0000 2260.6200 3370.4200 2261.4800 ;
      RECT 1017.4800 2260.3600 3370.4200 2260.6200 ;
      RECT 2436.3200 2259.8400 3370.4200 2260.3600 ;
      RECT 0.0000 2259.8400 1015.2800 2260.6200 ;
      RECT 1017.4800 2259.5400 1295.6000 2260.3600 ;
      RECT 1004.8200 2259.5400 1015.2800 2259.8400 ;
      RECT 2436.3200 2259.2800 2446.8800 2259.8400 ;
      RECT 2178.6800 2259.2800 2434.1200 2260.3600 ;
      RECT 1738.2400 2259.2800 2176.4800 2260.3600 ;
      RECT 1518.0200 2259.2800 1736.0400 2260.3600 ;
      RECT 1297.8000 2259.2800 1515.8200 2260.3600 ;
      RECT 1004.8200 2259.2800 1295.6000 2259.5400 ;
      RECT 3364.7200 2258.7600 3370.4200 2259.8400 ;
      RECT 3307.6200 2258.7600 3361.1200 2259.8400 ;
      RECT 2494.8200 2258.7600 3305.4200 2259.8400 ;
      RECT 2449.0800 2258.7600 2492.6200 2259.8400 ;
      RECT 1004.8200 2258.7600 2446.8800 2259.2800 ;
      RECT 9.3000 2258.7600 1002.6200 2259.8400 ;
      RECT 0.0000 2258.7600 5.7000 2259.8400 ;
      RECT 0.0000 2258.3300 3370.4200 2258.7600 ;
      RECT 1.1000 2257.4500 3370.4200 2258.3300 ;
      RECT 1.1000 2257.4300 1005.2200 2257.4500 ;
      RECT 1065.1600 2257.2900 3370.4200 2257.4500 ;
      RECT 2446.4800 2257.1200 3370.4200 2257.2900 ;
      RECT 0.0000 2257.1200 1005.2200 2257.4300 ;
      RECT 3368.7200 2256.0400 3370.4200 2257.1200 ;
      RECT 3305.0200 2256.0400 3365.1200 2257.1200 ;
      RECT 2497.4200 2256.0400 3302.8200 2257.1200 ;
      RECT 2446.4800 2256.0400 2495.2200 2257.1200 ;
      RECT 5.3000 2256.0400 1005.2200 2257.1200 ;
      RECT 0.0000 2256.0400 1.7000 2257.1200 ;
      RECT 1065.1600 2255.2500 1283.0400 2257.2900 ;
      RECT 1011.2200 2255.2500 1059.1600 2257.4500 ;
      RECT 0.0000 2255.2500 1005.2200 2256.0400 ;
      RECT 2446.4800 2255.0900 3370.4200 2256.0400 ;
      RECT 2392.5400 2255.0900 2440.4800 2257.2900 ;
      RECT 2172.3200 2255.0900 2380.3400 2257.2900 ;
      RECT 1945.9000 2255.0900 2163.9200 2257.2900 ;
      RECT 1731.8800 2255.0900 1939.9000 2257.2900 ;
      RECT 1511.6600 2255.0900 1719.6800 2257.2900 ;
      RECT 1291.4400 2255.0900 1499.4600 2257.2900 ;
      RECT 0.0000 2255.0900 1283.0400 2255.2500 ;
      RECT 0.0000 2255.0500 3370.4200 2255.0900 ;
      RECT 1067.7600 2254.6900 3370.4200 2255.0500 ;
      RECT 2449.0800 2254.4000 3370.4200 2254.6900 ;
      RECT 0.0000 2254.4000 1002.6200 2255.0500 ;
      RECT 3364.7200 2253.3200 3370.4200 2254.4000 ;
      RECT 3307.6200 2253.3200 3361.1200 2254.4000 ;
      RECT 2494.8200 2253.3200 3305.4200 2254.4000 ;
      RECT 2449.0800 2253.3200 2492.6200 2254.4000 ;
      RECT 9.3000 2253.3200 1002.6200 2254.4000 ;
      RECT 0.0000 2253.3200 5.7000 2254.4000 ;
      RECT 1067.7600 2252.8500 1285.6400 2254.6900 ;
      RECT 1011.2200 2252.8500 1059.1600 2255.0500 ;
      RECT 0.0000 2252.8500 1002.6200 2253.3200 ;
      RECT 2449.0800 2252.4900 3370.4200 2253.3200 ;
      RECT 2392.5400 2252.4900 2440.4800 2254.6900 ;
      RECT 2172.3200 2252.4900 2386.7400 2254.6900 ;
      RECT 1948.5000 2252.4900 2166.5200 2254.6900 ;
      RECT 1731.8800 2252.4900 1939.9000 2254.6900 ;
      RECT 1511.6600 2252.4900 1719.6800 2254.6900 ;
      RECT 1291.4400 2252.4900 1499.4600 2254.6900 ;
      RECT 0.0000 2252.4900 1285.6400 2252.8500 ;
      RECT 0.0000 2251.6800 3370.4200 2252.4900 ;
      RECT 3368.7200 2250.6000 3370.4200 2251.6800 ;
      RECT 3305.0200 2250.6000 3365.1200 2251.6800 ;
      RECT 2497.4200 2250.6000 3302.8200 2251.6800 ;
      RECT 2446.4800 2250.6000 2495.2200 2251.6800 ;
      RECT 1007.4200 2250.6000 2444.2800 2251.6800 ;
      RECT 5.3000 2250.6000 1005.2200 2251.6800 ;
      RECT 0.0000 2250.6000 1.7000 2251.6800 ;
      RECT 0.0000 2248.9600 3370.4200 2250.6000 ;
      RECT 3364.7200 2247.8800 3370.4200 2248.9600 ;
      RECT 3307.6200 2247.8800 3361.1200 2248.9600 ;
      RECT 2494.8200 2247.8800 3305.4200 2248.9600 ;
      RECT 2449.0800 2247.8800 2492.6200 2248.9600 ;
      RECT 1004.8200 2247.8800 2446.8800 2248.9600 ;
      RECT 9.3000 2247.8800 1002.6200 2248.9600 ;
      RECT 0.0000 2247.8800 5.7000 2248.9600 ;
      RECT 0.0000 2247.5200 3370.4200 2247.8800 ;
      RECT 0.0000 2247.3500 1.7000 2247.5200 ;
      RECT 1065.1600 2247.2600 3370.4200 2247.5200 ;
      RECT 1.1000 2246.4500 1.7000 2247.3500 ;
      RECT 2446.4800 2246.2400 3370.4200 2247.2600 ;
      RECT 1065.1600 2245.3200 1283.0400 2247.2600 ;
      RECT 3368.7200 2245.1600 3370.4200 2246.2400 ;
      RECT 3305.0200 2245.1600 3365.1200 2246.2400 ;
      RECT 2497.4200 2245.1600 3302.8200 2246.2400 ;
      RECT 2446.4800 2245.1600 2495.2200 2246.2400 ;
      RECT 1007.4200 2245.1600 1283.0400 2245.3200 ;
      RECT 5.3000 2245.1600 1005.2200 2245.3200 ;
      RECT 0.0000 2245.1600 1.7000 2246.4500 ;
      RECT 2446.4800 2245.0600 3370.4200 2245.1600 ;
      RECT 1945.9000 2245.0600 2163.9200 2247.2600 ;
      RECT 0.0000 2245.0600 1283.0400 2245.1600 ;
      RECT 0.0000 2244.9200 3370.4200 2245.0600 ;
      RECT 1067.7600 2244.6600 3370.4200 2244.9200 ;
      RECT 2449.0800 2243.5200 3370.4200 2244.6600 ;
      RECT 1067.7600 2242.7200 1285.6400 2244.6600 ;
      RECT 1948.5000 2242.4600 2166.5200 2244.6600 ;
      RECT 1004.8200 2242.4600 1285.6400 2242.7200 ;
      RECT 3364.7200 2242.4400 3370.4200 2243.5200 ;
      RECT 3307.6200 2242.4400 3361.1200 2243.5200 ;
      RECT 2494.8200 2242.4400 3305.4200 2243.5200 ;
      RECT 2449.0800 2242.4400 2492.6200 2243.5200 ;
      RECT 1004.8200 2242.4400 2446.8800 2242.4600 ;
      RECT 9.3000 2242.4400 1002.6200 2242.7200 ;
      RECT 0.0000 2242.4400 5.7000 2244.9200 ;
      RECT 0.0000 2240.8000 3370.4200 2242.4400 ;
      RECT 3368.7200 2239.7200 3370.4200 2240.8000 ;
      RECT 3305.0200 2239.7200 3365.1200 2240.8000 ;
      RECT 2497.4200 2239.7200 3302.8200 2240.8000 ;
      RECT 2446.4800 2239.7200 2495.2200 2240.8000 ;
      RECT 1007.4200 2239.7200 2444.2800 2240.8000 ;
      RECT 5.3000 2239.7200 1005.2200 2240.8000 ;
      RECT 0.0000 2239.7200 1.7000 2240.8000 ;
      RECT 0.0000 2238.0800 3370.4200 2239.7200 ;
      RECT 3364.7200 2237.0000 3370.4200 2238.0800 ;
      RECT 3307.6200 2237.0000 3361.1200 2238.0800 ;
      RECT 2494.8200 2237.0000 3305.4200 2238.0800 ;
      RECT 2449.0800 2237.0000 2492.6200 2238.0800 ;
      RECT 1004.8200 2237.0000 2446.8800 2238.0800 ;
      RECT 9.3000 2237.0000 1002.6200 2238.0800 ;
      RECT 0.0000 2237.0000 5.7000 2238.0800 ;
      RECT 0.0000 2236.9100 3370.4200 2237.0000 ;
      RECT 1067.7600 2236.7500 3370.4200 2236.9100 ;
      RECT 0.0000 2236.3700 1002.6200 2236.9100 ;
      RECT 1.1000 2235.4700 1002.6200 2236.3700 ;
      RECT 2449.0800 2235.3600 3370.4200 2236.7500 ;
      RECT 0.0000 2235.3600 1002.6200 2235.4700 ;
      RECT 1067.7600 2234.7100 1285.6400 2236.7500 ;
      RECT 1011.2200 2234.7100 1059.1600 2236.9100 ;
      RECT 5.3000 2234.7100 1002.6200 2235.3600 ;
      RECT 2449.0800 2234.5500 2495.2200 2235.3600 ;
      RECT 2392.5400 2234.5500 2440.4800 2236.7500 ;
      RECT 2172.3200 2234.5500 2380.3400 2236.7500 ;
      RECT 1948.5000 2234.5500 2166.5200 2236.7500 ;
      RECT 1731.8800 2234.5500 1939.9000 2236.7500 ;
      RECT 1511.6600 2234.5500 1719.6800 2236.7500 ;
      RECT 1291.4400 2234.5500 1499.4600 2236.7500 ;
      RECT 1007.4200 2234.5500 1285.6400 2234.7100 ;
      RECT 1007.4200 2234.5100 2444.2800 2234.5500 ;
      RECT 3368.7200 2234.2800 3370.4200 2235.3600 ;
      RECT 3305.0200 2234.2800 3365.1200 2235.3600 ;
      RECT 2497.4200 2234.2800 3302.8200 2235.3600 ;
      RECT 2446.4800 2234.2800 2495.2200 2234.5500 ;
      RECT 5.3000 2234.2800 1005.2200 2234.7100 ;
      RECT 0.0000 2234.2800 1.7000 2235.3600 ;
      RECT 1065.1600 2234.1500 2444.2800 2234.5100 ;
      RECT 2446.4800 2232.6400 3370.4200 2234.2800 ;
      RECT 0.0000 2232.6400 1005.2200 2234.2800 ;
      RECT 1065.1600 2232.3100 1283.0400 2234.1500 ;
      RECT 1011.2200 2232.3100 1059.1600 2234.5100 ;
      RECT 1004.8200 2232.3100 1005.2200 2232.6400 ;
      RECT 2446.4800 2231.9500 2446.8800 2232.6400 ;
      RECT 2392.5400 2231.9500 2440.4800 2234.1500 ;
      RECT 2172.3200 2231.9500 2380.3400 2234.1500 ;
      RECT 1945.9000 2231.9500 2163.9200 2234.1500 ;
      RECT 1731.8800 2231.9500 1939.9000 2234.1500 ;
      RECT 1511.6600 2231.9500 1719.6800 2234.1500 ;
      RECT 1291.4400 2231.9500 1499.4600 2234.1500 ;
      RECT 1004.8200 2231.9500 1283.0400 2232.3100 ;
      RECT 3364.7200 2231.5600 3370.4200 2232.6400 ;
      RECT 3307.6200 2231.5600 3361.1200 2232.6400 ;
      RECT 2494.8200 2231.5600 3305.4200 2232.6400 ;
      RECT 2449.0800 2231.5600 2492.6200 2232.6400 ;
      RECT 1004.8200 2231.5600 2446.8800 2231.9500 ;
      RECT 9.3000 2231.5600 1002.6200 2232.6400 ;
      RECT 0.0000 2231.5600 5.7000 2232.6400 ;
      RECT 0.0000 2229.9200 3370.4200 2231.5600 ;
      RECT 1007.4200 2229.5400 2444.2800 2229.9200 ;
      RECT 1057.5000 2229.2800 2444.2800 2229.5400 ;
      RECT 3368.7200 2228.8400 3370.4200 2229.9200 ;
      RECT 3305.0200 2228.8400 3365.1200 2229.9200 ;
      RECT 2497.4200 2228.8400 3302.8200 2229.9200 ;
      RECT 2446.4800 2228.8400 2495.2200 2229.9200 ;
      RECT 2396.3000 2228.8400 2444.2800 2229.2800 ;
      RECT 1007.4200 2228.8400 1055.3000 2229.5400 ;
      RECT 5.3000 2228.8400 1005.2200 2229.9200 ;
      RECT 0.0000 2228.8400 1.7000 2229.9200 ;
      RECT 1057.5000 2228.4600 1293.0000 2229.2800 ;
      RECT 0.0000 2228.4600 1055.3000 2228.8400 ;
      RECT 2396.3000 2228.2000 3370.4200 2228.8400 ;
      RECT 2176.0800 2228.2000 2394.1000 2229.2800 ;
      RECT 1735.6400 2228.2000 2173.8800 2229.2800 ;
      RECT 1515.4200 2228.2000 1733.4400 2229.2800 ;
      RECT 1295.2000 2228.2000 1513.2200 2229.2800 ;
      RECT 0.0000 2228.2000 1293.0000 2228.4600 ;
      RECT 0.0000 2227.2000 3370.4200 2228.2000 ;
      RECT 3364.7200 2226.1200 3370.4200 2227.2000 ;
      RECT 3307.6200 2226.1200 3361.1200 2227.2000 ;
      RECT 2494.8200 2226.1200 3305.4200 2227.2000 ;
      RECT 2449.0800 2226.1200 2492.6200 2227.2000 ;
      RECT 1004.8200 2226.1200 2446.8800 2227.2000 ;
      RECT 9.3000 2226.1200 1002.6200 2227.2000 ;
      RECT 0.0000 2226.1200 5.7000 2227.2000 ;
      RECT 0.0000 2225.3900 3370.4200 2226.1200 ;
      RECT 1.1000 2224.4900 3370.4200 2225.3900 ;
      RECT 0.0000 2224.4800 3370.4200 2224.4900 ;
      RECT 3368.7200 2223.4000 3370.4200 2224.4800 ;
      RECT 3305.0200 2223.4000 3365.1200 2224.4800 ;
      RECT 2497.4200 2223.4000 3302.8200 2224.4800 ;
      RECT 2446.4800 2223.4000 2495.2200 2224.4800 ;
      RECT 1007.4200 2223.4000 2444.2800 2224.4800 ;
      RECT 5.3000 2223.4000 1005.2200 2224.4800 ;
      RECT 0.0000 2223.4000 1.7000 2224.4800 ;
      RECT 0.0000 2221.7600 3370.4200 2223.4000 ;
      RECT 3364.7200 2220.6800 3370.4200 2221.7600 ;
      RECT 3307.6200 2220.6800 3361.1200 2221.7600 ;
      RECT 2494.8200 2220.6800 3305.4200 2221.7600 ;
      RECT 2449.0800 2220.6800 2492.6200 2221.7600 ;
      RECT 1004.8200 2220.6800 2446.8800 2221.7600 ;
      RECT 9.3000 2220.6800 1002.6200 2221.7600 ;
      RECT 0.0000 2220.6800 5.7000 2221.7600 ;
      RECT 0.0000 2219.0400 3370.4200 2220.6800 ;
      RECT 3368.7200 2217.9600 3370.4200 2219.0400 ;
      RECT 3305.0200 2217.9600 3365.1200 2219.0400 ;
      RECT 2497.4200 2217.9600 3302.8200 2219.0400 ;
      RECT 2446.4800 2217.9600 2495.2200 2219.0400 ;
      RECT 1007.4200 2217.9600 2444.2800 2219.0400 ;
      RECT 5.3000 2217.9600 1005.2200 2219.0400 ;
      RECT 0.0000 2217.9600 1.7000 2219.0400 ;
      RECT 0.0000 2216.3200 3370.4200 2217.9600 ;
      RECT 3364.7200 2215.2400 3370.4200 2216.3200 ;
      RECT 3307.6200 2215.2400 3361.1200 2216.3200 ;
      RECT 2494.8200 2215.2400 3305.4200 2216.3200 ;
      RECT 2449.0800 2215.2400 2492.6200 2216.3200 ;
      RECT 1004.8200 2215.2400 2446.8800 2216.3200 ;
      RECT 9.3000 2215.2400 1002.6200 2216.3200 ;
      RECT 0.0000 2215.2400 5.7000 2216.3200 ;
      RECT 0.0000 2214.4100 3370.4200 2215.2400 ;
      RECT 1.1000 2213.6000 3370.4200 2214.4100 ;
      RECT 1.1000 2213.5100 1.7000 2213.6000 ;
      RECT 3368.7200 2212.5200 3370.4200 2213.6000 ;
      RECT 3305.0200 2212.5200 3365.1200 2213.6000 ;
      RECT 2497.4200 2212.5200 3302.8200 2213.6000 ;
      RECT 2446.4800 2212.5200 2495.2200 2213.6000 ;
      RECT 1007.4200 2212.5200 2444.2800 2213.6000 ;
      RECT 5.3000 2212.5200 1005.2200 2213.6000 ;
      RECT 0.0000 2212.5200 1.7000 2213.5100 ;
      RECT 0.0000 2210.8800 3370.4200 2212.5200 ;
      RECT 3364.7200 2209.8000 3370.4200 2210.8800 ;
      RECT 3307.6200 2209.8000 3361.1200 2210.8800 ;
      RECT 2494.8200 2209.8000 3305.4200 2210.8800 ;
      RECT 2449.0800 2209.8000 2492.6200 2210.8800 ;
      RECT 1004.8200 2209.8000 2446.8800 2210.8800 ;
      RECT 9.3000 2209.8000 1002.6200 2210.8800 ;
      RECT 0.0000 2209.8000 5.7000 2210.8800 ;
      RECT 0.0000 2208.1600 3370.4200 2209.8000 ;
      RECT 3368.7200 2207.0800 3370.4200 2208.1600 ;
      RECT 3305.0200 2207.0800 3365.1200 2208.1600 ;
      RECT 2497.4200 2207.0800 3302.8200 2208.1600 ;
      RECT 2446.4800 2207.0800 2495.2200 2208.1600 ;
      RECT 1007.4200 2207.0800 2444.2800 2208.1600 ;
      RECT 5.3000 2207.0800 1005.2200 2208.1600 ;
      RECT 0.0000 2207.0800 1.7000 2208.1600 ;
      RECT 0.0000 2205.4400 3370.4200 2207.0800 ;
      RECT 3364.7200 2204.3600 3370.4200 2205.4400 ;
      RECT 3307.6200 2204.3600 3361.1200 2205.4400 ;
      RECT 2494.8200 2204.3600 3305.4200 2205.4400 ;
      RECT 2449.0800 2204.3600 2492.6200 2205.4400 ;
      RECT 1004.8200 2204.3600 2446.8800 2205.4400 ;
      RECT 9.3000 2204.3600 1002.6200 2205.4400 ;
      RECT 0.0000 2204.3600 5.7000 2205.4400 ;
      RECT 0.0000 2204.0400 3370.4200 2204.3600 ;
      RECT 1.1000 2203.1400 3370.4200 2204.0400 ;
      RECT 0.0000 2202.7200 3370.4200 2203.1400 ;
      RECT 3368.7200 2201.6400 3370.4200 2202.7200 ;
      RECT 3305.0200 2201.6400 3365.1200 2202.7200 ;
      RECT 2497.4200 2201.6400 3302.8200 2202.7200 ;
      RECT 2446.4800 2201.6400 2495.2200 2202.7200 ;
      RECT 1007.4200 2201.6400 2444.2800 2202.7200 ;
      RECT 5.3000 2201.6400 1005.2200 2202.7200 ;
      RECT 0.0000 2201.6400 1.7000 2202.7200 ;
      RECT 0.0000 2200.0000 3370.4200 2201.6400 ;
      RECT 3364.7200 2198.9200 3370.4200 2200.0000 ;
      RECT 3307.6200 2198.9200 3361.1200 2200.0000 ;
      RECT 2494.8200 2198.9200 3305.4200 2200.0000 ;
      RECT 2449.0800 2198.9200 2492.6200 2200.0000 ;
      RECT 1004.8200 2198.9200 2446.8800 2200.0000 ;
      RECT 9.3000 2198.9200 1002.6200 2200.0000 ;
      RECT 0.0000 2198.9200 5.7000 2200.0000 ;
      RECT 0.0000 2197.2800 3370.4200 2198.9200 ;
      RECT 3368.7200 2196.2000 3370.4200 2197.2800 ;
      RECT 3305.0200 2196.2000 3365.1200 2197.2800 ;
      RECT 2497.4200 2196.2000 3302.8200 2197.2800 ;
      RECT 2446.4800 2196.2000 2495.2200 2197.2800 ;
      RECT 1007.4200 2196.2000 2444.2800 2197.2800 ;
      RECT 5.3000 2196.2000 1005.2200 2197.2800 ;
      RECT 0.0000 2196.2000 1.7000 2197.2800 ;
      RECT 0.0000 2194.5600 3370.4200 2196.2000 ;
      RECT 3364.7200 2193.4800 3370.4200 2194.5600 ;
      RECT 3307.6200 2193.4800 3361.1200 2194.5600 ;
      RECT 2494.8200 2193.4800 3305.4200 2194.5600 ;
      RECT 2449.0800 2193.4800 2492.6200 2194.5600 ;
      RECT 1004.8200 2193.4800 2446.8800 2194.5600 ;
      RECT 9.3000 2193.4800 1002.6200 2194.5600 ;
      RECT 0.0000 2193.4800 5.7000 2194.5600 ;
      RECT 0.0000 2193.0600 3370.4200 2193.4800 ;
      RECT 1.1000 2192.1600 3370.4200 2193.0600 ;
      RECT 0.0000 2191.8400 3370.4200 2192.1600 ;
      RECT 3368.7200 2190.7600 3370.4200 2191.8400 ;
      RECT 3305.0200 2190.7600 3365.1200 2191.8400 ;
      RECT 2497.4200 2190.7600 3302.8200 2191.8400 ;
      RECT 2446.4800 2190.7600 2495.2200 2191.8400 ;
      RECT 1007.4200 2190.7600 2444.2800 2191.8400 ;
      RECT 5.3000 2190.7600 1005.2200 2191.8400 ;
      RECT 0.0000 2190.7600 1.7000 2191.8400 ;
      RECT 0.0000 2189.1200 3370.4200 2190.7600 ;
      RECT 3364.7200 2188.0400 3370.4200 2189.1200 ;
      RECT 3307.6200 2188.0400 3361.1200 2189.1200 ;
      RECT 2494.8200 2188.0400 3305.4200 2189.1200 ;
      RECT 2449.0800 2188.0400 2492.6200 2189.1200 ;
      RECT 1004.8200 2188.0400 2446.8800 2189.1200 ;
      RECT 9.3000 2188.0400 1002.6200 2189.1200 ;
      RECT 0.0000 2188.0400 5.7000 2189.1200 ;
      RECT 0.0000 2186.4000 3370.4200 2188.0400 ;
      RECT 3368.7200 2185.3200 3370.4200 2186.4000 ;
      RECT 3305.0200 2185.3200 3365.1200 2186.4000 ;
      RECT 2497.4200 2185.3200 3302.8200 2186.4000 ;
      RECT 2446.4800 2185.3200 2495.2200 2186.4000 ;
      RECT 1007.4200 2185.3200 2444.2800 2186.4000 ;
      RECT 5.3000 2185.3200 1005.2200 2186.4000 ;
      RECT 0.0000 2185.3200 1.7000 2186.4000 ;
      RECT 0.0000 2183.6800 3370.4200 2185.3200 ;
      RECT 3364.7200 2182.6000 3370.4200 2183.6800 ;
      RECT 3307.6200 2182.6000 3361.1200 2183.6800 ;
      RECT 2494.8200 2182.6000 3305.4200 2183.6800 ;
      RECT 2449.0800 2182.6000 2492.6200 2183.6800 ;
      RECT 1004.8200 2182.6000 2446.8800 2183.6800 ;
      RECT 9.3000 2182.6000 1002.6200 2183.6800 ;
      RECT 0.0000 2182.6000 5.7000 2183.6800 ;
      RECT 0.0000 2182.0800 3370.4200 2182.6000 ;
      RECT 1.1000 2181.1800 3370.4200 2182.0800 ;
      RECT 0.0000 2180.9600 3370.4200 2181.1800 ;
      RECT 3368.7200 2179.8800 3370.4200 2180.9600 ;
      RECT 3305.0200 2179.8800 3365.1200 2180.9600 ;
      RECT 2497.4200 2179.8800 3302.8200 2180.9600 ;
      RECT 2446.4800 2179.8800 2495.2200 2180.9600 ;
      RECT 1007.4200 2179.8800 2444.2800 2180.9600 ;
      RECT 5.3000 2179.8800 1005.2200 2180.9600 ;
      RECT 0.0000 2179.8800 1.7000 2180.9600 ;
      RECT 0.0000 2178.2400 3370.4200 2179.8800 ;
      RECT 3364.7200 2177.1600 3370.4200 2178.2400 ;
      RECT 3307.6200 2177.1600 3361.1200 2178.2400 ;
      RECT 2494.8200 2177.1600 3305.4200 2178.2400 ;
      RECT 2449.0800 2177.1600 2492.6200 2178.2400 ;
      RECT 1004.8200 2177.1600 2446.8800 2178.2400 ;
      RECT 9.3000 2177.1600 1002.6200 2178.2400 ;
      RECT 0.0000 2177.1600 5.7000 2178.2400 ;
      RECT 0.0000 2175.5200 3370.4200 2177.1600 ;
      RECT 3368.7200 2174.4400 3370.4200 2175.5200 ;
      RECT 3305.0200 2174.4400 3365.1200 2175.5200 ;
      RECT 2497.4200 2174.4400 3302.8200 2175.5200 ;
      RECT 2446.4800 2174.4400 2495.2200 2175.5200 ;
      RECT 1007.4200 2174.4400 2444.2800 2175.5200 ;
      RECT 5.3000 2174.4400 1005.2200 2175.5200 ;
      RECT 0.0000 2174.4400 1.7000 2175.5200 ;
      RECT 0.0000 2172.8000 3370.4200 2174.4400 ;
      RECT 3364.7200 2171.7200 3370.4200 2172.8000 ;
      RECT 3307.6200 2171.7200 3361.1200 2172.8000 ;
      RECT 2494.8200 2171.7200 3305.4200 2172.8000 ;
      RECT 2449.0800 2171.7200 2492.6200 2172.8000 ;
      RECT 1004.8200 2171.7200 2446.8800 2172.8000 ;
      RECT 9.3000 2171.7200 1002.6200 2172.8000 ;
      RECT 0.0000 2171.7200 5.7000 2172.8000 ;
      RECT 0.0000 2171.1000 3370.4200 2171.7200 ;
      RECT 1.1000 2170.2000 3370.4200 2171.1000 ;
      RECT 0.0000 2170.0800 3370.4200 2170.2000 ;
      RECT 3368.7200 2169.0000 3370.4200 2170.0800 ;
      RECT 3305.0200 2169.0000 3365.1200 2170.0800 ;
      RECT 2497.4200 2169.0000 3302.8200 2170.0800 ;
      RECT 2446.4800 2169.0000 2495.2200 2170.0800 ;
      RECT 1007.4200 2169.0000 2444.2800 2170.0800 ;
      RECT 5.3000 2169.0000 1005.2200 2170.0800 ;
      RECT 0.0000 2169.0000 1.7000 2170.0800 ;
      RECT 0.0000 2167.3600 3370.4200 2169.0000 ;
      RECT 3364.7200 2166.2800 3370.4200 2167.3600 ;
      RECT 3307.6200 2166.2800 3361.1200 2167.3600 ;
      RECT 2494.8200 2166.2800 3305.4200 2167.3600 ;
      RECT 2449.0800 2166.2800 2492.6200 2167.3600 ;
      RECT 1004.8200 2166.2800 2446.8800 2167.3600 ;
      RECT 9.3000 2166.2800 1002.6200 2167.3600 ;
      RECT 0.0000 2166.2800 5.7000 2167.3600 ;
      RECT 0.0000 2164.6400 3370.4200 2166.2800 ;
      RECT 3368.7200 2163.5600 3370.4200 2164.6400 ;
      RECT 3305.0200 2163.5600 3365.1200 2164.6400 ;
      RECT 2497.4200 2163.5600 3302.8200 2164.6400 ;
      RECT 2446.4800 2163.5600 2495.2200 2164.6400 ;
      RECT 1007.4200 2163.5600 2444.2800 2164.6400 ;
      RECT 5.3000 2163.5600 1005.2200 2164.6400 ;
      RECT 0.0000 2163.5600 1.7000 2164.6400 ;
      RECT 0.0000 2161.9200 3370.4200 2163.5600 ;
      RECT 3364.7200 2160.8400 3370.4200 2161.9200 ;
      RECT 3307.6200 2160.8400 3361.1200 2161.9200 ;
      RECT 2494.8200 2160.8400 3305.4200 2161.9200 ;
      RECT 2449.0800 2160.8400 2492.6200 2161.9200 ;
      RECT 1004.8200 2160.8400 2446.8800 2161.9200 ;
      RECT 9.3000 2160.8400 1002.6200 2161.9200 ;
      RECT 0.0000 2160.8400 5.7000 2161.9200 ;
      RECT 0.0000 2160.1200 3370.4200 2160.8400 ;
      RECT 1.1000 2159.2200 3370.4200 2160.1200 ;
      RECT 0.0000 2159.2000 3370.4200 2159.2200 ;
      RECT 3368.7200 2158.1200 3370.4200 2159.2000 ;
      RECT 3305.0200 2158.1200 3365.1200 2159.2000 ;
      RECT 2497.4200 2158.1200 3302.8200 2159.2000 ;
      RECT 2446.4800 2158.1200 2495.2200 2159.2000 ;
      RECT 1007.4200 2158.1200 2444.2800 2159.2000 ;
      RECT 5.3000 2158.1200 1005.2200 2159.2000 ;
      RECT 0.0000 2158.1200 1.7000 2159.2000 ;
      RECT 0.0000 2156.4800 3370.4200 2158.1200 ;
      RECT 3364.7200 2155.4000 3370.4200 2156.4800 ;
      RECT 3307.6200 2155.4000 3361.1200 2156.4800 ;
      RECT 2494.8200 2155.4000 3305.4200 2156.4800 ;
      RECT 2449.0800 2155.4000 2492.6200 2156.4800 ;
      RECT 1004.8200 2155.4000 2446.8800 2156.4800 ;
      RECT 9.3000 2155.4000 1002.6200 2156.4800 ;
      RECT 0.0000 2155.4000 5.7000 2156.4800 ;
      RECT 0.0000 2153.7600 3370.4200 2155.4000 ;
      RECT 3368.7200 2152.6800 3370.4200 2153.7600 ;
      RECT 3305.0200 2152.6800 3365.1200 2153.7600 ;
      RECT 2497.4200 2152.6800 3302.8200 2153.7600 ;
      RECT 2446.4800 2152.6800 2495.2200 2153.7600 ;
      RECT 1007.4200 2152.6800 2444.2800 2153.7600 ;
      RECT 5.3000 2152.6800 1005.2200 2153.7600 ;
      RECT 0.0000 2152.6800 1.7000 2153.7600 ;
      RECT 0.0000 2151.0400 3370.4200 2152.6800 ;
      RECT 3364.7200 2149.9600 3370.4200 2151.0400 ;
      RECT 3307.6200 2149.9600 3361.1200 2151.0400 ;
      RECT 2494.8200 2149.9600 3305.4200 2151.0400 ;
      RECT 2449.0800 2149.9600 2492.6200 2151.0400 ;
      RECT 1004.8200 2149.9600 2446.8800 2151.0400 ;
      RECT 9.3000 2149.9600 1002.6200 2151.0400 ;
      RECT 0.0000 2149.9600 5.7000 2151.0400 ;
      RECT 0.0000 2149.7500 3370.4200 2149.9600 ;
      RECT 1.1000 2148.8500 3370.4200 2149.7500 ;
      RECT 0.0000 2148.3200 3370.4200 2148.8500 ;
      RECT 3368.7200 2147.2400 3370.4200 2148.3200 ;
      RECT 3305.0200 2147.2400 3365.1200 2148.3200 ;
      RECT 2497.4200 2147.2400 3302.8200 2148.3200 ;
      RECT 2446.4800 2147.2400 2495.2200 2148.3200 ;
      RECT 1007.4200 2147.2400 2444.2800 2148.3200 ;
      RECT 5.3000 2147.2400 1005.2200 2148.3200 ;
      RECT 0.0000 2147.2400 1.7000 2148.3200 ;
      RECT 0.0000 2145.6000 3370.4200 2147.2400 ;
      RECT 3364.7200 2144.5200 3370.4200 2145.6000 ;
      RECT 3307.6200 2144.5200 3361.1200 2145.6000 ;
      RECT 2494.8200 2144.5200 3305.4200 2145.6000 ;
      RECT 2449.0800 2144.5200 2492.6200 2145.6000 ;
      RECT 1004.8200 2144.5200 2446.8800 2145.6000 ;
      RECT 9.3000 2144.5200 1002.6200 2145.6000 ;
      RECT 0.0000 2144.5200 5.7000 2145.6000 ;
      RECT 0.0000 2142.8800 3370.4200 2144.5200 ;
      RECT 3368.7200 2141.8000 3370.4200 2142.8800 ;
      RECT 3305.0200 2141.8000 3365.1200 2142.8800 ;
      RECT 2497.4200 2141.8000 3302.8200 2142.8800 ;
      RECT 2446.4800 2141.8000 2495.2200 2142.8800 ;
      RECT 1007.4200 2141.8000 2444.2800 2142.8800 ;
      RECT 5.3000 2141.8000 1005.2200 2142.8800 ;
      RECT 0.0000 2141.8000 1.7000 2142.8800 ;
      RECT 0.0000 2140.1600 3370.4200 2141.8000 ;
      RECT 3364.7200 2139.0800 3370.4200 2140.1600 ;
      RECT 3307.6200 2139.0800 3361.1200 2140.1600 ;
      RECT 2494.8200 2139.0800 3305.4200 2140.1600 ;
      RECT 2449.0800 2139.0800 2492.6200 2140.1600 ;
      RECT 1004.8200 2139.0800 2446.8800 2140.1600 ;
      RECT 9.3000 2139.0800 1002.6200 2140.1600 ;
      RECT 0.0000 2139.0800 5.7000 2140.1600 ;
      RECT 0.0000 2138.7700 3370.4200 2139.0800 ;
      RECT 1.1000 2137.8700 3370.4200 2138.7700 ;
      RECT 0.0000 2137.4400 3370.4200 2137.8700 ;
      RECT 3368.7200 2136.3600 3370.4200 2137.4400 ;
      RECT 3305.0200 2136.3600 3365.1200 2137.4400 ;
      RECT 2497.4200 2136.3600 3302.8200 2137.4400 ;
      RECT 2446.4800 2136.3600 2495.2200 2137.4400 ;
      RECT 1007.4200 2136.3600 2444.2800 2137.4400 ;
      RECT 5.3000 2136.3600 1005.2200 2137.4400 ;
      RECT 0.0000 2136.3600 1.7000 2137.4400 ;
      RECT 0.0000 2134.7200 3370.4200 2136.3600 ;
      RECT 3364.7200 2133.6400 3370.4200 2134.7200 ;
      RECT 3307.6200 2133.6400 3361.1200 2134.7200 ;
      RECT 2494.8200 2133.6400 3305.4200 2134.7200 ;
      RECT 2449.0800 2133.6400 2492.6200 2134.7200 ;
      RECT 1004.8200 2133.6400 2446.8800 2134.7200 ;
      RECT 9.3000 2133.6400 1002.6200 2134.7200 ;
      RECT 0.0000 2133.6400 5.7000 2134.7200 ;
      RECT 0.0000 2132.0000 3370.4200 2133.6400 ;
      RECT 3368.7200 2130.9200 3370.4200 2132.0000 ;
      RECT 3305.0200 2130.9200 3365.1200 2132.0000 ;
      RECT 2497.4200 2130.9200 3302.8200 2132.0000 ;
      RECT 2446.4800 2130.9200 2495.2200 2132.0000 ;
      RECT 1007.4200 2130.9200 2444.2800 2132.0000 ;
      RECT 5.3000 2130.9200 1005.2200 2132.0000 ;
      RECT 0.0000 2130.9200 1.7000 2132.0000 ;
      RECT 0.0000 2129.2800 3370.4200 2130.9200 ;
      RECT 3364.7200 2128.2000 3370.4200 2129.2800 ;
      RECT 3307.6200 2128.2000 3361.1200 2129.2800 ;
      RECT 2494.8200 2128.2000 3305.4200 2129.2800 ;
      RECT 2449.0800 2128.2000 2492.6200 2129.2800 ;
      RECT 1004.8200 2128.2000 2446.8800 2129.2800 ;
      RECT 9.3000 2128.2000 1002.6200 2129.2800 ;
      RECT 0.0000 2128.2000 5.7000 2129.2800 ;
      RECT 0.0000 2127.7900 3370.4200 2128.2000 ;
      RECT 1.1000 2126.8900 3370.4200 2127.7900 ;
      RECT 0.0000 2126.5600 3370.4200 2126.8900 ;
      RECT 3368.7200 2125.4800 3370.4200 2126.5600 ;
      RECT 3305.0200 2125.4800 3365.1200 2126.5600 ;
      RECT 2497.4200 2125.4800 3302.8200 2126.5600 ;
      RECT 2446.4800 2125.4800 2495.2200 2126.5600 ;
      RECT 1007.4200 2125.4800 2444.2800 2126.5600 ;
      RECT 5.3000 2125.4800 1005.2200 2126.5600 ;
      RECT 0.0000 2125.4800 1.7000 2126.5600 ;
      RECT 0.0000 2123.8400 3370.4200 2125.4800 ;
      RECT 3364.7200 2122.7600 3370.4200 2123.8400 ;
      RECT 3307.6200 2122.7600 3361.1200 2123.8400 ;
      RECT 2494.8200 2122.7600 3305.4200 2123.8400 ;
      RECT 2449.0800 2122.7600 2492.6200 2123.8400 ;
      RECT 1004.8200 2122.7600 2446.8800 2123.8400 ;
      RECT 9.3000 2122.7600 1002.6200 2123.8400 ;
      RECT 0.0000 2122.7600 5.7000 2123.8400 ;
      RECT 0.0000 2121.1200 3370.4200 2122.7600 ;
      RECT 3368.7200 2120.0400 3370.4200 2121.1200 ;
      RECT 3305.0200 2120.0400 3365.1200 2121.1200 ;
      RECT 2497.4200 2120.0400 3302.8200 2121.1200 ;
      RECT 2446.4800 2120.0400 2495.2200 2121.1200 ;
      RECT 1007.4200 2120.0400 2444.2800 2121.1200 ;
      RECT 5.3000 2120.0400 1005.2200 2121.1200 ;
      RECT 0.0000 2120.0400 1.7000 2121.1200 ;
      RECT 0.0000 2118.4000 3370.4200 2120.0400 ;
      RECT 3364.7200 2117.3200 3370.4200 2118.4000 ;
      RECT 3307.6200 2117.3200 3361.1200 2118.4000 ;
      RECT 2494.8200 2117.3200 3305.4200 2118.4000 ;
      RECT 2449.0800 2117.3200 2492.6200 2118.4000 ;
      RECT 1004.8200 2117.3200 2446.8800 2118.4000 ;
      RECT 9.3000 2117.3200 1002.6200 2118.4000 ;
      RECT 0.0000 2117.3200 5.7000 2118.4000 ;
      RECT 0.0000 2116.8100 3370.4200 2117.3200 ;
      RECT 1.1000 2115.9100 3370.4200 2116.8100 ;
      RECT 0.0000 2115.6800 3370.4200 2115.9100 ;
      RECT 3368.7200 2114.6000 3370.4200 2115.6800 ;
      RECT 3305.0200 2114.6000 3365.1200 2115.6800 ;
      RECT 2497.4200 2114.6000 3302.8200 2115.6800 ;
      RECT 2446.4800 2114.6000 2495.2200 2115.6800 ;
      RECT 1007.4200 2114.6000 2444.2800 2115.6800 ;
      RECT 5.3000 2114.6000 1005.2200 2115.6800 ;
      RECT 0.0000 2114.6000 1.7000 2115.6800 ;
      RECT 0.0000 2112.9600 3370.4200 2114.6000 ;
      RECT 3364.7200 2111.8800 3370.4200 2112.9600 ;
      RECT 3307.6200 2111.8800 3361.1200 2112.9600 ;
      RECT 2494.8200 2111.8800 3305.4200 2112.9600 ;
      RECT 2449.0800 2111.8800 2492.6200 2112.9600 ;
      RECT 1004.8200 2111.8800 2446.8800 2112.9600 ;
      RECT 9.3000 2111.8800 1002.6200 2112.9600 ;
      RECT 0.0000 2111.8800 5.7000 2112.9600 ;
      RECT 0.0000 2110.2400 3370.4200 2111.8800 ;
      RECT 3368.7200 2109.1600 3370.4200 2110.2400 ;
      RECT 3305.0200 2109.1600 3365.1200 2110.2400 ;
      RECT 2497.4200 2109.1600 3302.8200 2110.2400 ;
      RECT 2446.4800 2109.1600 2495.2200 2110.2400 ;
      RECT 1007.4200 2109.1600 2444.2800 2110.2400 ;
      RECT 5.3000 2109.1600 1005.2200 2110.2400 ;
      RECT 0.0000 2109.1600 1.7000 2110.2400 ;
      RECT 0.0000 2107.5200 3370.4200 2109.1600 ;
      RECT 3364.7200 2106.4400 3370.4200 2107.5200 ;
      RECT 3307.6200 2106.4400 3361.1200 2107.5200 ;
      RECT 2494.8200 2106.4400 3305.4200 2107.5200 ;
      RECT 2449.0800 2106.4400 2492.6200 2107.5200 ;
      RECT 1004.8200 2106.4400 2446.8800 2107.5200 ;
      RECT 9.3000 2106.4400 1002.6200 2107.5200 ;
      RECT 0.0000 2106.4400 5.7000 2107.5200 ;
      RECT 0.0000 2105.8300 3370.4200 2106.4400 ;
      RECT 1.1000 2104.9300 3370.4200 2105.8300 ;
      RECT 0.0000 2104.8000 3370.4200 2104.9300 ;
      RECT 3368.7200 2103.7200 3370.4200 2104.8000 ;
      RECT 3305.0200 2103.7200 3365.1200 2104.8000 ;
      RECT 2497.4200 2103.7200 3302.8200 2104.8000 ;
      RECT 2446.4800 2103.7200 2495.2200 2104.8000 ;
      RECT 1007.4200 2103.7200 2444.2800 2104.8000 ;
      RECT 5.3000 2103.7200 1005.2200 2104.8000 ;
      RECT 0.0000 2103.7200 1.7000 2104.8000 ;
      RECT 0.0000 2102.0800 3370.4200 2103.7200 ;
      RECT 3364.7200 2101.0000 3370.4200 2102.0800 ;
      RECT 3307.6200 2101.0000 3361.1200 2102.0800 ;
      RECT 2494.8200 2101.0000 3305.4200 2102.0800 ;
      RECT 2449.0800 2101.0000 2492.6200 2102.0800 ;
      RECT 1004.8200 2101.0000 2446.8800 2102.0800 ;
      RECT 9.3000 2101.0000 1002.6200 2102.0800 ;
      RECT 0.0000 2101.0000 5.7000 2102.0800 ;
      RECT 0.0000 2099.3600 3370.4200 2101.0000 ;
      RECT 3368.7200 2098.2800 3370.4200 2099.3600 ;
      RECT 3305.0200 2098.2800 3365.1200 2099.3600 ;
      RECT 2497.4200 2098.2800 3302.8200 2099.3600 ;
      RECT 2446.4800 2098.2800 2495.2200 2099.3600 ;
      RECT 1007.4200 2098.2800 2444.2800 2099.3600 ;
      RECT 5.3000 2098.2800 1005.2200 2099.3600 ;
      RECT 0.0000 2098.2800 1.7000 2099.3600 ;
      RECT 0.0000 2096.6400 3370.4200 2098.2800 ;
      RECT 3364.7200 2095.5600 3370.4200 2096.6400 ;
      RECT 3307.6200 2095.5600 3361.1200 2096.6400 ;
      RECT 2494.8200 2095.5600 3305.4200 2096.6400 ;
      RECT 2449.0800 2095.5600 2492.6200 2096.6400 ;
      RECT 1004.8200 2095.5600 2446.8800 2096.6400 ;
      RECT 9.3000 2095.5600 1002.6200 2096.6400 ;
      RECT 0.0000 2095.5600 5.7000 2096.6400 ;
      RECT 0.0000 2095.4600 3370.4200 2095.5600 ;
      RECT 1.1000 2094.5600 3370.4200 2095.4600 ;
      RECT 0.0000 2093.9200 3370.4200 2094.5600 ;
      RECT 3368.7200 2092.8400 3370.4200 2093.9200 ;
      RECT 3305.0200 2092.8400 3365.1200 2093.9200 ;
      RECT 2497.4200 2092.8400 3302.8200 2093.9200 ;
      RECT 2446.4800 2092.8400 2495.2200 2093.9200 ;
      RECT 1007.4200 2092.8400 2444.2800 2093.9200 ;
      RECT 5.3000 2092.8400 1005.2200 2093.9200 ;
      RECT 0.0000 2092.8400 1.7000 2093.9200 ;
      RECT 0.0000 2091.2000 3370.4200 2092.8400 ;
      RECT 3364.7200 2090.1200 3370.4200 2091.2000 ;
      RECT 3307.6200 2090.1200 3361.1200 2091.2000 ;
      RECT 2494.8200 2090.1200 3305.4200 2091.2000 ;
      RECT 2449.0800 2090.1200 2492.6200 2091.2000 ;
      RECT 1004.8200 2090.1200 2446.8800 2091.2000 ;
      RECT 9.3000 2090.1200 1002.6200 2091.2000 ;
      RECT 0.0000 2090.1200 5.7000 2091.2000 ;
      RECT 0.0000 2088.4800 3370.4200 2090.1200 ;
      RECT 3368.7200 2087.4000 3370.4200 2088.4800 ;
      RECT 3305.0200 2087.4000 3365.1200 2088.4800 ;
      RECT 2497.4200 2087.4000 3302.8200 2088.4800 ;
      RECT 2446.4800 2087.4000 2495.2200 2088.4800 ;
      RECT 1007.4200 2087.4000 2444.2800 2088.4800 ;
      RECT 5.3000 2087.4000 1005.2200 2088.4800 ;
      RECT 0.0000 2087.4000 1.7000 2088.4800 ;
      RECT 0.0000 2085.7600 3370.4200 2087.4000 ;
      RECT 3364.7200 2084.6800 3370.4200 2085.7600 ;
      RECT 3307.6200 2084.6800 3361.1200 2085.7600 ;
      RECT 2494.8200 2084.6800 3305.4200 2085.7600 ;
      RECT 2449.0800 2084.6800 2492.6200 2085.7600 ;
      RECT 1004.8200 2084.6800 2446.8800 2085.7600 ;
      RECT 9.3000 2084.6800 1002.6200 2085.7600 ;
      RECT 0.0000 2084.6800 5.7000 2085.7600 ;
      RECT 0.0000 2084.4800 3370.4200 2084.6800 ;
      RECT 1.1000 2083.5800 3370.4200 2084.4800 ;
      RECT 0.0000 2083.0400 3370.4200 2083.5800 ;
      RECT 3368.7200 2081.9600 3370.4200 2083.0400 ;
      RECT 3305.0200 2081.9600 3365.1200 2083.0400 ;
      RECT 2497.4200 2081.9600 3302.8200 2083.0400 ;
      RECT 2446.4800 2081.9600 2495.2200 2083.0400 ;
      RECT 1007.4200 2081.9600 2444.2800 2083.0400 ;
      RECT 5.3000 2081.9600 1005.2200 2083.0400 ;
      RECT 0.0000 2081.9600 1.7000 2083.0400 ;
      RECT 0.0000 2080.3200 3370.4200 2081.9600 ;
      RECT 3364.7200 2079.2400 3370.4200 2080.3200 ;
      RECT 3307.6200 2079.2400 3361.1200 2080.3200 ;
      RECT 2494.8200 2079.2400 3305.4200 2080.3200 ;
      RECT 2449.0800 2079.2400 2492.6200 2080.3200 ;
      RECT 1004.8200 2079.2400 2446.8800 2080.3200 ;
      RECT 9.3000 2079.2400 1002.6200 2080.3200 ;
      RECT 0.0000 2079.2400 5.7000 2080.3200 ;
      RECT 0.0000 2077.6000 3370.4200 2079.2400 ;
      RECT 3368.7200 2076.5200 3370.4200 2077.6000 ;
      RECT 3305.0200 2076.5200 3365.1200 2077.6000 ;
      RECT 2497.4200 2076.5200 3302.8200 2077.6000 ;
      RECT 2446.4800 2076.5200 2495.2200 2077.6000 ;
      RECT 1007.4200 2076.5200 2444.2800 2077.6000 ;
      RECT 5.3000 2076.5200 1005.2200 2077.6000 ;
      RECT 0.0000 2076.5200 1.7000 2077.6000 ;
      RECT 0.0000 2074.8800 3370.4200 2076.5200 ;
      RECT 3364.7200 2073.8000 3370.4200 2074.8800 ;
      RECT 3307.6200 2073.8000 3361.1200 2074.8800 ;
      RECT 2494.8200 2073.8000 3305.4200 2074.8800 ;
      RECT 2449.0800 2073.8000 2492.6200 2074.8800 ;
      RECT 1004.8200 2073.8000 2446.8800 2074.8800 ;
      RECT 9.3000 2073.8000 1002.6200 2074.8800 ;
      RECT 0.0000 2073.8000 5.7000 2074.8800 ;
      RECT 0.0000 2073.5000 3370.4200 2073.8000 ;
      RECT 1.1000 2072.6000 3370.4200 2073.5000 ;
      RECT 0.0000 2072.1600 3370.4200 2072.6000 ;
      RECT 3368.7200 2071.0800 3370.4200 2072.1600 ;
      RECT 3305.0200 2071.0800 3365.1200 2072.1600 ;
      RECT 2497.4200 2071.0800 3302.8200 2072.1600 ;
      RECT 2446.4800 2071.0800 2495.2200 2072.1600 ;
      RECT 1007.4200 2071.0800 2444.2800 2072.1600 ;
      RECT 5.3000 2071.0800 1005.2200 2072.1600 ;
      RECT 0.0000 2071.0800 1.7000 2072.1600 ;
      RECT 0.0000 2069.4400 3370.4200 2071.0800 ;
      RECT 3364.7200 2068.3600 3370.4200 2069.4400 ;
      RECT 3307.6200 2068.3600 3361.1200 2069.4400 ;
      RECT 2494.8200 2068.3600 3305.4200 2069.4400 ;
      RECT 2449.0800 2068.3600 2492.6200 2069.4400 ;
      RECT 1004.8200 2068.3600 2446.8800 2069.4400 ;
      RECT 9.3000 2068.3600 1002.6200 2069.4400 ;
      RECT 0.0000 2068.3600 5.7000 2069.4400 ;
      RECT 0.0000 2066.7200 3370.4200 2068.3600 ;
      RECT 3368.7200 2065.6400 3370.4200 2066.7200 ;
      RECT 3305.0200 2065.6400 3365.1200 2066.7200 ;
      RECT 2497.4200 2065.6400 3302.8200 2066.7200 ;
      RECT 2446.4800 2065.6400 2495.2200 2066.7200 ;
      RECT 1007.4200 2065.6400 2444.2800 2066.7200 ;
      RECT 5.3000 2065.6400 1005.2200 2066.7200 ;
      RECT 0.0000 2065.6400 1.7000 2066.7200 ;
      RECT 0.0000 2064.0000 3370.4200 2065.6400 ;
      RECT 3364.7200 2062.9200 3370.4200 2064.0000 ;
      RECT 3307.6200 2062.9200 3361.1200 2064.0000 ;
      RECT 2494.8200 2062.9200 3305.4200 2064.0000 ;
      RECT 2449.0800 2062.9200 2492.6200 2064.0000 ;
      RECT 1004.8200 2062.9200 2446.8800 2064.0000 ;
      RECT 9.3000 2062.9200 1002.6200 2064.0000 ;
      RECT 0.0000 2062.9200 5.7000 2064.0000 ;
      RECT 0.0000 2062.5200 3370.4200 2062.9200 ;
      RECT 1.1000 2061.6200 3370.4200 2062.5200 ;
      RECT 0.0000 2061.2800 3370.4200 2061.6200 ;
      RECT 3368.7200 2060.2000 3370.4200 2061.2800 ;
      RECT 3305.0200 2060.2000 3365.1200 2061.2800 ;
      RECT 2497.4200 2060.2000 3302.8200 2061.2800 ;
      RECT 2446.4800 2060.2000 2495.2200 2061.2800 ;
      RECT 1007.4200 2060.2000 2444.2800 2061.2800 ;
      RECT 5.3000 2060.2000 1005.2200 2061.2800 ;
      RECT 0.0000 2060.2000 1.7000 2061.2800 ;
      RECT 0.0000 2058.5600 3370.4200 2060.2000 ;
      RECT 3364.7200 2057.4800 3370.4200 2058.5600 ;
      RECT 3307.6200 2057.4800 3361.1200 2058.5600 ;
      RECT 2494.8200 2057.4800 3305.4200 2058.5600 ;
      RECT 2449.0800 2057.4800 2492.6200 2058.5600 ;
      RECT 1004.8200 2057.4800 2446.8800 2058.5600 ;
      RECT 9.3000 2057.4800 1002.6200 2058.5600 ;
      RECT 0.0000 2057.4800 5.7000 2058.5600 ;
      RECT 0.0000 2055.8400 3370.4200 2057.4800 ;
      RECT 3368.7200 2054.7600 3370.4200 2055.8400 ;
      RECT 3305.0200 2054.7600 3365.1200 2055.8400 ;
      RECT 2497.4200 2054.7600 3302.8200 2055.8400 ;
      RECT 2446.4800 2054.7600 2495.2200 2055.8400 ;
      RECT 1007.4200 2054.7600 2444.2800 2055.8400 ;
      RECT 5.3000 2054.7600 1005.2200 2055.8400 ;
      RECT 0.0000 2054.7600 1.7000 2055.8400 ;
      RECT 0.0000 2053.1200 3370.4200 2054.7600 ;
      RECT 3364.7200 2052.0400 3370.4200 2053.1200 ;
      RECT 3307.6200 2052.0400 3361.1200 2053.1200 ;
      RECT 2494.8200 2052.0400 3305.4200 2053.1200 ;
      RECT 2449.0800 2052.0400 2492.6200 2053.1200 ;
      RECT 1004.8200 2052.0400 2446.8800 2053.1200 ;
      RECT 9.3000 2052.0400 1002.6200 2053.1200 ;
      RECT 0.0000 2052.0400 5.7000 2053.1200 ;
      RECT 0.0000 2051.5400 3370.4200 2052.0400 ;
      RECT 1.1000 2050.6400 3370.4200 2051.5400 ;
      RECT 0.0000 2050.4000 3370.4200 2050.6400 ;
      RECT 3368.7200 2049.3200 3370.4200 2050.4000 ;
      RECT 3305.0200 2049.3200 3365.1200 2050.4000 ;
      RECT 2497.4200 2049.3200 3302.8200 2050.4000 ;
      RECT 2446.4800 2049.3200 2495.2200 2050.4000 ;
      RECT 1007.4200 2049.3200 2444.2800 2050.4000 ;
      RECT 5.3000 2049.3200 1005.2200 2050.4000 ;
      RECT 0.0000 2049.3200 1.7000 2050.4000 ;
      RECT 0.0000 2047.6800 3370.4200 2049.3200 ;
      RECT 3364.7200 2046.6000 3370.4200 2047.6800 ;
      RECT 3307.6200 2046.6000 3361.1200 2047.6800 ;
      RECT 2494.8200 2046.6000 3305.4200 2047.6800 ;
      RECT 2449.0800 2046.6000 2492.6200 2047.6800 ;
      RECT 1004.8200 2046.6000 2446.8800 2047.6800 ;
      RECT 9.3000 2046.6000 1002.6200 2047.6800 ;
      RECT 0.0000 2046.6000 5.7000 2047.6800 ;
      RECT 0.0000 2044.9600 3370.4200 2046.6000 ;
      RECT 3368.7200 2043.8800 3370.4200 2044.9600 ;
      RECT 3305.0200 2043.8800 3365.1200 2044.9600 ;
      RECT 2497.4200 2043.8800 3302.8200 2044.9600 ;
      RECT 2446.4800 2043.8800 2495.2200 2044.9600 ;
      RECT 1007.4200 2043.8800 2444.2800 2044.9600 ;
      RECT 5.3000 2043.8800 1005.2200 2044.9600 ;
      RECT 0.0000 2043.8800 1.7000 2044.9600 ;
      RECT 0.0000 2042.2400 3370.4200 2043.8800 ;
      RECT 0.0000 2041.1700 5.7000 2042.2400 ;
      RECT 3364.7200 2041.1600 3370.4200 2042.2400 ;
      RECT 3307.6200 2041.1600 3361.1200 2042.2400 ;
      RECT 2494.8200 2041.1600 3305.4200 2042.2400 ;
      RECT 2449.0800 2041.1600 2492.6200 2042.2400 ;
      RECT 1004.8200 2041.1600 2446.8800 2042.2400 ;
      RECT 9.3000 2041.1600 1002.6200 2042.2400 ;
      RECT 1.1000 2041.1600 5.7000 2041.1700 ;
      RECT 1.1000 2040.2700 3370.4200 2041.1600 ;
      RECT 0.0000 2039.5200 3370.4200 2040.2700 ;
      RECT 3368.7200 2038.4400 3370.4200 2039.5200 ;
      RECT 3305.0200 2038.4400 3365.1200 2039.5200 ;
      RECT 2497.4200 2038.4400 3302.8200 2039.5200 ;
      RECT 2446.4800 2038.4400 2495.2200 2039.5200 ;
      RECT 1007.4200 2038.4400 2444.2800 2039.5200 ;
      RECT 5.3000 2038.4400 1005.2200 2039.5200 ;
      RECT 0.0000 2038.4400 1.7000 2039.5200 ;
      RECT 0.0000 2036.8000 3370.4200 2038.4400 ;
      RECT 3364.7200 2035.7200 3370.4200 2036.8000 ;
      RECT 3307.6200 2035.7200 3361.1200 2036.8000 ;
      RECT 2494.8200 2035.7200 3305.4200 2036.8000 ;
      RECT 2449.0800 2035.7200 2492.6200 2036.8000 ;
      RECT 1004.8200 2035.7200 2446.8800 2036.8000 ;
      RECT 9.3000 2035.7200 1002.6200 2036.8000 ;
      RECT 0.0000 2035.7200 5.7000 2036.8000 ;
      RECT 0.0000 2034.0800 3370.4200 2035.7200 ;
      RECT 3368.7200 2033.0000 3370.4200 2034.0800 ;
      RECT 3305.0200 2033.0000 3365.1200 2034.0800 ;
      RECT 2497.4200 2033.0000 3302.8200 2034.0800 ;
      RECT 2446.4800 2033.0000 2495.2200 2034.0800 ;
      RECT 1007.4200 2033.0000 2444.2800 2034.0800 ;
      RECT 5.3000 2033.0000 1005.2200 2034.0800 ;
      RECT 0.0000 2033.0000 1.7000 2034.0800 ;
      RECT 0.0000 2031.3600 3370.4200 2033.0000 ;
      RECT 1004.8200 2030.9800 2446.8800 2031.3600 ;
      RECT 1077.7200 2030.7200 2446.8800 2030.9800 ;
      RECT 3364.7200 2030.2800 3370.4200 2031.3600 ;
      RECT 3307.6200 2030.2800 3361.1200 2031.3600 ;
      RECT 2494.8200 2030.2800 3305.4200 2031.3600 ;
      RECT 2449.0800 2030.2800 2492.6200 2031.3600 ;
      RECT 2436.3200 2030.2800 2446.8800 2030.7200 ;
      RECT 1004.8200 2030.2800 1015.2800 2030.9800 ;
      RECT 9.3000 2030.2800 1002.6200 2031.3600 ;
      RECT 0.0000 2030.2800 5.7000 2031.3600 ;
      RECT 0.0000 2030.1900 1015.2800 2030.2800 ;
      RECT 1077.7200 2029.9000 1295.6000 2030.7200 ;
      RECT 1017.4800 2029.9000 1075.5200 2030.9800 ;
      RECT 1.1000 2029.9000 1015.2800 2030.1900 ;
      RECT 2436.3200 2029.6400 3370.4200 2030.2800 ;
      RECT 2178.6800 2029.6400 2434.1200 2030.7200 ;
      RECT 1958.4600 2029.6400 2176.4800 2030.7200 ;
      RECT 1738.2400 2029.6400 1956.2600 2030.7200 ;
      RECT 1518.0200 2029.6400 1736.0400 2030.7200 ;
      RECT 1297.8000 2029.6400 1515.8200 2030.7200 ;
      RECT 1.1000 2029.6400 1295.6000 2029.9000 ;
      RECT 1.1000 2029.2900 3370.4200 2029.6400 ;
      RECT 0.0000 2028.6400 3370.4200 2029.2900 ;
      RECT 1007.4200 2027.9100 2444.2800 2028.6400 ;
      RECT 1007.4200 2027.8100 1062.9600 2027.9100 ;
      RECT 1285.3800 2027.6500 2444.2800 2027.9100 ;
      RECT 3368.7200 2027.5600 3370.4200 2028.6400 ;
      RECT 3305.0200 2027.5600 3365.1200 2028.6400 ;
      RECT 2497.4200 2027.5600 3302.8200 2028.6400 ;
      RECT 2446.4800 2027.5600 2495.2200 2028.6400 ;
      RECT 5.3000 2027.5600 1005.2200 2028.6400 ;
      RECT 0.0000 2027.5600 1.7000 2028.6400 ;
      RECT 2446.4800 2025.9200 3370.4200 2027.5600 ;
      RECT 0.0000 2025.9200 1005.2200 2027.5600 ;
      RECT 1071.3600 2025.7100 1279.3800 2027.9100 ;
      RECT 1065.1600 2025.6100 1283.0400 2025.7100 ;
      RECT 1011.2200 2025.6100 1059.1600 2027.8100 ;
      RECT 1002.1300 2025.6100 1005.2200 2025.9200 ;
      RECT 2446.4800 2025.4500 2446.8800 2025.9200 ;
      RECT 2392.5400 2025.4500 2440.4800 2027.6500 ;
      RECT 2172.3200 2025.4500 2380.3400 2027.6500 ;
      RECT 1952.1000 2025.4500 2160.1200 2027.6500 ;
      RECT 1731.8800 2025.4500 1939.9000 2027.6500 ;
      RECT 1511.6600 2025.4500 1719.6800 2027.6500 ;
      RECT 1291.4400 2025.4500 1499.4600 2027.6500 ;
      RECT 1002.1300 2025.4500 1283.0400 2025.6100 ;
      RECT 1002.1300 2025.4100 2446.8800 2025.4500 ;
      RECT 1011.2200 2025.3100 2446.8800 2025.4100 ;
      RECT 1287.9800 2025.0500 2446.8800 2025.3100 ;
      RECT 3364.7200 2024.8400 3370.4200 2025.9200 ;
      RECT 3307.6200 2024.8400 3361.1200 2025.9200 ;
      RECT 2494.8200 2024.8400 3305.4200 2025.9200 ;
      RECT 2449.0800 2024.8400 2492.6200 2025.9200 ;
      RECT 1002.1300 2024.8400 1002.6200 2025.4100 ;
      RECT 9.3000 2024.8400 1001.0300 2025.9200 ;
      RECT 0.0000 2024.8400 5.7000 2025.9200 ;
      RECT 1011.2200 2023.2100 1065.5600 2025.3100 ;
      RECT 0.0000 2023.2100 1002.6200 2024.8400 ;
      RECT 2449.0800 2023.2000 3370.4200 2024.8400 ;
      RECT 0.0000 2023.2000 1065.5600 2023.2100 ;
      RECT 1071.3600 2023.1100 1279.3800 2025.3100 ;
      RECT 1007.4200 2023.1100 1065.5600 2023.2000 ;
      RECT 2449.0800 2022.8500 2495.2200 2023.2000 ;
      RECT 2392.5400 2022.8500 2440.4800 2025.0500 ;
      RECT 2172.3200 2022.8500 2380.3400 2025.0500 ;
      RECT 1952.1000 2022.8500 2166.5200 2025.0500 ;
      RECT 1731.8800 2022.8500 1939.9000 2025.0500 ;
      RECT 1511.6600 2022.8500 1719.6800 2025.0500 ;
      RECT 1291.4400 2022.8500 1499.4600 2025.0500 ;
      RECT 1007.4200 2022.8500 1285.6400 2023.1100 ;
      RECT 3368.7200 2022.1200 3370.4200 2023.2000 ;
      RECT 3305.0200 2022.1200 3365.1200 2023.2000 ;
      RECT 2497.4200 2022.1200 3302.8200 2023.2000 ;
      RECT 2446.4800 2022.1200 2495.2200 2022.8500 ;
      RECT 1007.4200 2022.1200 2444.2800 2022.8500 ;
      RECT 5.3000 2022.1200 1005.2200 2023.2000 ;
      RECT 0.0000 2022.1200 1.7000 2023.2000 ;
      RECT 2446.4800 2021.9500 3370.4200 2022.1200 ;
      RECT 0.0000 2021.9500 2444.2800 2022.1200 ;
      RECT 0.0000 2020.4800 3370.4200 2021.9500 ;
      RECT 3364.7200 2019.4000 3370.4200 2020.4800 ;
      RECT 3307.6200 2019.4000 3361.1200 2020.4800 ;
      RECT 2494.8200 2019.4000 3305.4200 2020.4800 ;
      RECT 2449.0800 2019.4000 2492.6200 2020.4800 ;
      RECT 1004.8200 2019.4000 2446.8800 2020.4800 ;
      RECT 9.3000 2019.4000 1002.6200 2020.4800 ;
      RECT 0.0000 2019.4000 5.7000 2020.4800 ;
      RECT 0.0000 2019.2100 3370.4200 2019.4000 ;
      RECT 1.1000 2018.3100 3370.4200 2019.2100 ;
      RECT 0.0000 2017.8800 3370.4200 2018.3100 ;
      RECT 1285.3800 2017.7600 3370.4200 2017.8800 ;
      RECT 1285.3800 2017.6200 2444.2800 2017.7600 ;
      RECT 3368.7200 2016.6800 3370.4200 2017.7600 ;
      RECT 3305.0200 2016.6800 3365.1200 2017.7600 ;
      RECT 2497.4200 2016.6800 3302.8200 2017.7600 ;
      RECT 2446.4800 2016.6800 2495.2200 2017.7600 ;
      RECT 0.0000 2015.6800 1.7000 2017.8800 ;
      RECT 2446.4800 2015.4200 3370.4200 2016.6800 ;
      RECT 0.0000 2015.4200 1283.0400 2015.6800 ;
      RECT 0.0000 2015.3800 3370.4200 2015.4200 ;
      RECT 1065.0600 2015.2800 3370.4200 2015.3800 ;
      RECT 0.0000 2015.2800 1062.6600 2015.3800 ;
      RECT 1287.9800 2015.1200 3370.4200 2015.2800 ;
      RECT 1945.8000 2015.0400 3370.4200 2015.1200 ;
      RECT 1945.8000 2015.0200 2446.8800 2015.0400 ;
      RECT 1287.9800 2015.0200 1943.4000 2015.1200 ;
      RECT 3364.7200 2013.9600 3370.4200 2015.0400 ;
      RECT 3307.6200 2013.9600 3361.1200 2015.0400 ;
      RECT 2494.8200 2013.9600 3305.4200 2015.0400 ;
      RECT 2449.0800 2013.9600 2492.6200 2015.0400 ;
      RECT 0.0000 2013.0800 5.7000 2015.2800 ;
      RECT 2449.0800 2012.8200 3370.4200 2013.9600 ;
      RECT 1065.0600 2012.8200 1285.6400 2013.0800 ;
      RECT 1945.8000 2012.3200 3370.4200 2012.8200 ;
      RECT 0.0000 2012.3200 1062.6600 2013.0800 ;
      RECT 1065.0600 2011.3800 1943.4000 2012.8200 ;
      RECT 1007.4200 2011.3800 1062.6600 2012.3200 ;
      RECT 3368.7200 2011.2400 3370.4200 2012.3200 ;
      RECT 3305.0200 2011.2400 3365.1200 2012.3200 ;
      RECT 2497.4200 2011.2400 3302.8200 2012.3200 ;
      RECT 2446.4800 2011.2400 2495.2200 2012.3200 ;
      RECT 1945.8000 2011.2400 2444.2800 2012.3200 ;
      RECT 1007.4200 2011.2400 1943.4000 2011.3800 ;
      RECT 965.0200 2011.2400 1005.2200 2012.3200 ;
      RECT 157.4200 2011.2400 962.8200 2012.3200 ;
      RECT 5.3000 2011.2400 155.2200 2012.3200 ;
      RECT 0.0000 2011.2400 1.7000 2012.3200 ;
      RECT 1945.8000 2011.1200 3370.4200 2011.2400 ;
      RECT 0.0000 2011.1200 1943.4000 2011.2400 ;
      RECT 0.0000 2009.6000 3370.4200 2011.1200 ;
      RECT 3364.7200 2008.5200 3370.4200 2009.6000 ;
      RECT 3307.6200 2008.5200 3361.1200 2009.6000 ;
      RECT 2494.8200 2008.5200 3305.4200 2009.6000 ;
      RECT 2449.0800 2008.5200 2492.6200 2009.6000 ;
      RECT 1004.8200 2008.5200 2446.8800 2009.6000 ;
      RECT 967.6200 2008.5200 1002.6200 2009.6000 ;
      RECT 154.8200 2008.5200 965.4200 2009.6000 ;
      RECT 9.3000 2008.5200 152.6200 2009.6000 ;
      RECT 0.0000 2008.5200 5.7000 2009.6000 ;
      RECT 0.0000 2008.4200 3370.4200 2008.5200 ;
      RECT 0.0000 2008.2300 1065.5600 2008.4200 ;
      RECT 1287.9800 2008.1600 3370.4200 2008.4200 ;
      RECT 2168.7200 2008.0700 3370.4200 2008.1600 ;
      RECT 1.1000 2008.0700 1065.5600 2008.2300 ;
      RECT 1.1000 2007.3300 1005.2200 2008.0700 ;
      RECT 1007.4200 2007.2700 1065.5600 2008.0700 ;
      RECT 0.0000 2007.2700 1005.2200 2007.3300 ;
      RECT 2446.4800 2007.1100 3370.4200 2008.0700 ;
      RECT 2168.7200 2007.1100 2444.2800 2008.0700 ;
      RECT 1287.9800 2007.1100 1946.3000 2008.1600 ;
      RECT 2449.0800 2006.8800 3370.4200 2007.1100 ;
      RECT 0.0000 2006.8800 1002.6200 2007.2700 ;
      RECT 1071.3600 2006.2200 1279.3800 2008.4200 ;
      RECT 1062.4600 2006.2200 1065.5600 2007.2700 ;
      RECT 1952.1000 2005.9600 2160.1200 2008.1600 ;
      RECT 1943.2000 2005.9600 1946.3000 2007.1100 ;
      RECT 1062.4600 2005.8200 1285.6400 2006.2200 ;
      RECT 3368.7200 2005.8000 3370.4200 2006.8800 ;
      RECT 3305.0200 2005.8000 3365.1200 2006.8800 ;
      RECT 2497.4200 2005.8000 3302.8200 2006.8800 ;
      RECT 2449.0800 2005.8000 2495.2200 2006.8800 ;
      RECT 965.0200 2005.8000 1002.6200 2006.8800 ;
      RECT 157.4200 2005.8000 962.8200 2006.8800 ;
      RECT 5.3000 2005.8000 155.2200 2006.8800 ;
      RECT 0.0000 2005.8000 1.7000 2006.8800 ;
      RECT 1943.2000 2005.5600 2166.5200 2005.9600 ;
      RECT 1062.4600 2005.0700 1062.9600 2005.8200 ;
      RECT 1011.2200 2005.0700 1059.1600 2007.2700 ;
      RECT 0.0000 2005.0700 1002.6200 2005.8000 ;
      RECT 2449.0800 2004.9100 3370.4200 2005.8000 ;
      RECT 2392.5400 2004.9100 2440.4800 2007.1100 ;
      RECT 2172.3200 2004.9100 2380.3400 2007.1100 ;
      RECT 2166.1200 2004.9100 2166.5200 2005.5600 ;
      RECT 1943.2000 2004.9100 1943.7000 2005.5600 ;
      RECT 1731.8800 2004.9100 1939.9000 2007.1100 ;
      RECT 1511.6600 2004.9100 1719.6800 2007.1100 ;
      RECT 1291.4400 2004.9100 1499.4600 2007.1100 ;
      RECT 1285.3800 2004.9100 1285.6400 2005.8200 ;
      RECT 0.0000 2004.8700 1062.9600 2005.0700 ;
      RECT 2166.1200 2004.5100 3370.4200 2004.9100 ;
      RECT 1285.3800 2004.5100 1943.7000 2004.9100 ;
      RECT 2446.4800 2004.1600 3370.4200 2004.5100 ;
      RECT 0.0000 2004.1600 1005.2200 2004.8700 ;
      RECT 1071.3600 2003.6200 1279.3800 2005.8200 ;
      RECT 1952.1000 2003.3600 2160.1200 2005.5600 ;
      RECT 3364.7200 2003.0800 3370.4200 2004.1600 ;
      RECT 3307.6200 2003.0800 3361.1200 2004.1600 ;
      RECT 2494.8200 2003.0800 3305.4200 2004.1600 ;
      RECT 2449.0800 2003.0800 2492.6200 2004.1600 ;
      RECT 2446.4800 2003.0800 2446.8800 2004.1600 ;
      RECT 1004.8200 2003.0800 1005.2200 2004.1600 ;
      RECT 967.6200 2003.0800 1002.6200 2004.1600 ;
      RECT 154.8200 2003.0800 965.4200 2004.1600 ;
      RECT 9.3000 2003.0800 152.6200 2004.1600 ;
      RECT 0.0000 2003.0800 5.7000 2004.1600 ;
      RECT 1065.1600 2002.6700 1283.0400 2003.6200 ;
      RECT 1011.2200 2002.6700 1059.1600 2004.8700 ;
      RECT 0.0000 2002.6700 1005.2200 2003.0800 ;
      RECT 2446.4800 2002.3100 3370.4200 2003.0800 ;
      RECT 2392.5400 2002.3100 2440.4800 2004.5100 ;
      RECT 2172.3200 2002.3100 2380.3400 2004.5100 ;
      RECT 1945.9000 2002.3100 2163.9200 2003.3600 ;
      RECT 1731.8800 2002.3100 1939.9000 2004.5100 ;
      RECT 1511.6600 2002.3100 1719.6800 2004.5100 ;
      RECT 1291.4400 2002.3100 1499.4600 2004.5100 ;
      RECT 0.0000 2002.3100 1283.0400 2002.6700 ;
      RECT 0.0000 2001.4400 3370.4200 2002.3100 ;
      RECT 3368.7200 2000.3600 3370.4200 2001.4400 ;
      RECT 3305.0200 2000.3600 3365.1200 2001.4400 ;
      RECT 2497.4200 2000.3600 3302.8200 2001.4400 ;
      RECT 2446.4800 2000.3600 2495.2200 2001.4400 ;
      RECT 1007.4200 2000.3600 2444.2800 2001.4400 ;
      RECT 965.0200 2000.3600 1005.2200 2001.4400 ;
      RECT 157.4200 2000.3600 962.8200 2001.4400 ;
      RECT 5.3000 2000.3600 155.2200 2001.4400 ;
      RECT 0.0000 2000.3600 1.7000 2001.4400 ;
      RECT 0.0000 1999.9000 3370.4200 2000.3600 ;
      RECT 1057.5000 1999.6400 3370.4200 1999.9000 ;
      RECT 1057.5000 1998.8200 1293.0000 1999.6400 ;
      RECT 0.0000 1998.8200 1055.3000 1999.9000 ;
      RECT 0.0000 1998.7400 1293.0000 1998.8200 ;
      RECT 2396.3000 1998.7200 3370.4200 1999.6400 ;
      RECT 0.0000 1998.7200 1072.9200 1998.7400 ;
      RECT 2396.3000 1998.5600 2446.8800 1998.7200 ;
      RECT 2176.0800 1998.5600 2394.1000 1999.6400 ;
      RECT 1735.6400 1998.5600 2173.8800 1999.6400 ;
      RECT 1515.4200 1998.5600 1733.4400 1999.6400 ;
      RECT 1295.2000 1998.5600 1513.2200 1999.6400 ;
      RECT 1075.1200 1998.5600 1293.0000 1998.7400 ;
      RECT 1075.1200 1998.4800 2446.8800 1998.5600 ;
      RECT 1075.1200 1997.6600 1953.6600 1998.4800 ;
      RECT 1004.8200 1997.6600 1072.9200 1998.7200 ;
      RECT 3364.7200 1997.6400 3370.4200 1998.7200 ;
      RECT 3307.6200 1997.6400 3361.1200 1998.7200 ;
      RECT 2494.8200 1997.6400 3305.4200 1998.7200 ;
      RECT 2449.0800 1997.6400 2492.6200 1998.7200 ;
      RECT 1955.8600 1997.6400 2446.8800 1998.4800 ;
      RECT 1004.8200 1997.6400 1953.6600 1997.6600 ;
      RECT 967.6200 1997.6400 1002.6200 1998.7200 ;
      RECT 154.8200 1997.6400 965.4200 1998.7200 ;
      RECT 9.3000 1997.6400 152.6200 1998.7200 ;
      RECT 0.0000 1997.6400 5.7000 1998.7200 ;
      RECT 1955.8600 1997.4000 3370.4200 1997.6400 ;
      RECT 0.0000 1997.4000 1953.6600 1997.6400 ;
      RECT 0.0000 1997.2500 3370.4200 1997.4000 ;
      RECT 1.1000 1996.3500 3370.4200 1997.2500 ;
      RECT 0.0000 1996.0000 3370.4200 1996.3500 ;
      RECT 3368.7200 1994.9200 3370.4200 1996.0000 ;
      RECT 3305.0200 1994.9200 3365.1200 1996.0000 ;
      RECT 2497.4200 1994.9200 3302.8200 1996.0000 ;
      RECT 2446.4800 1994.9200 2495.2200 1996.0000 ;
      RECT 1007.4200 1994.9200 2444.2800 1996.0000 ;
      RECT 965.0200 1994.9200 1005.2200 1996.0000 ;
      RECT 157.4200 1994.9200 962.8200 1996.0000 ;
      RECT 5.3000 1994.9200 155.2200 1996.0000 ;
      RECT 0.0000 1994.9200 1.7000 1996.0000 ;
      RECT 0.0000 1993.2800 3370.4200 1994.9200 ;
      RECT 3364.7200 1992.2000 3370.4200 1993.2800 ;
      RECT 3307.6200 1992.2000 3361.1200 1993.2800 ;
      RECT 2494.8200 1992.2000 3305.4200 1993.2800 ;
      RECT 2449.0800 1992.2000 2492.6200 1993.2800 ;
      RECT 1004.8200 1992.2000 2446.8800 1993.2800 ;
      RECT 967.6200 1992.2000 1002.6200 1993.2800 ;
      RECT 154.8200 1992.2000 965.4200 1993.2800 ;
      RECT 9.3000 1992.2000 152.6200 1993.2800 ;
      RECT 0.0000 1992.2000 5.7000 1993.2800 ;
      RECT 0.0000 1990.5600 3370.4200 1992.2000 ;
      RECT 3368.7200 1989.4800 3370.4200 1990.5600 ;
      RECT 3305.0200 1989.4800 3365.1200 1990.5600 ;
      RECT 2497.4200 1989.4800 3302.8200 1990.5600 ;
      RECT 2446.4800 1989.4800 2495.2200 1990.5600 ;
      RECT 1007.4200 1989.4800 2444.2800 1990.5600 ;
      RECT 965.0200 1989.4800 1005.2200 1990.5600 ;
      RECT 157.4200 1989.4800 962.8200 1990.5600 ;
      RECT 5.3000 1989.4800 155.2200 1990.5600 ;
      RECT 0.0000 1989.4800 1.7000 1990.5600 ;
      RECT 0.0000 1987.8400 3370.4200 1989.4800 ;
      RECT 0.0000 1986.8800 5.7000 1987.8400 ;
      RECT 3364.7200 1986.7600 3370.4200 1987.8400 ;
      RECT 3307.6200 1986.7600 3361.1200 1987.8400 ;
      RECT 2494.8200 1986.7600 3305.4200 1987.8400 ;
      RECT 2449.0800 1986.7600 2492.6200 1987.8400 ;
      RECT 1004.8200 1986.7600 2446.8800 1987.8400 ;
      RECT 967.6200 1986.7600 1002.6200 1987.8400 ;
      RECT 154.8200 1986.7600 965.4200 1987.8400 ;
      RECT 9.3000 1986.7600 152.6200 1987.8400 ;
      RECT 1.1000 1986.7600 5.7000 1986.8800 ;
      RECT 1.1000 1985.9800 3370.4200 1986.7600 ;
      RECT 0.0000 1985.1200 3370.4200 1985.9800 ;
      RECT 3368.7200 1984.0400 3370.4200 1985.1200 ;
      RECT 3305.0200 1984.0400 3365.1200 1985.1200 ;
      RECT 2497.4200 1984.0400 3302.8200 1985.1200 ;
      RECT 2446.4800 1984.0400 2495.2200 1985.1200 ;
      RECT 1007.4200 1984.0400 2444.2800 1985.1200 ;
      RECT 965.0200 1984.0400 1005.2200 1985.1200 ;
      RECT 157.4200 1984.0400 962.8200 1985.1200 ;
      RECT 5.3000 1984.0400 155.2200 1985.1200 ;
      RECT 0.0000 1984.0400 1.7000 1985.1200 ;
      RECT 0.0000 1982.4000 3370.4200 1984.0400 ;
      RECT 3364.7200 1981.3200 3370.4200 1982.4000 ;
      RECT 3307.6200 1981.3200 3361.1200 1982.4000 ;
      RECT 2494.8200 1981.3200 3305.4200 1982.4000 ;
      RECT 2449.0800 1981.3200 2492.6200 1982.4000 ;
      RECT 1004.8200 1981.3200 2446.8800 1982.4000 ;
      RECT 967.6200 1981.3200 1002.6200 1982.4000 ;
      RECT 154.8200 1981.3200 965.4200 1982.4000 ;
      RECT 9.3000 1981.3200 152.6200 1982.4000 ;
      RECT 0.0000 1981.3200 5.7000 1982.4000 ;
      RECT 0.0000 1979.6800 3370.4200 1981.3200 ;
      RECT 3368.7200 1978.6000 3370.4200 1979.6800 ;
      RECT 3305.0200 1978.6000 3365.1200 1979.6800 ;
      RECT 2497.4200 1978.6000 3302.8200 1979.6800 ;
      RECT 2446.4800 1978.6000 2495.2200 1979.6800 ;
      RECT 1007.4200 1978.6000 2444.2800 1979.6800 ;
      RECT 965.0200 1978.6000 1005.2200 1979.6800 ;
      RECT 157.4200 1978.6000 962.8200 1979.6800 ;
      RECT 5.3000 1978.6000 155.2200 1979.6800 ;
      RECT 0.0000 1978.6000 1.7000 1979.6800 ;
      RECT 0.0000 1976.9600 3370.4200 1978.6000 ;
      RECT 0.0000 1975.9000 5.7000 1976.9600 ;
      RECT 3364.7200 1975.8800 3370.4200 1976.9600 ;
      RECT 3307.6200 1975.8800 3361.1200 1976.9600 ;
      RECT 2494.8200 1975.8800 3305.4200 1976.9600 ;
      RECT 2449.0800 1975.8800 2492.6200 1976.9600 ;
      RECT 1004.8200 1975.8800 2446.8800 1976.9600 ;
      RECT 967.6200 1975.8800 1002.6200 1976.9600 ;
      RECT 154.8200 1975.8800 965.4200 1976.9600 ;
      RECT 9.3000 1975.8800 152.6200 1976.9600 ;
      RECT 1.1000 1975.8800 5.7000 1975.9000 ;
      RECT 1.1000 1975.0000 3370.4200 1975.8800 ;
      RECT 0.0000 1974.2400 3370.4200 1975.0000 ;
      RECT 3368.7200 1973.1600 3370.4200 1974.2400 ;
      RECT 3305.0200 1973.1600 3365.1200 1974.2400 ;
      RECT 2497.4200 1973.1600 3302.8200 1974.2400 ;
      RECT 2446.4800 1973.1600 2495.2200 1974.2400 ;
      RECT 1007.4200 1973.1600 2444.2800 1974.2400 ;
      RECT 965.0200 1973.1600 1005.2200 1974.2400 ;
      RECT 157.4200 1973.1600 962.8200 1974.2400 ;
      RECT 5.3000 1973.1600 155.2200 1974.2400 ;
      RECT 0.0000 1973.1600 1.7000 1974.2400 ;
      RECT 0.0000 1971.5200 3370.4200 1973.1600 ;
      RECT 3364.7200 1970.4400 3370.4200 1971.5200 ;
      RECT 3307.6200 1970.4400 3361.1200 1971.5200 ;
      RECT 2494.8200 1970.4400 3305.4200 1971.5200 ;
      RECT 2449.0800 1970.4400 2492.6200 1971.5200 ;
      RECT 1004.8200 1970.4400 2446.8800 1971.5200 ;
      RECT 967.6200 1970.4400 1002.6200 1971.5200 ;
      RECT 154.8200 1970.4400 965.4200 1971.5200 ;
      RECT 9.3000 1970.4400 152.6200 1971.5200 ;
      RECT 0.0000 1970.4400 5.7000 1971.5200 ;
      RECT 0.0000 1968.8000 3370.4200 1970.4400 ;
      RECT 3368.7200 1967.7200 3370.4200 1968.8000 ;
      RECT 3305.0200 1967.7200 3365.1200 1968.8000 ;
      RECT 157.4200 1967.7200 3302.8200 1968.8000 ;
      RECT 5.3000 1967.7200 155.2200 1968.8000 ;
      RECT 0.0000 1967.7200 1.7000 1968.8000 ;
      RECT 0.0000 1966.0800 3370.4200 1967.7200 ;
      RECT 3364.7200 1965.0000 3370.4200 1966.0800 ;
      RECT 3307.6200 1965.0000 3361.1200 1966.0800 ;
      RECT 154.8200 1965.0000 3305.4200 1966.0800 ;
      RECT 9.3000 1965.0000 152.6200 1966.0800 ;
      RECT 0.0000 1965.0000 5.7000 1966.0800 ;
      RECT 0.0000 1964.9200 3370.4200 1965.0000 ;
      RECT 1.1000 1964.0200 3370.4200 1964.9200 ;
      RECT 0.0000 1963.3600 3370.4200 1964.0200 ;
      RECT 3368.7200 1962.2800 3370.4200 1963.3600 ;
      RECT 3305.0200 1962.2800 3365.1200 1963.3600 ;
      RECT 157.4200 1962.2800 3302.8200 1963.3600 ;
      RECT 5.3000 1962.2800 155.2200 1963.3600 ;
      RECT 0.0000 1962.2800 1.7000 1963.3600 ;
      RECT 0.0000 1960.6400 3370.4200 1962.2800 ;
      RECT 3364.7200 1959.5600 3370.4200 1960.6400 ;
      RECT 3307.6200 1959.5600 3361.1200 1960.6400 ;
      RECT 154.8200 1959.5600 3305.4200 1960.6400 ;
      RECT 9.3000 1959.5600 152.6200 1960.6400 ;
      RECT 0.0000 1959.5600 5.7000 1960.6400 ;
      RECT 0.0000 1957.9200 3370.4200 1959.5600 ;
      RECT 3368.7200 1956.8400 3370.4200 1957.9200 ;
      RECT 3305.0200 1956.8400 3365.1200 1957.9200 ;
      RECT 157.4200 1956.8400 3302.8200 1957.9200 ;
      RECT 5.3000 1956.8400 155.2200 1957.9200 ;
      RECT 0.0000 1956.8400 1.7000 1957.9200 ;
      RECT 0.0000 1955.2000 3370.4200 1956.8400 ;
      RECT 3364.7200 1954.1200 3370.4200 1955.2000 ;
      RECT 3307.6200 1954.1200 3361.1200 1955.2000 ;
      RECT 154.8200 1954.1200 3305.4200 1955.2000 ;
      RECT 9.3000 1954.1200 152.6200 1955.2000 ;
      RECT 0.0000 1954.1200 5.7000 1955.2000 ;
      RECT 0.0000 1953.9400 3370.4200 1954.1200 ;
      RECT 1.1000 1953.0400 3370.4200 1953.9400 ;
      RECT 0.0000 1952.4800 3370.4200 1953.0400 ;
      RECT 3368.7200 1951.4000 3370.4200 1952.4800 ;
      RECT 3305.0200 1951.4000 3365.1200 1952.4800 ;
      RECT 157.4200 1951.4000 3302.8200 1952.4800 ;
      RECT 5.3000 1951.4000 155.2200 1952.4800 ;
      RECT 0.0000 1951.4000 1.7000 1952.4800 ;
      RECT 0.0000 1949.7600 3370.4200 1951.4000 ;
      RECT 3364.7200 1948.6800 3370.4200 1949.7600 ;
      RECT 3307.6200 1948.6800 3361.1200 1949.7600 ;
      RECT 154.8200 1948.6800 3305.4200 1949.7600 ;
      RECT 9.3000 1948.6800 152.6200 1949.7600 ;
      RECT 0.0000 1948.6800 5.7000 1949.7600 ;
      RECT 0.0000 1947.0400 3370.4200 1948.6800 ;
      RECT 3368.7200 1945.9600 3370.4200 1947.0400 ;
      RECT 3305.0200 1945.9600 3365.1200 1947.0400 ;
      RECT 157.4200 1945.9600 3302.8200 1947.0400 ;
      RECT 5.3000 1945.9600 155.2200 1947.0400 ;
      RECT 0.0000 1945.9600 1.7000 1947.0400 ;
      RECT 0.0000 1944.3200 3370.4200 1945.9600 ;
      RECT 3364.7200 1943.2400 3370.4200 1944.3200 ;
      RECT 3307.6200 1943.2400 3361.1200 1944.3200 ;
      RECT 154.8200 1943.2400 3305.4200 1944.3200 ;
      RECT 9.3000 1943.2400 152.6200 1944.3200 ;
      RECT 0.0000 1943.2400 5.7000 1944.3200 ;
      RECT 0.0000 1942.9600 3370.4200 1943.2400 ;
      RECT 1.1000 1942.0600 3370.4200 1942.9600 ;
      RECT 0.0000 1941.6000 3370.4200 1942.0600 ;
      RECT 3368.7200 1940.5200 3370.4200 1941.6000 ;
      RECT 3305.0200 1940.5200 3365.1200 1941.6000 ;
      RECT 157.4200 1940.5200 3302.8200 1941.6000 ;
      RECT 5.3000 1940.5200 155.2200 1941.6000 ;
      RECT 0.0000 1940.5200 1.7000 1941.6000 ;
      RECT 0.0000 1938.8800 3370.4200 1940.5200 ;
      RECT 3364.7200 1937.8000 3370.4200 1938.8800 ;
      RECT 3307.6200 1937.8000 3361.1200 1938.8800 ;
      RECT 154.8200 1937.8000 3305.4200 1938.8800 ;
      RECT 9.3000 1937.8000 152.6200 1938.8800 ;
      RECT 0.0000 1937.8000 5.7000 1938.8800 ;
      RECT 0.0000 1936.1600 3370.4200 1937.8000 ;
      RECT 3368.7200 1935.0800 3370.4200 1936.1600 ;
      RECT 3305.0200 1935.0800 3365.1200 1936.1600 ;
      RECT 157.4200 1935.0800 3302.8200 1936.1600 ;
      RECT 5.3000 1935.0800 155.2200 1936.1600 ;
      RECT 0.0000 1935.0800 1.7000 1936.1600 ;
      RECT 0.0000 1933.4400 3370.4200 1935.0800 ;
      RECT 0.0000 1932.5900 5.7000 1933.4400 ;
      RECT 3364.7200 1932.3600 3370.4200 1933.4400 ;
      RECT 3307.6200 1932.3600 3361.1200 1933.4400 ;
      RECT 154.8200 1932.3600 3305.4200 1933.4400 ;
      RECT 9.3000 1932.3600 152.6200 1933.4400 ;
      RECT 1.1000 1932.3600 5.7000 1932.5900 ;
      RECT 1.1000 1931.6900 3370.4200 1932.3600 ;
      RECT 0.0000 1930.7200 3370.4200 1931.6900 ;
      RECT 3368.7200 1929.6400 3370.4200 1930.7200 ;
      RECT 3305.0200 1929.6400 3365.1200 1930.7200 ;
      RECT 157.4200 1929.6400 3302.8200 1930.7200 ;
      RECT 5.3000 1929.6400 155.2200 1930.7200 ;
      RECT 0.0000 1929.6400 1.7000 1930.7200 ;
      RECT 0.0000 1928.0000 3370.4200 1929.6400 ;
      RECT 3364.7200 1926.9200 3370.4200 1928.0000 ;
      RECT 3307.6200 1926.9200 3361.1200 1928.0000 ;
      RECT 154.8200 1926.9200 3305.4200 1928.0000 ;
      RECT 9.3000 1926.9200 152.6200 1928.0000 ;
      RECT 0.0000 1926.9200 5.7000 1928.0000 ;
      RECT 0.0000 1925.2800 3370.4200 1926.9200 ;
      RECT 3368.7200 1924.2000 3370.4200 1925.2800 ;
      RECT 3305.0200 1924.2000 3365.1200 1925.2800 ;
      RECT 157.4200 1924.2000 3302.8200 1925.2800 ;
      RECT 5.3000 1924.2000 155.2200 1925.2800 ;
      RECT 0.0000 1924.2000 1.7000 1925.2800 ;
      RECT 0.0000 1922.5600 3370.4200 1924.2000 ;
      RECT 0.0000 1921.6100 5.7000 1922.5600 ;
      RECT 3364.7200 1921.4800 3370.4200 1922.5600 ;
      RECT 3307.6200 1921.4800 3361.1200 1922.5600 ;
      RECT 154.8200 1921.4800 3305.4200 1922.5600 ;
      RECT 9.3000 1921.4800 152.6200 1922.5600 ;
      RECT 1.1000 1921.4800 5.7000 1921.6100 ;
      RECT 1.1000 1920.7100 3370.4200 1921.4800 ;
      RECT 0.0000 1919.8400 3370.4200 1920.7100 ;
      RECT 3368.7200 1918.7600 3370.4200 1919.8400 ;
      RECT 3305.0200 1918.7600 3365.1200 1919.8400 ;
      RECT 157.4200 1918.7600 3302.8200 1919.8400 ;
      RECT 5.3000 1918.7600 155.2200 1919.8400 ;
      RECT 0.0000 1918.7600 1.7000 1919.8400 ;
      RECT 0.0000 1917.1200 3370.4200 1918.7600 ;
      RECT 3364.7200 1916.0400 3370.4200 1917.1200 ;
      RECT 3307.6200 1916.0400 3361.1200 1917.1200 ;
      RECT 154.8200 1916.0400 3305.4200 1917.1200 ;
      RECT 9.3000 1916.0400 152.6200 1917.1200 ;
      RECT 0.0000 1916.0400 5.7000 1917.1200 ;
      RECT 0.0000 1914.4000 3370.4200 1916.0400 ;
      RECT 3368.7200 1913.3200 3370.4200 1914.4000 ;
      RECT 3305.0200 1913.3200 3365.1200 1914.4000 ;
      RECT 157.4200 1913.3200 3302.8200 1914.4000 ;
      RECT 5.3000 1913.3200 155.2200 1914.4000 ;
      RECT 0.0000 1913.3200 1.7000 1914.4000 ;
      RECT 0.0000 1911.6800 3370.4200 1913.3200 ;
      RECT 0.0000 1910.6300 5.7000 1911.6800 ;
      RECT 3364.7200 1910.6000 3370.4200 1911.6800 ;
      RECT 3307.6200 1910.6000 3361.1200 1911.6800 ;
      RECT 154.8200 1910.6000 3305.4200 1911.6800 ;
      RECT 9.3000 1910.6000 152.6200 1911.6800 ;
      RECT 1.1000 1910.6000 5.7000 1910.6300 ;
      RECT 1.1000 1909.7300 3370.4200 1910.6000 ;
      RECT 0.0000 1908.9600 3370.4200 1909.7300 ;
      RECT 3368.7200 1907.8800 3370.4200 1908.9600 ;
      RECT 3305.0200 1907.8800 3365.1200 1908.9600 ;
      RECT 157.4200 1907.8800 3302.8200 1908.9600 ;
      RECT 5.3000 1907.8800 155.2200 1908.9600 ;
      RECT 0.0000 1907.8800 1.7000 1908.9600 ;
      RECT 0.0000 1906.2400 3370.4200 1907.8800 ;
      RECT 3364.7200 1905.1600 3370.4200 1906.2400 ;
      RECT 3307.6200 1905.1600 3361.1200 1906.2400 ;
      RECT 154.8200 1905.1600 3305.4200 1906.2400 ;
      RECT 9.3000 1905.1600 152.6200 1906.2400 ;
      RECT 0.0000 1905.1600 5.7000 1906.2400 ;
      RECT 0.0000 1903.5200 3370.4200 1905.1600 ;
      RECT 3368.7200 1902.4400 3370.4200 1903.5200 ;
      RECT 3305.0200 1902.4400 3365.1200 1903.5200 ;
      RECT 157.4200 1902.4400 3302.8200 1903.5200 ;
      RECT 5.3000 1902.4400 155.2200 1903.5200 ;
      RECT 0.0000 1902.4400 1.7000 1903.5200 ;
      RECT 0.0000 1900.8000 3370.4200 1902.4400 ;
      RECT 3364.7200 1899.7200 3370.4200 1900.8000 ;
      RECT 3307.6200 1899.7200 3361.1200 1900.8000 ;
      RECT 154.8200 1899.7200 3305.4200 1900.8000 ;
      RECT 9.3000 1899.7200 152.6200 1900.8000 ;
      RECT 0.0000 1899.7200 5.7000 1900.8000 ;
      RECT 0.0000 1899.6500 3370.4200 1899.7200 ;
      RECT 1.1000 1898.7500 3370.4200 1899.6500 ;
      RECT 0.0000 1898.0800 3370.4200 1898.7500 ;
      RECT 3368.7200 1897.0000 3370.4200 1898.0800 ;
      RECT 3305.0200 1897.0000 3365.1200 1898.0800 ;
      RECT 157.4200 1897.0000 3302.8200 1898.0800 ;
      RECT 5.3000 1897.0000 155.2200 1898.0800 ;
      RECT 0.0000 1897.0000 1.7000 1898.0800 ;
      RECT 0.0000 1895.3600 3370.4200 1897.0000 ;
      RECT 3364.7200 1894.2800 3370.4200 1895.3600 ;
      RECT 3307.6200 1894.2800 3361.1200 1895.3600 ;
      RECT 154.8200 1894.2800 3305.4200 1895.3600 ;
      RECT 9.3000 1894.2800 152.6200 1895.3600 ;
      RECT 0.0000 1894.2800 5.7000 1895.3600 ;
      RECT 0.0000 1892.6400 3370.4200 1894.2800 ;
      RECT 3368.7200 1891.5600 3370.4200 1892.6400 ;
      RECT 3305.0200 1891.5600 3365.1200 1892.6400 ;
      RECT 157.4200 1891.5600 3302.8200 1892.6400 ;
      RECT 5.3000 1891.5600 155.2200 1892.6400 ;
      RECT 0.0000 1891.5600 1.7000 1892.6400 ;
      RECT 0.0000 1889.9200 3370.4200 1891.5600 ;
      RECT 3364.7200 1888.8400 3370.4200 1889.9200 ;
      RECT 3307.6200 1888.8400 3361.1200 1889.9200 ;
      RECT 154.8200 1888.8400 3305.4200 1889.9200 ;
      RECT 9.3000 1888.8400 152.6200 1889.9200 ;
      RECT 0.0000 1888.8400 5.7000 1889.9200 ;
      RECT 0.0000 1888.6700 3370.4200 1888.8400 ;
      RECT 1.1000 1887.7700 3370.4200 1888.6700 ;
      RECT 0.0000 1887.2000 3370.4200 1887.7700 ;
      RECT 3368.7200 1886.1200 3370.4200 1887.2000 ;
      RECT 3305.0200 1886.1200 3365.1200 1887.2000 ;
      RECT 157.4200 1886.1200 3302.8200 1887.2000 ;
      RECT 5.3000 1886.1200 155.2200 1887.2000 ;
      RECT 0.0000 1886.1200 1.7000 1887.2000 ;
      RECT 0.0000 1884.4800 3370.4200 1886.1200 ;
      RECT 3364.7200 1883.4000 3370.4200 1884.4800 ;
      RECT 3307.6200 1883.4000 3361.1200 1884.4800 ;
      RECT 154.8200 1883.4000 3305.4200 1884.4800 ;
      RECT 9.3000 1883.4000 152.6200 1884.4800 ;
      RECT 0.0000 1883.4000 5.7000 1884.4800 ;
      RECT 0.0000 1881.7600 3370.4200 1883.4000 ;
      RECT 3368.7200 1880.6800 3370.4200 1881.7600 ;
      RECT 3305.0200 1880.6800 3365.1200 1881.7600 ;
      RECT 157.4200 1880.6800 3302.8200 1881.7600 ;
      RECT 5.3000 1880.6800 155.2200 1881.7600 ;
      RECT 0.0000 1880.6800 1.7000 1881.7600 ;
      RECT 0.0000 1879.0400 3370.4200 1880.6800 ;
      RECT 0.0000 1878.3000 5.7000 1879.0400 ;
      RECT 3364.7200 1877.9600 3370.4200 1879.0400 ;
      RECT 3307.6200 1877.9600 3361.1200 1879.0400 ;
      RECT 154.8200 1877.9600 3305.4200 1879.0400 ;
      RECT 9.3000 1877.9600 152.6200 1879.0400 ;
      RECT 1.1000 1877.9600 5.7000 1878.3000 ;
      RECT 1.1000 1877.4000 3370.4200 1877.9600 ;
      RECT 0.0000 1876.3200 3370.4200 1877.4000 ;
      RECT 3368.7200 1875.2400 3370.4200 1876.3200 ;
      RECT 3305.0200 1875.2400 3365.1200 1876.3200 ;
      RECT 157.4200 1875.2400 3302.8200 1876.3200 ;
      RECT 5.3000 1875.2400 155.2200 1876.3200 ;
      RECT 0.0000 1875.2400 1.7000 1876.3200 ;
      RECT 0.0000 1873.6000 3370.4200 1875.2400 ;
      RECT 3364.7200 1872.5200 3370.4200 1873.6000 ;
      RECT 3307.6200 1872.5200 3361.1200 1873.6000 ;
      RECT 154.8200 1872.5200 3305.4200 1873.6000 ;
      RECT 9.3000 1872.5200 152.6200 1873.6000 ;
      RECT 0.0000 1872.5200 5.7000 1873.6000 ;
      RECT 0.0000 1870.8800 3370.4200 1872.5200 ;
      RECT 3368.7200 1869.8000 3370.4200 1870.8800 ;
      RECT 3305.0200 1869.8000 3365.1200 1870.8800 ;
      RECT 157.4200 1869.8000 3302.8200 1870.8800 ;
      RECT 5.3000 1869.8000 155.2200 1870.8800 ;
      RECT 0.0000 1869.8000 1.7000 1870.8800 ;
      RECT 0.0000 1868.1600 3370.4200 1869.8000 ;
      RECT 0.0000 1867.3200 5.7000 1868.1600 ;
      RECT 3364.7200 1867.0800 3370.4200 1868.1600 ;
      RECT 3307.6200 1867.0800 3361.1200 1868.1600 ;
      RECT 154.8200 1867.0800 3305.4200 1868.1600 ;
      RECT 9.3000 1867.0800 152.6200 1868.1600 ;
      RECT 1.1000 1867.0800 5.7000 1867.3200 ;
      RECT 1.1000 1866.4200 3370.4200 1867.0800 ;
      RECT 0.0000 1865.4400 3370.4200 1866.4200 ;
      RECT 3368.7200 1864.3600 3370.4200 1865.4400 ;
      RECT 3305.0200 1864.3600 3365.1200 1865.4400 ;
      RECT 157.4200 1864.3600 3302.8200 1865.4400 ;
      RECT 5.3000 1864.3600 155.2200 1865.4400 ;
      RECT 0.0000 1864.3600 1.7000 1865.4400 ;
      RECT 0.0000 1862.7200 3370.4200 1864.3600 ;
      RECT 3364.7200 1861.6400 3370.4200 1862.7200 ;
      RECT 3307.6200 1861.6400 3361.1200 1862.7200 ;
      RECT 154.8200 1861.6400 3305.4200 1862.7200 ;
      RECT 9.3000 1861.6400 152.6200 1862.7200 ;
      RECT 0.0000 1861.6400 5.7000 1862.7200 ;
      RECT 0.0000 1860.0000 3370.4200 1861.6400 ;
      RECT 3368.7200 1858.9200 3370.4200 1860.0000 ;
      RECT 3305.0200 1858.9200 3365.1200 1860.0000 ;
      RECT 157.4200 1858.9200 3302.8200 1860.0000 ;
      RECT 5.3000 1858.9200 155.2200 1860.0000 ;
      RECT 0.0000 1858.9200 1.7000 1860.0000 ;
      RECT 0.0000 1857.2800 3370.4200 1858.9200 ;
      RECT 0.0000 1856.3400 5.7000 1857.2800 ;
      RECT 3364.7200 1856.2000 3370.4200 1857.2800 ;
      RECT 3307.6200 1856.2000 3361.1200 1857.2800 ;
      RECT 154.8200 1856.2000 3305.4200 1857.2800 ;
      RECT 9.3000 1856.2000 152.6200 1857.2800 ;
      RECT 1.1000 1856.2000 5.7000 1856.3400 ;
      RECT 1.1000 1855.4400 3370.4200 1856.2000 ;
      RECT 0.0000 1854.5600 3370.4200 1855.4400 ;
      RECT 3368.7200 1853.4800 3370.4200 1854.5600 ;
      RECT 3305.0200 1853.4800 3365.1200 1854.5600 ;
      RECT 157.4200 1853.4800 3302.8200 1854.5600 ;
      RECT 5.3000 1853.4800 155.2200 1854.5600 ;
      RECT 0.0000 1853.4800 1.7000 1854.5600 ;
      RECT 0.0000 1851.8400 3370.4200 1853.4800 ;
      RECT 3364.7200 1850.7600 3370.4200 1851.8400 ;
      RECT 3307.6200 1850.7600 3361.1200 1851.8400 ;
      RECT 154.8200 1850.7600 3305.4200 1851.8400 ;
      RECT 9.3000 1850.7600 152.6200 1851.8400 ;
      RECT 0.0000 1850.7600 5.7000 1851.8400 ;
      RECT 0.0000 1849.1200 3370.4200 1850.7600 ;
      RECT 3368.7200 1848.0400 3370.4200 1849.1200 ;
      RECT 3305.0200 1848.0400 3365.1200 1849.1200 ;
      RECT 157.4200 1848.0400 3302.8200 1849.1200 ;
      RECT 5.3000 1848.0400 155.2200 1849.1200 ;
      RECT 0.0000 1848.0400 1.7000 1849.1200 ;
      RECT 0.0000 1846.4000 3370.4200 1848.0400 ;
      RECT 0.0000 1845.3600 5.7000 1846.4000 ;
      RECT 3364.7200 1845.3200 3370.4200 1846.4000 ;
      RECT 3307.6200 1845.3200 3361.1200 1846.4000 ;
      RECT 154.8200 1845.3200 3305.4200 1846.4000 ;
      RECT 9.3000 1845.3200 152.6200 1846.4000 ;
      RECT 1.1000 1845.3200 5.7000 1845.3600 ;
      RECT 1.1000 1844.4600 3370.4200 1845.3200 ;
      RECT 0.0000 1843.6800 3370.4200 1844.4600 ;
      RECT 3368.7200 1842.6000 3370.4200 1843.6800 ;
      RECT 3305.0200 1842.6000 3365.1200 1843.6800 ;
      RECT 157.4200 1842.6000 3302.8200 1843.6800 ;
      RECT 5.3000 1842.6000 155.2200 1843.6800 ;
      RECT 0.0000 1842.6000 1.7000 1843.6800 ;
      RECT 0.0000 1840.9600 3370.4200 1842.6000 ;
      RECT 3364.7200 1839.8800 3370.4200 1840.9600 ;
      RECT 3307.6200 1839.8800 3361.1200 1840.9600 ;
      RECT 154.8200 1839.8800 3305.4200 1840.9600 ;
      RECT 9.3000 1839.8800 152.6200 1840.9600 ;
      RECT 0.0000 1839.8800 5.7000 1840.9600 ;
      RECT 0.0000 1838.2400 3370.4200 1839.8800 ;
      RECT 3368.7200 1837.1600 3370.4200 1838.2400 ;
      RECT 3305.0200 1837.1600 3365.1200 1838.2400 ;
      RECT 157.4200 1837.1600 3302.8200 1838.2400 ;
      RECT 5.3000 1837.1600 155.2200 1838.2400 ;
      RECT 0.0000 1837.1600 1.7000 1838.2400 ;
      RECT 0.0000 1835.5200 3370.4200 1837.1600 ;
      RECT 3364.7200 1834.4400 3370.4200 1835.5200 ;
      RECT 3307.6200 1834.4400 3361.1200 1835.5200 ;
      RECT 154.8200 1834.4400 3305.4200 1835.5200 ;
      RECT 9.3000 1834.4400 152.6200 1835.5200 ;
      RECT 0.0000 1834.4400 5.7000 1835.5200 ;
      RECT 0.0000 1834.3800 3370.4200 1834.4400 ;
      RECT 1.1000 1833.4800 3370.4200 1834.3800 ;
      RECT 0.0000 1832.8000 3370.4200 1833.4800 ;
      RECT 3368.7200 1831.7200 3370.4200 1832.8000 ;
      RECT 3305.0200 1831.7200 3365.1200 1832.8000 ;
      RECT 157.4200 1831.7200 3302.8200 1832.8000 ;
      RECT 5.3000 1831.7200 155.2200 1832.8000 ;
      RECT 0.0000 1831.7200 1.7000 1832.8000 ;
      RECT 0.0000 1830.0800 3370.4200 1831.7200 ;
      RECT 3364.7200 1829.0000 3370.4200 1830.0800 ;
      RECT 3307.6200 1829.0000 3361.1200 1830.0800 ;
      RECT 154.8200 1829.0000 3305.4200 1830.0800 ;
      RECT 9.3000 1829.0000 152.6200 1830.0800 ;
      RECT 0.0000 1829.0000 5.7000 1830.0800 ;
      RECT 0.0000 1827.3600 3370.4200 1829.0000 ;
      RECT 3368.7200 1826.2800 3370.4200 1827.3600 ;
      RECT 3305.0200 1826.2800 3365.1200 1827.3600 ;
      RECT 157.4200 1826.2800 3302.8200 1827.3600 ;
      RECT 5.3000 1826.2800 155.2200 1827.3600 ;
      RECT 0.0000 1826.2800 1.7000 1827.3600 ;
      RECT 0.0000 1824.6400 3370.4200 1826.2800 ;
      RECT 0.0000 1824.0100 5.7000 1824.6400 ;
      RECT 3364.7200 1823.5600 3370.4200 1824.6400 ;
      RECT 3307.6200 1823.5600 3361.1200 1824.6400 ;
      RECT 154.8200 1823.5600 3305.4200 1824.6400 ;
      RECT 9.3000 1823.5600 152.6200 1824.6400 ;
      RECT 1.1000 1823.5600 5.7000 1824.0100 ;
      RECT 1.1000 1823.1100 3370.4200 1823.5600 ;
      RECT 0.0000 1821.9200 3370.4200 1823.1100 ;
      RECT 3368.7200 1820.8400 3370.4200 1821.9200 ;
      RECT 3305.0200 1820.8400 3365.1200 1821.9200 ;
      RECT 157.4200 1820.8400 3302.8200 1821.9200 ;
      RECT 5.3000 1820.8400 155.2200 1821.9200 ;
      RECT 0.0000 1820.8400 1.7000 1821.9200 ;
      RECT 0.0000 1819.2000 3370.4200 1820.8400 ;
      RECT 3364.7200 1818.1200 3370.4200 1819.2000 ;
      RECT 3307.6200 1818.1200 3361.1200 1819.2000 ;
      RECT 154.8200 1818.1200 3305.4200 1819.2000 ;
      RECT 9.3000 1818.1200 152.6200 1819.2000 ;
      RECT 0.0000 1818.1200 5.7000 1819.2000 ;
      RECT 0.0000 1816.4800 3370.4200 1818.1200 ;
      RECT 3368.7200 1815.4000 3370.4200 1816.4800 ;
      RECT 3305.0200 1815.4000 3365.1200 1816.4800 ;
      RECT 157.4200 1815.4000 3302.8200 1816.4800 ;
      RECT 5.3000 1815.4000 155.2200 1816.4800 ;
      RECT 0.0000 1815.4000 1.7000 1816.4800 ;
      RECT 0.0000 1813.7600 3370.4200 1815.4000 ;
      RECT 0.0000 1813.0300 5.7000 1813.7600 ;
      RECT 3364.7200 1812.6800 3370.4200 1813.7600 ;
      RECT 3307.6200 1812.6800 3361.1200 1813.7600 ;
      RECT 154.8200 1812.6800 3305.4200 1813.7600 ;
      RECT 9.3000 1812.6800 152.6200 1813.7600 ;
      RECT 1.1000 1812.6800 5.7000 1813.0300 ;
      RECT 1.1000 1812.1300 3370.4200 1812.6800 ;
      RECT 0.0000 1811.0400 3370.4200 1812.1300 ;
      RECT 3368.7200 1809.9600 3370.4200 1811.0400 ;
      RECT 3305.0200 1809.9600 3365.1200 1811.0400 ;
      RECT 157.4200 1809.9600 3302.8200 1811.0400 ;
      RECT 5.3000 1809.9600 155.2200 1811.0400 ;
      RECT 0.0000 1809.9600 1.7000 1811.0400 ;
      RECT 0.0000 1808.3200 3370.4200 1809.9600 ;
      RECT 3364.7200 1807.2400 3370.4200 1808.3200 ;
      RECT 3307.6200 1807.2400 3361.1200 1808.3200 ;
      RECT 154.8200 1807.2400 3305.4200 1808.3200 ;
      RECT 9.3000 1807.2400 152.6200 1808.3200 ;
      RECT 0.0000 1807.2400 5.7000 1808.3200 ;
      RECT 0.0000 1805.6000 3370.4200 1807.2400 ;
      RECT 3368.7200 1804.5200 3370.4200 1805.6000 ;
      RECT 3305.0200 1804.5200 3365.1200 1805.6000 ;
      RECT 157.4200 1804.5200 3302.8200 1805.6000 ;
      RECT 5.3000 1804.5200 155.2200 1805.6000 ;
      RECT 0.0000 1804.5200 1.7000 1805.6000 ;
      RECT 0.0000 1802.8800 3370.4200 1804.5200 ;
      RECT 0.0000 1802.0500 5.7000 1802.8800 ;
      RECT 3364.7200 1801.8000 3370.4200 1802.8800 ;
      RECT 3307.6200 1801.8000 3361.1200 1802.8800 ;
      RECT 154.8200 1801.8000 3305.4200 1802.8800 ;
      RECT 9.3000 1801.8000 152.6200 1802.8800 ;
      RECT 1.1000 1801.8000 5.7000 1802.0500 ;
      RECT 1.1000 1801.3400 3370.4200 1801.8000 ;
      RECT 1.1000 1801.1500 1015.2800 1801.3400 ;
      RECT 1017.4800 1801.0800 3370.4200 1801.3400 ;
      RECT 1017.4800 1800.2600 1295.6000 1801.0800 ;
      RECT 0.0000 1800.2600 1015.2800 1801.1500 ;
      RECT 2436.3200 1800.1600 3370.4200 1801.0800 ;
      RECT 0.0000 1800.1600 1295.6000 1800.2600 ;
      RECT 2436.3200 1800.0000 3302.8200 1800.1600 ;
      RECT 2178.6800 1800.0000 2434.1200 1801.0800 ;
      RECT 1738.2400 1800.0000 2176.4800 1801.0800 ;
      RECT 1518.0200 1800.0000 1736.0400 1801.0800 ;
      RECT 1297.8000 1800.0000 1515.8200 1801.0800 ;
      RECT 157.4200 1800.0000 1295.6000 1800.1600 ;
      RECT 3368.7200 1799.0800 3370.4200 1800.1600 ;
      RECT 3305.0200 1799.0800 3365.1200 1800.1600 ;
      RECT 157.4200 1799.0800 3302.8200 1800.0000 ;
      RECT 5.3000 1799.0800 155.2200 1800.1600 ;
      RECT 0.0000 1799.0800 1.7000 1800.1600 ;
      RECT 0.0000 1798.1700 3370.4200 1799.0800 ;
      RECT 1065.1600 1798.0100 3370.4200 1798.1700 ;
      RECT 2446.4800 1797.4400 3370.4200 1798.0100 ;
      RECT 0.0000 1797.4400 1005.2200 1798.1700 ;
      RECT 3364.7200 1796.3600 3370.4200 1797.4400 ;
      RECT 3307.6200 1796.3600 3361.1200 1797.4400 ;
      RECT 2446.4800 1796.3600 3305.4200 1797.4400 ;
      RECT 154.8200 1796.3600 1005.2200 1797.4400 ;
      RECT 9.3000 1796.3600 152.6200 1797.4400 ;
      RECT 0.0000 1796.3600 5.7000 1797.4400 ;
      RECT 1065.1600 1795.9700 1283.0400 1798.0100 ;
      RECT 1011.2200 1795.9700 1059.1600 1798.1700 ;
      RECT 0.0000 1795.9700 1005.2200 1796.3600 ;
      RECT 2446.4800 1795.8100 3370.4200 1796.3600 ;
      RECT 2392.5400 1795.8100 2440.4800 1798.0100 ;
      RECT 2172.3200 1795.8100 2380.3400 1798.0100 ;
      RECT 1945.9000 1795.8100 2163.9200 1798.0100 ;
      RECT 1731.8800 1795.8100 1939.9000 1798.0100 ;
      RECT 1511.6600 1795.8100 1719.6800 1798.0100 ;
      RECT 1291.4400 1795.8100 1499.4600 1798.0100 ;
      RECT 0.0000 1795.8100 1283.0400 1795.9700 ;
      RECT 0.0000 1795.7700 3370.4200 1795.8100 ;
      RECT 1067.7600 1795.4100 3370.4200 1795.7700 ;
      RECT 2449.0800 1794.7200 3370.4200 1795.4100 ;
      RECT 0.0000 1794.7200 1002.6200 1795.7700 ;
      RECT 3368.7200 1793.6400 3370.4200 1794.7200 ;
      RECT 3305.0200 1793.6400 3365.1200 1794.7200 ;
      RECT 2449.0800 1793.6400 3302.8200 1794.7200 ;
      RECT 157.4200 1793.6400 1002.6200 1794.7200 ;
      RECT 5.3000 1793.6400 155.2200 1794.7200 ;
      RECT 0.0000 1793.6400 1.7000 1794.7200 ;
      RECT 1067.7600 1793.5700 1285.6400 1795.4100 ;
      RECT 1011.2200 1793.5700 1059.1600 1795.7700 ;
      RECT 0.0000 1793.5700 1002.6200 1793.6400 ;
      RECT 2449.0800 1793.2100 3370.4200 1793.6400 ;
      RECT 2392.5400 1793.2100 2440.4800 1795.4100 ;
      RECT 2172.3200 1793.2100 2386.7400 1795.4100 ;
      RECT 1948.5000 1793.2100 2166.5200 1795.4100 ;
      RECT 1731.8800 1793.2100 1939.9000 1795.4100 ;
      RECT 1511.6600 1793.2100 1719.6800 1795.4100 ;
      RECT 1291.4400 1793.2100 1499.4600 1795.4100 ;
      RECT 0.0000 1793.2100 1285.6400 1793.5700 ;
      RECT 0.0000 1792.0000 3370.4200 1793.2100 ;
      RECT 0.0000 1791.0700 5.7000 1792.0000 ;
      RECT 3364.7200 1790.9200 3370.4200 1792.0000 ;
      RECT 3307.6200 1790.9200 3361.1200 1792.0000 ;
      RECT 154.8200 1790.9200 3305.4200 1792.0000 ;
      RECT 9.3000 1790.9200 152.6200 1792.0000 ;
      RECT 1.1000 1790.9200 5.7000 1791.0700 ;
      RECT 1.1000 1790.1700 3370.4200 1790.9200 ;
      RECT 0.0000 1789.2800 3370.4200 1790.1700 ;
      RECT 157.4200 1788.2400 3302.8200 1789.2800 ;
      RECT 5.3000 1788.2400 155.2200 1789.2800 ;
      RECT 3368.7200 1788.2000 3370.4200 1789.2800 ;
      RECT 3305.0200 1788.2000 3365.1200 1789.2800 ;
      RECT 1065.1600 1788.2000 3302.8200 1788.2400 ;
      RECT 1065.1600 1787.9800 3370.4200 1788.2000 ;
      RECT 2446.4800 1786.5600 3370.4200 1787.9800 ;
      RECT 1065.1600 1786.0400 1283.0400 1787.9800 ;
      RECT 167.4150 1786.0400 953.1450 1788.2400 ;
      RECT 0.0000 1786.0400 1.7000 1789.2800 ;
      RECT 2446.4800 1785.7800 3305.4200 1786.5600 ;
      RECT 1945.9000 1785.7800 2163.9200 1787.9800 ;
      RECT 154.8200 1785.7800 1283.0400 1786.0400 ;
      RECT 154.8200 1785.6400 3305.4200 1785.7800 ;
      RECT 9.3000 1785.6400 152.6200 1786.0400 ;
      RECT 3364.7200 1785.4800 3370.4200 1786.5600 ;
      RECT 3307.6200 1785.4800 3361.1200 1786.5600 ;
      RECT 1067.7600 1785.4800 3305.4200 1785.6400 ;
      RECT 1067.7600 1785.3800 3370.4200 1785.4800 ;
      RECT 2449.0800 1783.8400 3370.4200 1785.3800 ;
      RECT 0.0000 1783.8400 5.7000 1786.0400 ;
      RECT 1067.7600 1783.4400 1285.6400 1785.3800 ;
      RECT 167.4150 1783.4400 953.1450 1785.6400 ;
      RECT 5.3000 1783.4400 5.7000 1783.8400 ;
      RECT 2449.0800 1783.1800 3302.8200 1783.8400 ;
      RECT 1948.5000 1783.1800 2166.5200 1785.3800 ;
      RECT 157.4200 1783.1800 1285.6400 1783.4400 ;
      RECT 3368.7200 1782.7600 3370.4200 1783.8400 ;
      RECT 3305.0200 1782.7600 3365.1200 1783.8400 ;
      RECT 157.4200 1782.7600 3302.8200 1783.1800 ;
      RECT 5.3000 1782.7600 155.2200 1783.4400 ;
      RECT 0.0000 1782.7600 1.7000 1783.8400 ;
      RECT 157.4200 1782.5900 3370.4200 1782.7600 ;
      RECT 0.0000 1782.5900 155.2200 1782.7600 ;
      RECT 0.0000 1781.1200 3370.4200 1782.5900 ;
      RECT 0.0000 1780.0900 5.7000 1781.1200 ;
      RECT 3364.7200 1780.0400 3370.4200 1781.1200 ;
      RECT 3307.6200 1780.0400 3361.1200 1781.1200 ;
      RECT 154.8200 1780.0400 3305.4200 1781.1200 ;
      RECT 9.3000 1780.0400 152.6200 1781.1200 ;
      RECT 1.1000 1780.0400 5.7000 1780.0900 ;
      RECT 1.1000 1779.1900 3370.4200 1780.0400 ;
      RECT 0.0000 1778.4000 3370.4200 1779.1900 ;
      RECT 157.4200 1777.6300 3302.8200 1778.4000 ;
      RECT 1067.7600 1777.4700 3302.8200 1777.6300 ;
      RECT 3368.7200 1777.3200 3370.4200 1778.4000 ;
      RECT 3305.0200 1777.3200 3365.1200 1778.4000 ;
      RECT 2449.0800 1777.3200 3302.8200 1777.4700 ;
      RECT 157.4200 1777.3200 1002.6200 1777.6300 ;
      RECT 5.3000 1777.3200 155.2200 1778.4000 ;
      RECT 0.0000 1777.3200 1.7000 1778.4000 ;
      RECT 2449.0800 1775.6800 3370.4200 1777.3200 ;
      RECT 0.0000 1775.6800 1002.6200 1777.3200 ;
      RECT 1067.7600 1775.4300 1285.6400 1777.4700 ;
      RECT 1011.2200 1775.4300 1059.1600 1777.6300 ;
      RECT 154.8200 1775.4300 1002.6200 1775.6800 ;
      RECT 2449.0800 1775.2700 3305.4200 1775.6800 ;
      RECT 2392.5400 1775.2700 2440.4800 1777.4700 ;
      RECT 2172.3200 1775.2700 2380.3400 1777.4700 ;
      RECT 1948.5000 1775.2700 2166.5200 1777.4700 ;
      RECT 1731.8800 1775.2700 1939.9000 1777.4700 ;
      RECT 1511.6600 1775.2700 1719.6800 1777.4700 ;
      RECT 1291.4400 1775.2700 1499.4600 1777.4700 ;
      RECT 154.8200 1775.2700 1285.6400 1775.4300 ;
      RECT 154.8200 1775.2300 3305.4200 1775.2700 ;
      RECT 1065.1600 1774.8700 3305.4200 1775.2300 ;
      RECT 3364.7200 1774.6000 3370.4200 1775.6800 ;
      RECT 3307.6200 1774.6000 3361.1200 1775.6800 ;
      RECT 2446.4800 1774.6000 3305.4200 1774.8700 ;
      RECT 154.8200 1774.6000 1005.2200 1775.2300 ;
      RECT 9.3000 1774.6000 152.6200 1775.6800 ;
      RECT 0.0000 1774.6000 5.7000 1775.6800 ;
      RECT 1065.1600 1773.0300 1283.0400 1774.8700 ;
      RECT 1011.2200 1773.0300 1059.1600 1775.2300 ;
      RECT 0.0000 1773.0300 1005.2200 1774.6000 ;
      RECT 2446.4800 1772.9600 3370.4200 1774.6000 ;
      RECT 0.0000 1772.9600 1283.0400 1773.0300 ;
      RECT 2446.4800 1772.6700 3302.8200 1772.9600 ;
      RECT 2392.5400 1772.6700 2440.4800 1774.8700 ;
      RECT 2172.3200 1772.6700 2380.3400 1774.8700 ;
      RECT 1945.9000 1772.6700 2163.9200 1774.8700 ;
      RECT 1731.8800 1772.6700 1939.9000 1774.8700 ;
      RECT 1511.6600 1772.6700 1719.6800 1774.8700 ;
      RECT 1291.4400 1772.6700 1499.4600 1774.8700 ;
      RECT 157.4200 1772.6700 1283.0400 1772.9600 ;
      RECT 3368.7200 1771.8800 3370.4200 1772.9600 ;
      RECT 3305.0200 1771.8800 3365.1200 1772.9600 ;
      RECT 157.4200 1771.8800 3302.8200 1772.6700 ;
      RECT 5.3000 1771.8800 155.2200 1772.9600 ;
      RECT 0.0000 1771.8800 1.7000 1772.9600 ;
      RECT 0.0000 1770.2600 3370.4200 1771.8800 ;
      RECT 1015.0800 1770.2400 3370.4200 1770.2600 ;
      RECT 0.0000 1770.2400 1012.8800 1770.2600 ;
      RECT 1015.0800 1770.0000 3305.4200 1770.2400 ;
      RECT 0.0000 1769.7200 5.7000 1770.2400 ;
      RECT 1015.0800 1769.1800 1293.0000 1770.0000 ;
      RECT 154.8200 1769.1800 1012.8800 1770.2400 ;
      RECT 3364.7200 1769.1600 3370.4200 1770.2400 ;
      RECT 3307.6200 1769.1600 3361.1200 1770.2400 ;
      RECT 2396.3000 1769.1600 3305.4200 1770.0000 ;
      RECT 154.8200 1769.1600 1293.0000 1769.1800 ;
      RECT 9.3000 1769.1600 152.6200 1770.2400 ;
      RECT 1.1000 1769.1600 5.7000 1769.7200 ;
      RECT 2396.3000 1768.9200 3370.4200 1769.1600 ;
      RECT 2176.0800 1768.9200 2394.1000 1770.0000 ;
      RECT 1735.6400 1768.9200 2173.8800 1770.0000 ;
      RECT 1515.4200 1768.9200 1733.4400 1770.0000 ;
      RECT 1295.2000 1768.9200 1513.2200 1770.0000 ;
      RECT 1.1000 1768.9200 1293.0000 1769.1600 ;
      RECT 1.1000 1768.8200 3370.4200 1768.9200 ;
      RECT 0.0000 1767.5200 3370.4200 1768.8200 ;
      RECT 3368.7200 1766.4400 3370.4200 1767.5200 ;
      RECT 3305.0200 1766.4400 3365.1200 1767.5200 ;
      RECT 157.4200 1766.4400 3302.8200 1767.5200 ;
      RECT 5.3000 1766.4400 155.2200 1767.5200 ;
      RECT 0.0000 1766.4400 1.7000 1767.5200 ;
      RECT 0.0000 1764.8000 3370.4200 1766.4400 ;
      RECT 3364.7200 1763.7200 3370.4200 1764.8000 ;
      RECT 3307.6200 1763.7200 3361.1200 1764.8000 ;
      RECT 154.8200 1763.7200 3305.4200 1764.8000 ;
      RECT 9.3000 1763.7200 152.6200 1764.8000 ;
      RECT 0.0000 1763.7200 5.7000 1764.8000 ;
      RECT 0.0000 1762.0800 3370.4200 1763.7200 ;
      RECT 3368.7200 1761.0000 3370.4200 1762.0800 ;
      RECT 3305.0200 1761.0000 3365.1200 1762.0800 ;
      RECT 157.4200 1761.0000 3302.8200 1762.0800 ;
      RECT 5.3000 1761.0000 155.2200 1762.0800 ;
      RECT 0.0000 1761.0000 1.7000 1762.0800 ;
      RECT 0.0000 1759.3600 3370.4200 1761.0000 ;
      RECT 0.0000 1758.7400 5.7000 1759.3600 ;
      RECT 3364.7200 1758.2800 3370.4200 1759.3600 ;
      RECT 3307.6200 1758.2800 3361.1200 1759.3600 ;
      RECT 154.8200 1758.2800 3305.4200 1759.3600 ;
      RECT 9.3000 1758.2800 152.6200 1759.3600 ;
      RECT 1.1000 1758.2800 5.7000 1758.7400 ;
      RECT 1.1000 1757.8400 3370.4200 1758.2800 ;
      RECT 0.0000 1756.6400 3370.4200 1757.8400 ;
      RECT 3368.7200 1755.5600 3370.4200 1756.6400 ;
      RECT 3305.0200 1755.5600 3365.1200 1756.6400 ;
      RECT 157.4200 1755.5600 3302.8200 1756.6400 ;
      RECT 5.3000 1755.5600 155.2200 1756.6400 ;
      RECT 0.0000 1755.5600 1.7000 1756.6400 ;
      RECT 0.0000 1753.9200 3370.4200 1755.5600 ;
      RECT 3364.7200 1752.8400 3370.4200 1753.9200 ;
      RECT 3307.6200 1752.8400 3361.1200 1753.9200 ;
      RECT 154.8200 1752.8400 3305.4200 1753.9200 ;
      RECT 9.3000 1752.8400 152.6200 1753.9200 ;
      RECT 0.0000 1752.8400 5.7000 1753.9200 ;
      RECT 0.0000 1751.2000 3370.4200 1752.8400 ;
      RECT 3368.7200 1750.1200 3370.4200 1751.2000 ;
      RECT 3305.0200 1750.1200 3365.1200 1751.2000 ;
      RECT 157.4200 1750.1200 3302.8200 1751.2000 ;
      RECT 5.3000 1750.1200 155.2200 1751.2000 ;
      RECT 0.0000 1750.1200 1.7000 1751.2000 ;
      RECT 0.0000 1748.4800 3370.4200 1750.1200 ;
      RECT 0.0000 1747.7600 5.7000 1748.4800 ;
      RECT 3364.7200 1747.4000 3370.4200 1748.4800 ;
      RECT 3307.6200 1747.4000 3361.1200 1748.4800 ;
      RECT 154.8200 1747.4000 3305.4200 1748.4800 ;
      RECT 9.3000 1747.4000 152.6200 1748.4800 ;
      RECT 1.1000 1747.4000 5.7000 1747.7600 ;
      RECT 1.1000 1746.8600 3370.4200 1747.4000 ;
      RECT 0.0000 1745.7600 3370.4200 1746.8600 ;
      RECT 3368.7200 1744.6800 3370.4200 1745.7600 ;
      RECT 3305.0200 1744.6800 3365.1200 1745.7600 ;
      RECT 157.4200 1744.6800 3302.8200 1745.7600 ;
      RECT 5.3000 1744.6800 155.2200 1745.7600 ;
      RECT 0.0000 1744.6800 1.7000 1745.7600 ;
      RECT 0.0000 1743.0400 3370.4200 1744.6800 ;
      RECT 3364.7200 1741.9600 3370.4200 1743.0400 ;
      RECT 3307.6200 1741.9600 3361.1200 1743.0400 ;
      RECT 154.8200 1741.9600 3305.4200 1743.0400 ;
      RECT 9.3000 1741.9600 152.6200 1743.0400 ;
      RECT 0.0000 1741.9600 5.7000 1743.0400 ;
      RECT 0.0000 1740.3200 3370.4200 1741.9600 ;
      RECT 3368.7200 1739.2400 3370.4200 1740.3200 ;
      RECT 3305.0200 1739.2400 3365.1200 1740.3200 ;
      RECT 157.4200 1739.2400 3302.8200 1740.3200 ;
      RECT 5.3000 1739.2400 155.2200 1740.3200 ;
      RECT 0.0000 1739.2400 1.7000 1740.3200 ;
      RECT 0.0000 1737.6000 3370.4200 1739.2400 ;
      RECT 0.0000 1736.7800 5.7000 1737.6000 ;
      RECT 3364.7200 1736.5200 3370.4200 1737.6000 ;
      RECT 3307.6200 1736.5200 3361.1200 1737.6000 ;
      RECT 154.8200 1736.5200 3305.4200 1737.6000 ;
      RECT 9.3000 1736.5200 152.6200 1737.6000 ;
      RECT 1.1000 1736.5200 5.7000 1736.7800 ;
      RECT 1.1000 1735.8800 3370.4200 1736.5200 ;
      RECT 0.0000 1734.8800 3370.4200 1735.8800 ;
      RECT 3368.7200 1733.8000 3370.4200 1734.8800 ;
      RECT 3305.0200 1733.8000 3365.1200 1734.8800 ;
      RECT 157.4200 1733.8000 3302.8200 1734.8800 ;
      RECT 5.3000 1733.8000 155.2200 1734.8800 ;
      RECT 0.0000 1733.8000 1.7000 1734.8800 ;
      RECT 0.0000 1732.1600 3370.4200 1733.8000 ;
      RECT 3364.7200 1731.0800 3370.4200 1732.1600 ;
      RECT 3307.6200 1731.0800 3361.1200 1732.1600 ;
      RECT 154.8200 1731.0800 3305.4200 1732.1600 ;
      RECT 9.3000 1731.0800 152.6200 1732.1600 ;
      RECT 0.0000 1731.0800 5.7000 1732.1600 ;
      RECT 0.0000 1729.4400 3370.4200 1731.0800 ;
      RECT 3368.7200 1728.3600 3370.4200 1729.4400 ;
      RECT 3305.0200 1728.3600 3365.1200 1729.4400 ;
      RECT 157.4200 1728.3600 3302.8200 1729.4400 ;
      RECT 5.3000 1728.3600 155.2200 1729.4400 ;
      RECT 0.0000 1728.3600 1.7000 1729.4400 ;
      RECT 0.0000 1726.7200 3370.4200 1728.3600 ;
      RECT 0.0000 1725.8000 5.7000 1726.7200 ;
      RECT 3364.7200 1725.6400 3370.4200 1726.7200 ;
      RECT 3307.6200 1725.6400 3361.1200 1726.7200 ;
      RECT 154.8200 1725.6400 3305.4200 1726.7200 ;
      RECT 9.3000 1725.6400 152.6200 1726.7200 ;
      RECT 1.1000 1725.6400 5.7000 1725.8000 ;
      RECT 1.1000 1724.9000 3370.4200 1725.6400 ;
      RECT 0.0000 1724.0000 3370.4200 1724.9000 ;
      RECT 3368.7200 1722.9200 3370.4200 1724.0000 ;
      RECT 3305.0200 1722.9200 3365.1200 1724.0000 ;
      RECT 157.4200 1722.9200 3302.8200 1724.0000 ;
      RECT 5.3000 1722.9200 155.2200 1724.0000 ;
      RECT 0.0000 1722.9200 1.7000 1724.0000 ;
      RECT 0.0000 1721.2800 3370.4200 1722.9200 ;
      RECT 3364.7200 1720.2000 3370.4200 1721.2800 ;
      RECT 3307.6200 1720.2000 3361.1200 1721.2800 ;
      RECT 154.8200 1720.2000 3305.4200 1721.2800 ;
      RECT 9.3000 1720.2000 152.6200 1721.2800 ;
      RECT 0.0000 1720.2000 5.7000 1721.2800 ;
      RECT 0.0000 1718.5600 3370.4200 1720.2000 ;
      RECT 3368.7200 1717.4800 3370.4200 1718.5600 ;
      RECT 3305.0200 1717.4800 3365.1200 1718.5600 ;
      RECT 157.4200 1717.4800 3302.8200 1718.5600 ;
      RECT 5.3000 1717.4800 155.2200 1718.5600 ;
      RECT 0.0000 1717.4800 1.7000 1718.5600 ;
      RECT 0.0000 1715.8400 3370.4200 1717.4800 ;
      RECT 0.0000 1715.4300 5.7000 1715.8400 ;
      RECT 3364.7200 1714.7600 3370.4200 1715.8400 ;
      RECT 3307.6200 1714.7600 3361.1200 1715.8400 ;
      RECT 154.8200 1714.7600 3305.4200 1715.8400 ;
      RECT 9.3000 1714.7600 152.6200 1715.8400 ;
      RECT 1.1000 1714.7600 5.7000 1715.4300 ;
      RECT 1.1000 1714.5300 3370.4200 1714.7600 ;
      RECT 0.0000 1713.1200 3370.4200 1714.5300 ;
      RECT 3368.7200 1712.0400 3370.4200 1713.1200 ;
      RECT 3305.0200 1712.0400 3365.1200 1713.1200 ;
      RECT 157.4200 1712.0400 3302.8200 1713.1200 ;
      RECT 5.3000 1712.0400 155.2200 1713.1200 ;
      RECT 0.0000 1712.0400 1.7000 1713.1200 ;
      RECT 0.0000 1710.4000 3370.4200 1712.0400 ;
      RECT 3364.7200 1709.3200 3370.4200 1710.4000 ;
      RECT 3307.6200 1709.3200 3361.1200 1710.4000 ;
      RECT 154.8200 1709.3200 3305.4200 1710.4000 ;
      RECT 9.3000 1709.3200 152.6200 1710.4000 ;
      RECT 0.0000 1709.3200 5.7000 1710.4000 ;
      RECT 0.0000 1707.6800 3370.4200 1709.3200 ;
      RECT 3368.7200 1706.6000 3370.4200 1707.6800 ;
      RECT 3305.0200 1706.6000 3365.1200 1707.6800 ;
      RECT 157.4200 1706.6000 3302.8200 1707.6800 ;
      RECT 5.3000 1706.6000 155.2200 1707.6800 ;
      RECT 0.0000 1706.6000 1.7000 1707.6800 ;
      RECT 0.0000 1704.9600 3370.4200 1706.6000 ;
      RECT 0.0000 1704.4500 5.7000 1704.9600 ;
      RECT 3364.7200 1703.8800 3370.4200 1704.9600 ;
      RECT 3307.6200 1703.8800 3361.1200 1704.9600 ;
      RECT 154.8200 1703.8800 3305.4200 1704.9600 ;
      RECT 9.3000 1703.8800 152.6200 1704.9600 ;
      RECT 1.1000 1703.8800 5.7000 1704.4500 ;
      RECT 1.1000 1703.5500 3370.4200 1703.8800 ;
      RECT 0.0000 1702.2400 3370.4200 1703.5500 ;
      RECT 3368.7200 1701.1600 3370.4200 1702.2400 ;
      RECT 3305.0200 1701.1600 3365.1200 1702.2400 ;
      RECT 157.4200 1701.1600 3302.8200 1702.2400 ;
      RECT 5.3000 1701.1600 155.2200 1702.2400 ;
      RECT 0.0000 1701.1600 1.7000 1702.2400 ;
      RECT 0.0000 1699.5200 3370.4200 1701.1600 ;
      RECT 3364.7200 1698.4400 3370.4200 1699.5200 ;
      RECT 3307.6200 1698.4400 3361.1200 1699.5200 ;
      RECT 154.8200 1698.4400 3305.4200 1699.5200 ;
      RECT 9.3000 1698.4400 152.6200 1699.5200 ;
      RECT 0.0000 1698.4400 5.7000 1699.5200 ;
      RECT 0.0000 1696.8000 3370.4200 1698.4400 ;
      RECT 3368.7200 1695.7200 3370.4200 1696.8000 ;
      RECT 3305.0200 1695.7200 3365.1200 1696.8000 ;
      RECT 157.4200 1695.7200 3302.8200 1696.8000 ;
      RECT 5.3000 1695.7200 155.2200 1696.8000 ;
      RECT 0.0000 1695.7200 1.7000 1696.8000 ;
      RECT 0.0000 1694.0800 3370.4200 1695.7200 ;
      RECT 0.0000 1693.4700 5.7000 1694.0800 ;
      RECT 3364.7200 1693.0000 3370.4200 1694.0800 ;
      RECT 3307.6200 1693.0000 3361.1200 1694.0800 ;
      RECT 154.8200 1693.0000 3305.4200 1694.0800 ;
      RECT 9.3000 1693.0000 152.6200 1694.0800 ;
      RECT 1.1000 1693.0000 5.7000 1693.4700 ;
      RECT 1.1000 1692.5700 3370.4200 1693.0000 ;
      RECT 0.0000 1691.3600 3370.4200 1692.5700 ;
      RECT 3368.7200 1690.2800 3370.4200 1691.3600 ;
      RECT 3305.0200 1690.2800 3365.1200 1691.3600 ;
      RECT 157.4200 1690.2800 3302.8200 1691.3600 ;
      RECT 5.3000 1690.2800 155.2200 1691.3600 ;
      RECT 0.0000 1690.2800 1.7000 1691.3600 ;
      RECT 0.0000 1688.6400 3370.4200 1690.2800 ;
      RECT 3364.7200 1687.5600 3370.4200 1688.6400 ;
      RECT 3307.6200 1687.5600 3361.1200 1688.6400 ;
      RECT 154.8200 1687.5600 3305.4200 1688.6400 ;
      RECT 9.3000 1687.5600 152.6200 1688.6400 ;
      RECT 0.0000 1687.5600 5.7000 1688.6400 ;
      RECT 0.0000 1685.9200 3370.4200 1687.5600 ;
      RECT 3368.7200 1684.8400 3370.4200 1685.9200 ;
      RECT 3305.0200 1684.8400 3365.1200 1685.9200 ;
      RECT 157.4200 1684.8400 3302.8200 1685.9200 ;
      RECT 5.3000 1684.8400 155.2200 1685.9200 ;
      RECT 0.0000 1684.8400 1.7000 1685.9200 ;
      RECT 0.0000 1683.2000 3370.4200 1684.8400 ;
      RECT 0.0000 1682.4900 5.7000 1683.2000 ;
      RECT 3364.7200 1682.1200 3370.4200 1683.2000 ;
      RECT 3307.6200 1682.1200 3361.1200 1683.2000 ;
      RECT 154.8200 1682.1200 3305.4200 1683.2000 ;
      RECT 9.3000 1682.1200 152.6200 1683.2000 ;
      RECT 1.1000 1682.1200 5.7000 1682.4900 ;
      RECT 1.1000 1681.5900 3370.4200 1682.1200 ;
      RECT 0.0000 1680.4800 3370.4200 1681.5900 ;
      RECT 3368.7200 1679.4000 3370.4200 1680.4800 ;
      RECT 3305.0200 1679.4000 3365.1200 1680.4800 ;
      RECT 157.4200 1679.4000 3302.8200 1680.4800 ;
      RECT 5.3000 1679.4000 155.2200 1680.4800 ;
      RECT 0.0000 1679.4000 1.7000 1680.4800 ;
      RECT 0.0000 1677.7600 3370.4200 1679.4000 ;
      RECT 3364.7200 1676.6800 3370.4200 1677.7600 ;
      RECT 3307.6200 1676.6800 3361.1200 1677.7600 ;
      RECT 154.8200 1676.6800 3305.4200 1677.7600 ;
      RECT 9.3000 1676.6800 152.6200 1677.7600 ;
      RECT 0.0000 1676.6800 5.7000 1677.7600 ;
      RECT 0.0000 1675.0400 3370.4200 1676.6800 ;
      RECT 3368.7200 1673.9600 3370.4200 1675.0400 ;
      RECT 3305.0200 1673.9600 3365.1200 1675.0400 ;
      RECT 157.4200 1673.9600 3302.8200 1675.0400 ;
      RECT 5.3000 1673.9600 155.2200 1675.0400 ;
      RECT 0.0000 1673.9600 1.7000 1675.0400 ;
      RECT 0.0000 1672.3200 3370.4200 1673.9600 ;
      RECT 0.0000 1671.5100 5.7000 1672.3200 ;
      RECT 3364.7200 1671.2400 3370.4200 1672.3200 ;
      RECT 3307.6200 1671.2400 3361.1200 1672.3200 ;
      RECT 154.8200 1671.2400 3305.4200 1672.3200 ;
      RECT 9.3000 1671.2400 152.6200 1672.3200 ;
      RECT 1.1000 1671.2400 5.7000 1671.5100 ;
      RECT 1.1000 1670.6100 3370.4200 1671.2400 ;
      RECT 0.0000 1669.6000 3370.4200 1670.6100 ;
      RECT 3368.7200 1668.5200 3370.4200 1669.6000 ;
      RECT 3305.0200 1668.5200 3365.1200 1669.6000 ;
      RECT 157.4200 1668.5200 3302.8200 1669.6000 ;
      RECT 5.3000 1668.5200 155.2200 1669.6000 ;
      RECT 0.0000 1668.5200 1.7000 1669.6000 ;
      RECT 0.0000 1666.8800 3370.4200 1668.5200 ;
      RECT 3364.7200 1665.8000 3370.4200 1666.8800 ;
      RECT 3307.6200 1665.8000 3361.1200 1666.8800 ;
      RECT 154.8200 1665.8000 3305.4200 1666.8800 ;
      RECT 9.3000 1665.8000 152.6200 1666.8800 ;
      RECT 0.0000 1665.8000 5.7000 1666.8800 ;
      RECT 0.0000 1664.1600 3370.4200 1665.8000 ;
      RECT 3368.7200 1663.0800 3370.4200 1664.1600 ;
      RECT 3305.0200 1663.0800 3365.1200 1664.1600 ;
      RECT 157.4200 1663.0800 3302.8200 1664.1600 ;
      RECT 5.3000 1663.0800 155.2200 1664.1600 ;
      RECT 0.0000 1663.0800 1.7000 1664.1600 ;
      RECT 0.0000 1661.4400 3370.4200 1663.0800 ;
      RECT 0.0000 1661.1400 5.7000 1661.4400 ;
      RECT 3364.7200 1660.3600 3370.4200 1661.4400 ;
      RECT 3307.6200 1660.3600 3361.1200 1661.4400 ;
      RECT 154.8200 1660.3600 3305.4200 1661.4400 ;
      RECT 9.3000 1660.3600 152.6200 1661.4400 ;
      RECT 1.1000 1660.3600 5.7000 1661.1400 ;
      RECT 1.1000 1660.2400 3370.4200 1660.3600 ;
      RECT 0.0000 1658.7200 3370.4200 1660.2400 ;
      RECT 3368.7200 1657.6400 3370.4200 1658.7200 ;
      RECT 3305.0200 1657.6400 3365.1200 1658.7200 ;
      RECT 157.4200 1657.6400 3302.8200 1658.7200 ;
      RECT 5.3000 1657.6400 155.2200 1658.7200 ;
      RECT 0.0000 1657.6400 1.7000 1658.7200 ;
      RECT 0.0000 1656.0000 3370.4200 1657.6400 ;
      RECT 3364.7200 1654.9200 3370.4200 1656.0000 ;
      RECT 3307.6200 1654.9200 3361.1200 1656.0000 ;
      RECT 154.8200 1654.9200 3305.4200 1656.0000 ;
      RECT 9.3000 1654.9200 152.6200 1656.0000 ;
      RECT 0.0000 1654.9200 5.7000 1656.0000 ;
      RECT 0.0000 1653.2800 3370.4200 1654.9200 ;
      RECT 3368.7200 1652.2000 3370.4200 1653.2800 ;
      RECT 3305.0200 1652.2000 3365.1200 1653.2800 ;
      RECT 157.4200 1652.2000 3302.8200 1653.2800 ;
      RECT 5.3000 1652.2000 155.2200 1653.2800 ;
      RECT 0.0000 1652.2000 1.7000 1653.2800 ;
      RECT 0.0000 1650.5600 3370.4200 1652.2000 ;
      RECT 0.0000 1650.1600 5.7000 1650.5600 ;
      RECT 3364.7200 1649.4800 3370.4200 1650.5600 ;
      RECT 3307.6200 1649.4800 3361.1200 1650.5600 ;
      RECT 154.8200 1649.4800 3305.4200 1650.5600 ;
      RECT 9.3000 1649.4800 152.6200 1650.5600 ;
      RECT 1.1000 1649.4800 5.7000 1650.1600 ;
      RECT 1.1000 1649.2600 3370.4200 1649.4800 ;
      RECT 0.0000 1647.8400 3370.4200 1649.2600 ;
      RECT 3368.7200 1646.7600 3370.4200 1647.8400 ;
      RECT 3305.0200 1646.7600 3365.1200 1647.8400 ;
      RECT 157.4200 1646.7600 3302.8200 1647.8400 ;
      RECT 5.3000 1646.7600 155.2200 1647.8400 ;
      RECT 0.0000 1646.7600 1.7000 1647.8400 ;
      RECT 0.0000 1645.1200 3370.4200 1646.7600 ;
      RECT 3364.7200 1644.0400 3370.4200 1645.1200 ;
      RECT 3307.6200 1644.0400 3361.1200 1645.1200 ;
      RECT 154.8200 1644.0400 3305.4200 1645.1200 ;
      RECT 9.3000 1644.0400 152.6200 1645.1200 ;
      RECT 0.0000 1644.0400 5.7000 1645.1200 ;
      RECT 0.0000 1642.4000 3370.4200 1644.0400 ;
      RECT 3368.7200 1641.3200 3370.4200 1642.4000 ;
      RECT 3305.0200 1641.3200 3365.1200 1642.4000 ;
      RECT 157.4200 1641.3200 3302.8200 1642.4000 ;
      RECT 5.3000 1641.3200 155.2200 1642.4000 ;
      RECT 0.0000 1641.3200 1.7000 1642.4000 ;
      RECT 0.0000 1639.6800 3370.4200 1641.3200 ;
      RECT 0.0000 1639.1800 5.7000 1639.6800 ;
      RECT 3364.7200 1638.6000 3370.4200 1639.6800 ;
      RECT 3307.6200 1638.6000 3361.1200 1639.6800 ;
      RECT 154.8200 1638.6000 3305.4200 1639.6800 ;
      RECT 9.3000 1638.6000 152.6200 1639.6800 ;
      RECT 1.1000 1638.6000 5.7000 1639.1800 ;
      RECT 1.1000 1638.2800 3370.4200 1638.6000 ;
      RECT 0.0000 1636.9600 3370.4200 1638.2800 ;
      RECT 3368.7200 1635.8800 3370.4200 1636.9600 ;
      RECT 3305.0200 1635.8800 3365.1200 1636.9600 ;
      RECT 157.4200 1635.8800 3302.8200 1636.9600 ;
      RECT 5.3000 1635.8800 155.2200 1636.9600 ;
      RECT 0.0000 1635.8800 1.7000 1636.9600 ;
      RECT 0.0000 1634.2400 3370.4200 1635.8800 ;
      RECT 3364.7200 1633.1600 3370.4200 1634.2400 ;
      RECT 3307.6200 1633.1600 3361.1200 1634.2400 ;
      RECT 154.8200 1633.1600 3305.4200 1634.2400 ;
      RECT 9.3000 1633.1600 152.6200 1634.2400 ;
      RECT 0.0000 1633.1600 5.7000 1634.2400 ;
      RECT 0.0000 1631.5200 3370.4200 1633.1600 ;
      RECT 3368.7200 1630.4400 3370.4200 1631.5200 ;
      RECT 3305.0200 1630.4400 3365.1200 1631.5200 ;
      RECT 157.4200 1630.4400 3302.8200 1631.5200 ;
      RECT 5.3000 1630.4400 155.2200 1631.5200 ;
      RECT 0.0000 1630.4400 1.7000 1631.5200 ;
      RECT 0.0000 1628.8000 3370.4200 1630.4400 ;
      RECT 0.0000 1628.2000 5.7000 1628.8000 ;
      RECT 3364.7200 1627.7200 3370.4200 1628.8000 ;
      RECT 3307.6200 1627.7200 3361.1200 1628.8000 ;
      RECT 154.8200 1627.7200 3305.4200 1628.8000 ;
      RECT 9.3000 1627.7200 152.6200 1628.8000 ;
      RECT 1.1000 1627.7200 5.7000 1628.2000 ;
      RECT 1.1000 1627.3000 3370.4200 1627.7200 ;
      RECT 0.0000 1626.0800 3370.4200 1627.3000 ;
      RECT 3368.7200 1625.0000 3370.4200 1626.0800 ;
      RECT 3305.0200 1625.0000 3365.1200 1626.0800 ;
      RECT 157.4200 1625.0000 3302.8200 1626.0800 ;
      RECT 5.3000 1625.0000 155.2200 1626.0800 ;
      RECT 0.0000 1625.0000 1.7000 1626.0800 ;
      RECT 0.0000 1623.3600 3370.4200 1625.0000 ;
      RECT 3364.7200 1622.2800 3370.4200 1623.3600 ;
      RECT 3307.6200 1622.2800 3361.1200 1623.3600 ;
      RECT 154.8200 1622.2800 3305.4200 1623.3600 ;
      RECT 9.3000 1622.2800 152.6200 1623.3600 ;
      RECT 0.0000 1622.2800 5.7000 1623.3600 ;
      RECT 0.0000 1620.6400 3370.4200 1622.2800 ;
      RECT 3368.7200 1619.5600 3370.4200 1620.6400 ;
      RECT 3305.0200 1619.5600 3365.1200 1620.6400 ;
      RECT 157.4200 1619.5600 3302.8200 1620.6400 ;
      RECT 5.3000 1619.5600 155.2200 1620.6400 ;
      RECT 0.0000 1619.5600 1.7000 1620.6400 ;
      RECT 0.0000 1617.9200 3370.4200 1619.5600 ;
      RECT 0.0000 1617.2200 5.7000 1617.9200 ;
      RECT 3364.7200 1616.8400 3370.4200 1617.9200 ;
      RECT 3307.6200 1616.8400 3361.1200 1617.9200 ;
      RECT 154.8200 1616.8400 3305.4200 1617.9200 ;
      RECT 9.3000 1616.8400 152.6200 1617.9200 ;
      RECT 1.1000 1616.8400 5.7000 1617.2200 ;
      RECT 1.1000 1616.3200 3370.4200 1616.8400 ;
      RECT 0.0000 1615.2000 3370.4200 1616.3200 ;
      RECT 3368.7200 1614.1200 3370.4200 1615.2000 ;
      RECT 3305.0200 1614.1200 3365.1200 1615.2000 ;
      RECT 157.4200 1614.1200 3302.8200 1615.2000 ;
      RECT 5.3000 1614.1200 155.2200 1615.2000 ;
      RECT 0.0000 1614.1200 1.7000 1615.2000 ;
      RECT 0.0000 1612.4800 3370.4200 1614.1200 ;
      RECT 3364.7200 1611.4000 3370.4200 1612.4800 ;
      RECT 3307.6200 1611.4000 3361.1200 1612.4800 ;
      RECT 154.8200 1611.4000 3305.4200 1612.4800 ;
      RECT 9.3000 1611.4000 152.6200 1612.4800 ;
      RECT 0.0000 1611.4000 5.7000 1612.4800 ;
      RECT 0.0000 1609.7600 3370.4200 1611.4000 ;
      RECT 3368.7200 1608.6800 3370.4200 1609.7600 ;
      RECT 3305.0200 1608.6800 3365.1200 1609.7600 ;
      RECT 157.4200 1608.6800 3302.8200 1609.7600 ;
      RECT 5.3000 1608.6800 155.2200 1609.7600 ;
      RECT 0.0000 1608.6800 1.7000 1609.7600 ;
      RECT 0.0000 1607.0400 3370.4200 1608.6800 ;
      RECT 0.0000 1606.8500 5.7000 1607.0400 ;
      RECT 3364.7200 1605.9600 3370.4200 1607.0400 ;
      RECT 3307.6200 1605.9600 3361.1200 1607.0400 ;
      RECT 154.8200 1605.9600 3305.4200 1607.0400 ;
      RECT 9.3000 1605.9600 152.6200 1607.0400 ;
      RECT 1.1000 1605.9600 5.7000 1606.8500 ;
      RECT 1.1000 1605.9500 3370.4200 1605.9600 ;
      RECT 0.0000 1604.3200 3370.4200 1605.9500 ;
      RECT 3368.7200 1603.2400 3370.4200 1604.3200 ;
      RECT 3305.0200 1603.2400 3365.1200 1604.3200 ;
      RECT 157.4200 1603.2400 3302.8200 1604.3200 ;
      RECT 5.3000 1603.2400 155.2200 1604.3200 ;
      RECT 0.0000 1603.2400 1.7000 1604.3200 ;
      RECT 0.0000 1601.6000 3370.4200 1603.2400 ;
      RECT 3364.7200 1600.5200 3370.4200 1601.6000 ;
      RECT 3307.6200 1600.5200 3361.1200 1601.6000 ;
      RECT 154.8200 1600.5200 3305.4200 1601.6000 ;
      RECT 9.3000 1600.5200 152.6200 1601.6000 ;
      RECT 0.0000 1600.5200 5.7000 1601.6000 ;
      RECT 0.0000 1598.8800 3370.4200 1600.5200 ;
      RECT 3368.7200 1597.8000 3370.4200 1598.8800 ;
      RECT 3305.0200 1597.8000 3365.1200 1598.8800 ;
      RECT 157.4200 1597.8000 3302.8200 1598.8800 ;
      RECT 5.3000 1597.8000 155.2200 1598.8800 ;
      RECT 0.0000 1597.8000 1.7000 1598.8800 ;
      RECT 0.0000 1596.1600 3370.4200 1597.8000 ;
      RECT 0.0000 1595.8700 5.7000 1596.1600 ;
      RECT 3364.7200 1595.0800 3370.4200 1596.1600 ;
      RECT 3307.6200 1595.0800 3361.1200 1596.1600 ;
      RECT 154.8200 1595.0800 3305.4200 1596.1600 ;
      RECT 9.3000 1595.0800 152.6200 1596.1600 ;
      RECT 1.1000 1595.0800 5.7000 1595.8700 ;
      RECT 1.1000 1594.9700 3370.4200 1595.0800 ;
      RECT 0.0000 1593.4400 3370.4200 1594.9700 ;
      RECT 3368.7200 1592.3600 3370.4200 1593.4400 ;
      RECT 3305.0200 1592.3600 3365.1200 1593.4400 ;
      RECT 157.4200 1592.3600 3302.8200 1593.4400 ;
      RECT 5.3000 1592.3600 155.2200 1593.4400 ;
      RECT 0.0000 1592.3600 1.7000 1593.4400 ;
      RECT 0.0000 1590.7200 3370.4200 1592.3600 ;
      RECT 3364.7200 1589.6400 3370.4200 1590.7200 ;
      RECT 3307.6200 1589.6400 3361.1200 1590.7200 ;
      RECT 154.8200 1589.6400 3305.4200 1590.7200 ;
      RECT 9.3000 1589.6400 152.6200 1590.7200 ;
      RECT 0.0000 1589.6400 5.7000 1590.7200 ;
      RECT 0.0000 1588.0000 3370.4200 1589.6400 ;
      RECT 3368.7200 1586.9200 3370.4200 1588.0000 ;
      RECT 3305.0200 1586.9200 3365.1200 1588.0000 ;
      RECT 157.4200 1586.9200 3302.8200 1588.0000 ;
      RECT 5.3000 1586.9200 155.2200 1588.0000 ;
      RECT 0.0000 1586.9200 1.7000 1588.0000 ;
      RECT 0.0000 1585.2800 3370.4200 1586.9200 ;
      RECT 0.0000 1584.8900 5.7000 1585.2800 ;
      RECT 3364.7200 1584.2000 3370.4200 1585.2800 ;
      RECT 3307.6200 1584.2000 3361.1200 1585.2800 ;
      RECT 154.8200 1584.2000 3305.4200 1585.2800 ;
      RECT 9.3000 1584.2000 152.6200 1585.2800 ;
      RECT 1.1000 1584.2000 5.7000 1584.8900 ;
      RECT 1.1000 1583.9900 3370.4200 1584.2000 ;
      RECT 0.0000 1582.5600 3370.4200 1583.9900 ;
      RECT 3368.7200 1581.4800 3370.4200 1582.5600 ;
      RECT 3305.0200 1581.4800 3365.1200 1582.5600 ;
      RECT 157.4200 1581.4800 3302.8200 1582.5600 ;
      RECT 5.3000 1581.4800 155.2200 1582.5600 ;
      RECT 0.0000 1581.4800 1.7000 1582.5600 ;
      RECT 0.0000 1579.8400 3370.4200 1581.4800 ;
      RECT 3364.7200 1578.7600 3370.4200 1579.8400 ;
      RECT 3307.6200 1578.7600 3361.1200 1579.8400 ;
      RECT 154.8200 1578.7600 3305.4200 1579.8400 ;
      RECT 9.3000 1578.7600 152.6200 1579.8400 ;
      RECT 0.0000 1578.7600 5.7000 1579.8400 ;
      RECT 0.0000 1577.1200 3370.4200 1578.7600 ;
      RECT 3368.7200 1576.0400 3370.4200 1577.1200 ;
      RECT 3305.0200 1576.0400 3365.1200 1577.1200 ;
      RECT 157.4200 1576.0400 3302.8200 1577.1200 ;
      RECT 5.3000 1576.0400 155.2200 1577.1200 ;
      RECT 0.0000 1576.0400 1.7000 1577.1200 ;
      RECT 0.0000 1574.4000 3370.4200 1576.0400 ;
      RECT 0.0000 1573.9100 5.7000 1574.4000 ;
      RECT 3364.7200 1573.3200 3370.4200 1574.4000 ;
      RECT 3307.6200 1573.3200 3361.1200 1574.4000 ;
      RECT 154.8200 1573.3200 3305.4200 1574.4000 ;
      RECT 9.3000 1573.3200 152.6200 1574.4000 ;
      RECT 1.1000 1573.3200 5.7000 1573.9100 ;
      RECT 1.1000 1573.0100 3370.4200 1573.3200 ;
      RECT 0.0000 1571.7000 3370.4200 1573.0100 ;
      RECT 1077.7200 1571.6800 3370.4200 1571.7000 ;
      RECT 0.0000 1571.6800 1015.2800 1571.7000 ;
      RECT 1077.7200 1571.4400 3302.8200 1571.6800 ;
      RECT 1077.7200 1570.6200 1295.6000 1571.4400 ;
      RECT 1017.4800 1570.6200 1075.5200 1571.7000 ;
      RECT 157.4200 1570.6200 1015.2800 1571.6800 ;
      RECT 3368.7200 1570.6000 3370.4200 1571.6800 ;
      RECT 3305.0200 1570.6000 3365.1200 1571.6800 ;
      RECT 2436.3200 1570.6000 3302.8200 1571.4400 ;
      RECT 157.4200 1570.6000 1295.6000 1570.6200 ;
      RECT 5.3000 1570.6000 155.2200 1571.6800 ;
      RECT 0.0000 1570.6000 1.7000 1571.6800 ;
      RECT 2436.3200 1570.3600 3370.4200 1570.6000 ;
      RECT 2178.6800 1570.3600 2434.1200 1571.4400 ;
      RECT 1958.4600 1570.3600 2176.4800 1571.4400 ;
      RECT 1738.2400 1570.3600 1956.2600 1571.4400 ;
      RECT 1518.0200 1570.3600 1736.0400 1571.4400 ;
      RECT 1297.8000 1570.3600 1515.8200 1571.4400 ;
      RECT 0.0000 1570.3600 1295.6000 1570.6000 ;
      RECT 0.0000 1568.9600 3370.4200 1570.3600 ;
      RECT 154.8200 1568.6300 3305.4200 1568.9600 ;
      RECT 154.8200 1568.5300 1062.9600 1568.6300 ;
      RECT 1285.3800 1568.3700 3305.4200 1568.6300 ;
      RECT 3364.7200 1567.8800 3370.4200 1568.9600 ;
      RECT 3307.6200 1567.8800 3361.1200 1568.9600 ;
      RECT 2446.4800 1567.8800 3305.4200 1568.3700 ;
      RECT 154.8200 1567.8800 1005.2200 1568.5300 ;
      RECT 9.3000 1567.8800 152.6200 1568.9600 ;
      RECT 0.0000 1567.8800 5.7000 1568.9600 ;
      RECT 1071.3600 1566.4300 1279.3800 1568.6300 ;
      RECT 1065.1600 1566.3300 1283.0400 1566.4300 ;
      RECT 1011.2200 1566.3300 1059.1600 1568.5300 ;
      RECT 0.0000 1566.3300 1005.2200 1567.8800 ;
      RECT 2446.4800 1566.2400 3370.4200 1567.8800 ;
      RECT 0.0000 1566.2400 1283.0400 1566.3300 ;
      RECT 2446.4800 1566.1700 3302.8200 1566.2400 ;
      RECT 2392.5400 1566.1700 2440.4800 1568.3700 ;
      RECT 2172.3200 1566.1700 2380.3400 1568.3700 ;
      RECT 1952.1000 1566.1700 2160.1200 1568.3700 ;
      RECT 1731.8800 1566.1700 1939.9000 1568.3700 ;
      RECT 1511.6600 1566.1700 1719.6800 1568.3700 ;
      RECT 1291.4400 1566.1700 1499.4600 1568.3700 ;
      RECT 157.4200 1566.1700 1283.0400 1566.2400 ;
      RECT 157.4200 1566.1300 3302.8200 1566.1700 ;
      RECT 1067.7600 1566.0300 3302.8200 1566.1300 ;
      RECT 1287.9800 1565.7700 3302.8200 1566.0300 ;
      RECT 3368.7200 1565.1600 3370.4200 1566.2400 ;
      RECT 3305.0200 1565.1600 3365.1200 1566.2400 ;
      RECT 2449.0800 1565.1600 3302.8200 1565.7700 ;
      RECT 157.4200 1565.1600 1002.6200 1566.1300 ;
      RECT 5.3000 1565.1600 155.2200 1566.2400 ;
      RECT 0.0000 1565.1600 1.7000 1566.2400 ;
      RECT 1011.2200 1563.9300 1059.1600 1566.1300 ;
      RECT 0.0000 1563.9300 1002.6200 1565.1600 ;
      RECT 1071.3600 1563.8300 1279.3800 1566.0300 ;
      RECT 0.0000 1563.8300 1065.5600 1563.9300 ;
      RECT 2449.0800 1563.5700 3370.4200 1565.1600 ;
      RECT 2392.5400 1563.5700 2440.4800 1565.7700 ;
      RECT 2172.3200 1563.5700 2380.3400 1565.7700 ;
      RECT 1952.1000 1563.5700 2160.1200 1565.7700 ;
      RECT 1731.8800 1563.5700 1939.9000 1565.7700 ;
      RECT 1511.6600 1563.5700 1719.6800 1565.7700 ;
      RECT 1291.4400 1563.5700 1499.4600 1565.7700 ;
      RECT 0.0000 1563.5700 1285.6400 1563.8300 ;
      RECT 0.0000 1563.5200 3370.4200 1563.5700 ;
      RECT 0.0000 1562.9300 5.7000 1563.5200 ;
      RECT 3364.7200 1562.4400 3370.4200 1563.5200 ;
      RECT 3307.6200 1562.4400 3361.1200 1563.5200 ;
      RECT 154.8200 1562.4400 3305.4200 1563.5200 ;
      RECT 9.3000 1562.4400 152.6200 1563.5200 ;
      RECT 1.1000 1562.4400 5.7000 1562.9300 ;
      RECT 1.1000 1562.0300 3370.4200 1562.4400 ;
      RECT 0.0000 1560.8000 3370.4200 1562.0300 ;
      RECT 3368.7200 1559.7200 3370.4200 1560.8000 ;
      RECT 3305.0200 1559.7200 3365.1200 1560.8000 ;
      RECT 157.4200 1559.7200 3302.8200 1560.8000 ;
      RECT 5.3000 1559.7200 155.2200 1560.8000 ;
      RECT 0.0000 1559.7200 1.7000 1560.8000 ;
      RECT 0.0000 1559.6100 3370.4200 1559.7200 ;
      RECT 154.8200 1558.6000 3370.4200 1559.6100 ;
      RECT 9.3000 1558.6000 151.9400 1559.6100 ;
      RECT 0.0000 1558.6000 5.7000 1559.6100 ;
      RECT 1285.3800 1558.3400 3370.4200 1558.6000 ;
      RECT 2446.4800 1558.0800 3370.4200 1558.3400 ;
      RECT 3364.7200 1557.0000 3370.4200 1558.0800 ;
      RECT 3307.6200 1557.0000 3361.1200 1558.0800 ;
      RECT 2446.4800 1557.0000 3305.4200 1558.0800 ;
      RECT 167.4150 1556.4000 953.1450 1558.6000 ;
      RECT 0.0000 1556.4000 1.7000 1558.6000 ;
      RECT 2446.4800 1556.1400 3370.4200 1557.0000 ;
      RECT 0.0000 1556.1400 1283.0400 1556.4000 ;
      RECT 0.0000 1556.1000 3370.4200 1556.1400 ;
      RECT 1065.0600 1556.0000 3370.4200 1556.1000 ;
      RECT 0.0000 1556.0000 1062.6600 1556.1000 ;
      RECT 1287.9800 1555.8400 3370.4200 1556.0000 ;
      RECT 1945.8000 1555.7400 3370.4200 1555.8400 ;
      RECT 1287.9800 1555.7400 1943.4000 1555.8400 ;
      RECT 2449.0800 1555.3600 3370.4200 1555.7400 ;
      RECT 0.0000 1555.3600 5.7000 1556.0000 ;
      RECT 3368.7200 1554.2800 3370.4200 1555.3600 ;
      RECT 3305.0200 1554.2800 3365.1200 1555.3600 ;
      RECT 2449.0800 1554.2800 3302.8200 1555.3600 ;
      RECT 5.3000 1554.2800 5.7000 1555.3600 ;
      RECT 0.0000 1554.2800 1.7000 1555.3600 ;
      RECT 167.4150 1553.8000 953.1450 1556.0000 ;
      RECT 0.0000 1553.8000 5.7000 1554.2800 ;
      RECT 2449.0800 1553.5400 3370.4200 1554.2800 ;
      RECT 1065.0600 1553.5400 1285.6400 1553.8000 ;
      RECT 157.4200 1552.7900 1062.6600 1553.8000 ;
      RECT 0.0000 1552.7900 155.2200 1553.8000 ;
      RECT 1945.8000 1552.6400 3370.4200 1553.5400 ;
      RECT 0.0000 1552.6400 1062.6600 1552.7900 ;
      RECT 0.0000 1552.5600 5.7000 1552.6400 ;
      RECT 1065.0600 1552.1000 1943.4000 1553.5400 ;
      RECT 154.8200 1552.1000 1062.6600 1552.6400 ;
      RECT 1945.8000 1551.8400 3305.4200 1552.6400 ;
      RECT 154.8200 1551.8400 1943.4000 1552.1000 ;
      RECT 1.1000 1551.6600 5.7000 1552.5600 ;
      RECT 3364.7200 1551.5600 3370.4200 1552.6400 ;
      RECT 3307.6200 1551.5600 3361.1200 1552.6400 ;
      RECT 154.8200 1551.5600 3305.4200 1551.8400 ;
      RECT 9.3000 1551.5600 152.6200 1552.6400 ;
      RECT 0.0000 1551.5600 5.7000 1551.6600 ;
      RECT 0.0000 1549.9200 3370.4200 1551.5600 ;
      RECT 157.4200 1549.1400 3302.8200 1549.9200 ;
      RECT 1287.9800 1548.8800 3302.8200 1549.1400 ;
      RECT 3368.7200 1548.8400 3370.4200 1549.9200 ;
      RECT 3305.0200 1548.8400 3365.1200 1549.9200 ;
      RECT 2168.7200 1548.8400 3302.8200 1548.8800 ;
      RECT 157.4200 1548.8400 1065.5600 1549.1400 ;
      RECT 5.3000 1548.8400 155.2200 1549.9200 ;
      RECT 0.0000 1548.8400 1.7000 1549.9200 ;
      RECT 0.0000 1547.9900 1065.5600 1548.8400 ;
      RECT 2168.7200 1547.8300 3370.4200 1548.8400 ;
      RECT 1287.9800 1547.8300 1946.3000 1548.8800 ;
      RECT 2449.0800 1547.2000 3370.4200 1547.8300 ;
      RECT 0.0000 1547.2000 1002.6200 1547.9900 ;
      RECT 1071.3600 1546.9400 1279.3800 1549.1400 ;
      RECT 1062.4600 1546.9400 1065.5600 1547.9900 ;
      RECT 1952.1000 1546.6800 2160.1200 1548.8800 ;
      RECT 1943.2000 1546.6800 1946.3000 1547.8300 ;
      RECT 1062.4600 1546.5400 1285.6400 1546.9400 ;
      RECT 1943.2000 1546.2800 2166.5200 1546.6800 ;
      RECT 3364.7200 1546.1200 3370.4200 1547.2000 ;
      RECT 3307.6200 1546.1200 3361.1200 1547.2000 ;
      RECT 2449.0800 1546.1200 3305.4200 1547.2000 ;
      RECT 154.8200 1546.1200 1002.6200 1547.2000 ;
      RECT 9.3000 1546.1200 152.6200 1547.2000 ;
      RECT 0.0000 1546.1200 5.7000 1547.2000 ;
      RECT 1062.4600 1545.7900 1062.9600 1546.5400 ;
      RECT 1011.2200 1545.7900 1059.1600 1547.9900 ;
      RECT 0.0000 1545.7900 1002.6200 1546.1200 ;
      RECT 2449.0800 1545.6300 3370.4200 1546.1200 ;
      RECT 2392.5400 1545.6300 2440.4800 1547.8300 ;
      RECT 2172.3200 1545.6300 2380.3400 1547.8300 ;
      RECT 2166.1200 1545.6300 2166.5200 1546.2800 ;
      RECT 1943.2000 1545.6300 1943.7000 1546.2800 ;
      RECT 1731.8800 1545.6300 1939.9000 1547.8300 ;
      RECT 1511.6600 1545.6300 1719.6800 1547.8300 ;
      RECT 1291.4400 1545.6300 1499.4600 1547.8300 ;
      RECT 1285.3800 1545.6300 1285.6400 1546.5400 ;
      RECT 0.0000 1545.5900 1062.9600 1545.7900 ;
      RECT 2166.1200 1545.2300 3370.4200 1545.6300 ;
      RECT 1285.3800 1545.2300 1943.7000 1545.6300 ;
      RECT 2446.4800 1544.4800 3370.4200 1545.2300 ;
      RECT 0.0000 1544.4800 1005.2200 1545.5900 ;
      RECT 1071.3600 1544.3400 1279.3800 1546.5400 ;
      RECT 1952.1000 1544.0800 2160.1200 1546.2800 ;
      RECT 3368.7200 1543.4000 3370.4200 1544.4800 ;
      RECT 3305.0200 1543.4000 3365.1200 1544.4800 ;
      RECT 2446.4800 1543.4000 3302.8200 1544.4800 ;
      RECT 157.4200 1543.4000 1005.2200 1544.4800 ;
      RECT 5.3000 1543.4000 155.2200 1544.4800 ;
      RECT 0.0000 1543.4000 1.7000 1544.4800 ;
      RECT 1065.1600 1543.3900 1283.0400 1544.3400 ;
      RECT 1011.2200 1543.3900 1059.1600 1545.5900 ;
      RECT 0.0000 1543.3900 1005.2200 1543.4000 ;
      RECT 2446.4800 1543.0300 3370.4200 1543.4000 ;
      RECT 2392.5400 1543.0300 2440.4800 1545.2300 ;
      RECT 2172.3200 1543.0300 2380.3400 1545.2300 ;
      RECT 1945.9000 1543.0300 2163.9200 1544.0800 ;
      RECT 1731.8800 1543.0300 1939.9000 1545.2300 ;
      RECT 1511.6600 1543.0300 1719.6800 1545.2300 ;
      RECT 1291.4400 1543.0300 1499.4600 1545.2300 ;
      RECT 0.0000 1543.0300 1283.0400 1543.3900 ;
      RECT 0.0000 1541.7600 3370.4200 1543.0300 ;
      RECT 0.0000 1541.5800 5.7000 1541.7600 ;
      RECT 3364.7200 1540.6800 3370.4200 1541.7600 ;
      RECT 3307.6200 1540.6800 3361.1200 1541.7600 ;
      RECT 154.8200 1540.6800 3305.4200 1541.7600 ;
      RECT 9.3000 1540.6800 152.6200 1541.7600 ;
      RECT 1.1000 1540.6800 5.7000 1541.5800 ;
      RECT 0.0000 1540.6200 3370.4200 1540.6800 ;
      RECT 1057.5000 1540.3600 3370.4200 1540.6200 ;
      RECT 1057.5000 1539.5400 1293.0000 1540.3600 ;
      RECT 0.0000 1539.5400 1055.3000 1540.6200 ;
      RECT 0.0000 1539.4600 1293.0000 1539.5400 ;
      RECT 2396.3000 1539.2800 3370.4200 1540.3600 ;
      RECT 2176.0800 1539.2800 2394.1000 1540.3600 ;
      RECT 1735.6400 1539.2800 2173.8800 1540.3600 ;
      RECT 1515.4200 1539.2800 1733.4400 1540.3600 ;
      RECT 1295.2000 1539.2800 1513.2200 1540.3600 ;
      RECT 1075.1200 1539.2800 1293.0000 1539.4600 ;
      RECT 1075.1200 1539.2000 3370.4200 1539.2800 ;
      RECT 1955.8600 1539.0400 3370.4200 1539.2000 ;
      RECT 0.0000 1539.0400 1072.9200 1539.4600 ;
      RECT 1075.1200 1538.3800 1953.6600 1539.2000 ;
      RECT 157.4200 1538.3800 1072.9200 1539.0400 ;
      RECT 1955.8600 1538.1200 3302.8200 1539.0400 ;
      RECT 157.4200 1538.1200 1953.6600 1538.3800 ;
      RECT 3368.7200 1537.9600 3370.4200 1539.0400 ;
      RECT 3305.0200 1537.9600 3365.1200 1539.0400 ;
      RECT 157.4200 1537.9600 3302.8200 1538.1200 ;
      RECT 5.3000 1537.9600 155.2200 1539.0400 ;
      RECT 0.0000 1537.9600 1.7000 1539.0400 ;
      RECT 0.0000 1536.3200 3370.4200 1537.9600 ;
      RECT 3364.7200 1535.2400 3370.4200 1536.3200 ;
      RECT 3307.6200 1535.2400 3361.1200 1536.3200 ;
      RECT 154.8200 1535.2400 3305.4200 1536.3200 ;
      RECT 9.3000 1535.2400 152.6200 1536.3200 ;
      RECT 0.0000 1535.2400 5.7000 1536.3200 ;
      RECT 0.0000 1533.6000 3370.4200 1535.2400 ;
      RECT 3368.7200 1532.5200 3370.4200 1533.6000 ;
      RECT 3305.0200 1532.5200 3365.1200 1533.6000 ;
      RECT 157.4200 1532.5200 3302.8200 1533.6000 ;
      RECT 5.3000 1532.5200 155.2200 1533.6000 ;
      RECT 0.0000 1532.5200 1.7000 1533.6000 ;
      RECT 0.0000 1530.8800 3370.4200 1532.5200 ;
      RECT 0.0000 1530.6000 5.7000 1530.8800 ;
      RECT 3364.7200 1529.8000 3370.4200 1530.8800 ;
      RECT 3307.6200 1529.8000 3361.1200 1530.8800 ;
      RECT 154.8200 1529.8000 3305.4200 1530.8800 ;
      RECT 9.3000 1529.8000 152.6200 1530.8800 ;
      RECT 1.1000 1529.8000 5.7000 1530.6000 ;
      RECT 1.1000 1529.7000 3370.4200 1529.8000 ;
      RECT 0.0000 1528.1600 3370.4200 1529.7000 ;
      RECT 3368.7200 1527.0800 3370.4200 1528.1600 ;
      RECT 3305.0200 1527.0800 3365.1200 1528.1600 ;
      RECT 157.4200 1527.0800 3302.8200 1528.1600 ;
      RECT 5.3000 1527.0800 155.2200 1528.1600 ;
      RECT 0.0000 1527.0800 1.7000 1528.1600 ;
      RECT 0.0000 1525.4400 3370.4200 1527.0800 ;
      RECT 3364.7200 1524.3600 3370.4200 1525.4400 ;
      RECT 3307.6200 1524.3600 3361.1200 1525.4400 ;
      RECT 154.8200 1524.3600 3305.4200 1525.4400 ;
      RECT 9.3000 1524.3600 152.6200 1525.4400 ;
      RECT 0.0000 1524.3600 5.7000 1525.4400 ;
      RECT 0.0000 1522.7200 3370.4200 1524.3600 ;
      RECT 3368.7200 1521.6400 3370.4200 1522.7200 ;
      RECT 3305.0200 1521.6400 3365.1200 1522.7200 ;
      RECT 157.4200 1521.6400 3302.8200 1522.7200 ;
      RECT 5.3000 1521.6400 155.2200 1522.7200 ;
      RECT 0.0000 1521.6400 1.7000 1522.7200 ;
      RECT 0.0000 1520.0000 3370.4200 1521.6400 ;
      RECT 0.0000 1519.6200 5.7000 1520.0000 ;
      RECT 3364.7200 1518.9200 3370.4200 1520.0000 ;
      RECT 3307.6200 1518.9200 3361.1200 1520.0000 ;
      RECT 154.8200 1518.9200 3305.4200 1520.0000 ;
      RECT 9.3000 1518.9200 152.6200 1520.0000 ;
      RECT 1.1000 1518.9200 5.7000 1519.6200 ;
      RECT 1.1000 1518.7200 3370.4200 1518.9200 ;
      RECT 0.0000 1517.2800 3370.4200 1518.7200 ;
      RECT 3368.7200 1516.2000 3370.4200 1517.2800 ;
      RECT 3305.0200 1516.2000 3365.1200 1517.2800 ;
      RECT 157.4200 1516.2000 3302.8200 1517.2800 ;
      RECT 5.3000 1516.2000 155.2200 1517.2800 ;
      RECT 0.0000 1516.2000 1.7000 1517.2800 ;
      RECT 0.0000 1514.5600 3370.4200 1516.2000 ;
      RECT 3364.7200 1513.4800 3370.4200 1514.5600 ;
      RECT 3307.6200 1513.4800 3361.1200 1514.5600 ;
      RECT 154.8200 1513.4800 3305.4200 1514.5600 ;
      RECT 9.3000 1513.4800 152.6200 1514.5600 ;
      RECT 0.0000 1513.4800 5.7000 1514.5600 ;
      RECT 0.0000 1511.8400 3370.4200 1513.4800 ;
      RECT 3368.7200 1510.7600 3370.4200 1511.8400 ;
      RECT 3305.0200 1510.7600 3365.1200 1511.8400 ;
      RECT 157.4200 1510.7600 3302.8200 1511.8400 ;
      RECT 5.3000 1510.7600 155.2200 1511.8400 ;
      RECT 0.0000 1510.7600 1.7000 1511.8400 ;
      RECT 0.0000 1509.1200 3370.4200 1510.7600 ;
      RECT 0.0000 1508.6400 5.7000 1509.1200 ;
      RECT 3364.7200 1508.0400 3370.4200 1509.1200 ;
      RECT 3307.6200 1508.0400 3361.1200 1509.1200 ;
      RECT 154.8200 1508.0400 3305.4200 1509.1200 ;
      RECT 9.3000 1508.0400 152.6200 1509.1200 ;
      RECT 1.1000 1508.0400 5.7000 1508.6400 ;
      RECT 1.1000 1507.7400 3370.4200 1508.0400 ;
      RECT 0.0000 1506.4000 3370.4200 1507.7400 ;
      RECT 3368.7200 1505.3200 3370.4200 1506.4000 ;
      RECT 3305.0200 1505.3200 3365.1200 1506.4000 ;
      RECT 157.4200 1505.3200 3302.8200 1506.4000 ;
      RECT 5.3000 1505.3200 155.2200 1506.4000 ;
      RECT 0.0000 1505.3200 1.7000 1506.4000 ;
      RECT 0.0000 1503.6800 3370.4200 1505.3200 ;
      RECT 3364.7200 1502.6000 3370.4200 1503.6800 ;
      RECT 3307.6200 1502.6000 3361.1200 1503.6800 ;
      RECT 154.8200 1502.6000 3305.4200 1503.6800 ;
      RECT 9.3000 1502.6000 152.6200 1503.6800 ;
      RECT 0.0000 1502.6000 5.7000 1503.6800 ;
      RECT 0.0000 1500.9600 3370.4200 1502.6000 ;
      RECT 3368.7200 1499.8800 3370.4200 1500.9600 ;
      RECT 3305.0200 1499.8800 3365.1200 1500.9600 ;
      RECT 157.4200 1499.8800 3302.8200 1500.9600 ;
      RECT 5.3000 1499.8800 155.2200 1500.9600 ;
      RECT 0.0000 1499.8800 1.7000 1500.9600 ;
      RECT 0.0000 1498.2700 3370.4200 1499.8800 ;
      RECT 1.1000 1498.2400 3370.4200 1498.2700 ;
      RECT 1.1000 1497.3700 5.7000 1498.2400 ;
      RECT 3364.7200 1497.1600 3370.4200 1498.2400 ;
      RECT 3307.6200 1497.1600 3361.1200 1498.2400 ;
      RECT 154.8200 1497.1600 3305.4200 1498.2400 ;
      RECT 9.3000 1497.1600 152.6200 1498.2400 ;
      RECT 0.0000 1497.1600 5.7000 1497.3700 ;
      RECT 0.0000 1495.5200 3370.4200 1497.1600 ;
      RECT 3368.7200 1494.4400 3370.4200 1495.5200 ;
      RECT 3305.0200 1494.4400 3365.1200 1495.5200 ;
      RECT 157.4200 1494.4400 3302.8200 1495.5200 ;
      RECT 5.3000 1494.4400 155.2200 1495.5200 ;
      RECT 0.0000 1494.4400 1.7000 1495.5200 ;
      RECT 0.0000 1492.8000 3370.4200 1494.4400 ;
      RECT 3364.7200 1491.7200 3370.4200 1492.8000 ;
      RECT 3307.6200 1491.7200 3361.1200 1492.8000 ;
      RECT 154.8200 1491.7200 3305.4200 1492.8000 ;
      RECT 9.3000 1491.7200 152.6200 1492.8000 ;
      RECT 0.0000 1491.7200 5.7000 1492.8000 ;
      RECT 0.0000 1490.0800 3370.4200 1491.7200 ;
      RECT 3368.7200 1489.0000 3370.4200 1490.0800 ;
      RECT 3305.0200 1489.0000 3365.1200 1490.0800 ;
      RECT 157.4200 1489.0000 3302.8200 1490.0800 ;
      RECT 5.3000 1489.0000 155.2200 1490.0800 ;
      RECT 0.0000 1489.0000 1.7000 1490.0800 ;
      RECT 0.0000 1487.3600 3370.4200 1489.0000 ;
      RECT 0.0000 1487.2900 5.7000 1487.3600 ;
      RECT 1.1000 1486.3900 5.7000 1487.2900 ;
      RECT 3364.7200 1486.2800 3370.4200 1487.3600 ;
      RECT 3307.6200 1486.2800 3361.1200 1487.3600 ;
      RECT 154.8200 1486.2800 3305.4200 1487.3600 ;
      RECT 9.3000 1486.2800 152.6200 1487.3600 ;
      RECT 0.0000 1486.2800 5.7000 1486.3900 ;
      RECT 0.0000 1484.6400 3370.4200 1486.2800 ;
      RECT 3368.7200 1483.5600 3370.4200 1484.6400 ;
      RECT 3305.0200 1483.5600 3365.1200 1484.6400 ;
      RECT 157.4200 1483.5600 3302.8200 1484.6400 ;
      RECT 5.3000 1483.5600 155.2200 1484.6400 ;
      RECT 0.0000 1483.5600 1.7000 1484.6400 ;
      RECT 0.0000 1481.9200 3370.4200 1483.5600 ;
      RECT 3364.7200 1480.8400 3370.4200 1481.9200 ;
      RECT 3307.6200 1480.8400 3361.1200 1481.9200 ;
      RECT 154.8200 1480.8400 3305.4200 1481.9200 ;
      RECT 9.3000 1480.8400 152.6200 1481.9200 ;
      RECT 0.0000 1480.8400 5.7000 1481.9200 ;
      RECT 0.0000 1479.2000 3370.4200 1480.8400 ;
      RECT 3368.7200 1478.1200 3370.4200 1479.2000 ;
      RECT 3305.0200 1478.1200 3365.1200 1479.2000 ;
      RECT 157.4200 1478.1200 3302.8200 1479.2000 ;
      RECT 5.3000 1478.1200 155.2200 1479.2000 ;
      RECT 0.0000 1478.1200 1.7000 1479.2000 ;
      RECT 0.0000 1476.4800 3370.4200 1478.1200 ;
      RECT 0.0000 1476.3100 5.7000 1476.4800 ;
      RECT 1.1000 1475.4100 5.7000 1476.3100 ;
      RECT 3364.7200 1475.4000 3370.4200 1476.4800 ;
      RECT 3307.6200 1475.4000 3361.1200 1476.4800 ;
      RECT 154.8200 1475.4000 3305.4200 1476.4800 ;
      RECT 9.3000 1475.4000 152.6200 1476.4800 ;
      RECT 0.0000 1475.4000 5.7000 1475.4100 ;
      RECT 0.0000 1473.7600 3370.4200 1475.4000 ;
      RECT 3368.7200 1472.6800 3370.4200 1473.7600 ;
      RECT 3305.0200 1472.6800 3365.1200 1473.7600 ;
      RECT 157.4200 1472.6800 3302.8200 1473.7600 ;
      RECT 5.3000 1472.6800 155.2200 1473.7600 ;
      RECT 0.0000 1472.6800 1.7000 1473.7600 ;
      RECT 0.0000 1471.0400 3370.4200 1472.6800 ;
      RECT 3364.7200 1469.9600 3370.4200 1471.0400 ;
      RECT 3307.6200 1469.9600 3361.1200 1471.0400 ;
      RECT 154.8200 1469.9600 3305.4200 1471.0400 ;
      RECT 9.3000 1469.9600 152.6200 1471.0400 ;
      RECT 0.0000 1469.9600 5.7000 1471.0400 ;
      RECT 0.0000 1468.3200 3370.4200 1469.9600 ;
      RECT 3368.7200 1467.2400 3370.4200 1468.3200 ;
      RECT 3305.0200 1467.2400 3365.1200 1468.3200 ;
      RECT 157.4200 1467.2400 3302.8200 1468.3200 ;
      RECT 5.3000 1467.2400 155.2200 1468.3200 ;
      RECT 0.0000 1467.2400 1.7000 1468.3200 ;
      RECT 0.0000 1465.6000 3370.4200 1467.2400 ;
      RECT 0.0000 1465.3300 5.7000 1465.6000 ;
      RECT 3364.7200 1464.5200 3370.4200 1465.6000 ;
      RECT 3307.6200 1464.5200 3361.1200 1465.6000 ;
      RECT 154.8200 1464.5200 3305.4200 1465.6000 ;
      RECT 9.3000 1464.5200 152.6200 1465.6000 ;
      RECT 1.1000 1464.5200 5.7000 1465.3300 ;
      RECT 1.1000 1464.4300 3370.4200 1464.5200 ;
      RECT 0.0000 1462.8800 3370.4200 1464.4300 ;
      RECT 3368.7200 1461.8000 3370.4200 1462.8800 ;
      RECT 3305.0200 1461.8000 3365.1200 1462.8800 ;
      RECT 157.4200 1461.8000 3302.8200 1462.8800 ;
      RECT 5.3000 1461.8000 155.2200 1462.8800 ;
      RECT 0.0000 1461.8000 1.7000 1462.8800 ;
      RECT 0.0000 1460.1600 3370.4200 1461.8000 ;
      RECT 3364.7200 1459.0800 3370.4200 1460.1600 ;
      RECT 3307.6200 1459.0800 3361.1200 1460.1600 ;
      RECT 154.8200 1459.0800 3305.4200 1460.1600 ;
      RECT 9.3000 1459.0800 152.6200 1460.1600 ;
      RECT 0.0000 1459.0800 5.7000 1460.1600 ;
      RECT 0.0000 1457.4400 3370.4200 1459.0800 ;
      RECT 3368.7200 1456.3600 3370.4200 1457.4400 ;
      RECT 3305.0200 1456.3600 3365.1200 1457.4400 ;
      RECT 157.4200 1456.3600 3302.8200 1457.4400 ;
      RECT 5.3000 1456.3600 155.2200 1457.4400 ;
      RECT 0.0000 1456.3600 1.7000 1457.4400 ;
      RECT 0.0000 1454.7200 3370.4200 1456.3600 ;
      RECT 0.0000 1454.3500 5.7000 1454.7200 ;
      RECT 3364.7200 1453.6400 3370.4200 1454.7200 ;
      RECT 3307.6200 1453.6400 3361.1200 1454.7200 ;
      RECT 154.8200 1453.6400 3305.4200 1454.7200 ;
      RECT 9.3000 1453.6400 152.6200 1454.7200 ;
      RECT 1.1000 1453.6400 5.7000 1454.3500 ;
      RECT 1.1000 1453.4500 3370.4200 1453.6400 ;
      RECT 0.0000 1452.0000 3370.4200 1453.4500 ;
      RECT 3368.7200 1450.9200 3370.4200 1452.0000 ;
      RECT 3305.0200 1450.9200 3365.1200 1452.0000 ;
      RECT 157.4200 1450.9200 3302.8200 1452.0000 ;
      RECT 5.3000 1450.9200 155.2200 1452.0000 ;
      RECT 0.0000 1450.9200 1.7000 1452.0000 ;
      RECT 0.0000 1449.2800 3370.4200 1450.9200 ;
      RECT 3364.7200 1448.2000 3370.4200 1449.2800 ;
      RECT 3307.6200 1448.2000 3361.1200 1449.2800 ;
      RECT 154.8200 1448.2000 3305.4200 1449.2800 ;
      RECT 9.3000 1448.2000 152.6200 1449.2800 ;
      RECT 0.0000 1448.2000 5.7000 1449.2800 ;
      RECT 0.0000 1446.5600 3370.4200 1448.2000 ;
      RECT 3368.7200 1445.4800 3370.4200 1446.5600 ;
      RECT 3305.0200 1445.4800 3365.1200 1446.5600 ;
      RECT 157.4200 1445.4800 3302.8200 1446.5600 ;
      RECT 5.3000 1445.4800 155.2200 1446.5600 ;
      RECT 0.0000 1445.4800 1.7000 1446.5600 ;
      RECT 0.0000 1443.9800 3370.4200 1445.4800 ;
      RECT 1.1000 1443.8400 3370.4200 1443.9800 ;
      RECT 1.1000 1443.0800 5.7000 1443.8400 ;
      RECT 3364.7200 1442.7600 3370.4200 1443.8400 ;
      RECT 3307.6200 1442.7600 3361.1200 1443.8400 ;
      RECT 154.8200 1442.7600 3305.4200 1443.8400 ;
      RECT 9.3000 1442.7600 152.6200 1443.8400 ;
      RECT 0.0000 1442.7600 5.7000 1443.0800 ;
      RECT 0.0000 1441.1200 3370.4200 1442.7600 ;
      RECT 3368.7200 1440.0400 3370.4200 1441.1200 ;
      RECT 3305.0200 1440.0400 3365.1200 1441.1200 ;
      RECT 157.4200 1440.0400 3302.8200 1441.1200 ;
      RECT 5.3000 1440.0400 155.2200 1441.1200 ;
      RECT 0.0000 1440.0400 1.7000 1441.1200 ;
      RECT 0.0000 1438.4000 3370.4200 1440.0400 ;
      RECT 3364.7200 1437.3200 3370.4200 1438.4000 ;
      RECT 3307.6200 1437.3200 3361.1200 1438.4000 ;
      RECT 154.8200 1437.3200 3305.4200 1438.4000 ;
      RECT 9.3000 1437.3200 152.6200 1438.4000 ;
      RECT 0.0000 1437.3200 5.7000 1438.4000 ;
      RECT 0.0000 1435.6800 3370.4200 1437.3200 ;
      RECT 3368.7200 1434.6000 3370.4200 1435.6800 ;
      RECT 3305.0200 1434.6000 3365.1200 1435.6800 ;
      RECT 157.4200 1434.6000 3302.8200 1435.6800 ;
      RECT 5.3000 1434.6000 155.2200 1435.6800 ;
      RECT 0.0000 1434.6000 1.7000 1435.6800 ;
      RECT 0.0000 1433.0000 3370.4200 1434.6000 ;
      RECT 1.1000 1432.9600 3370.4200 1433.0000 ;
      RECT 1.1000 1432.1000 5.7000 1432.9600 ;
      RECT 3364.7200 1431.8800 3370.4200 1432.9600 ;
      RECT 3307.6200 1431.8800 3361.1200 1432.9600 ;
      RECT 154.8200 1431.8800 3305.4200 1432.9600 ;
      RECT 9.3000 1431.8800 152.6200 1432.9600 ;
      RECT 0.0000 1431.8800 5.7000 1432.1000 ;
      RECT 0.0000 1430.2400 3370.4200 1431.8800 ;
      RECT 3368.7200 1429.1600 3370.4200 1430.2400 ;
      RECT 3305.0200 1429.1600 3365.1200 1430.2400 ;
      RECT 157.4200 1429.1600 3302.8200 1430.2400 ;
      RECT 5.3000 1429.1600 155.2200 1430.2400 ;
      RECT 0.0000 1429.1600 1.7000 1430.2400 ;
      RECT 0.0000 1427.5200 3370.4200 1429.1600 ;
      RECT 3364.7200 1426.4400 3370.4200 1427.5200 ;
      RECT 3307.6200 1426.4400 3361.1200 1427.5200 ;
      RECT 154.8200 1426.4400 3305.4200 1427.5200 ;
      RECT 9.3000 1426.4400 152.6200 1427.5200 ;
      RECT 0.0000 1426.4400 5.7000 1427.5200 ;
      RECT 0.0000 1424.8000 3370.4200 1426.4400 ;
      RECT 3368.7200 1423.7200 3370.4200 1424.8000 ;
      RECT 3305.0200 1423.7200 3365.1200 1424.8000 ;
      RECT 157.4200 1423.7200 3302.8200 1424.8000 ;
      RECT 5.3000 1423.7200 155.2200 1424.8000 ;
      RECT 0.0000 1423.7200 1.7000 1424.8000 ;
      RECT 0.0000 1422.0800 3370.4200 1423.7200 ;
      RECT 0.0000 1422.0200 5.7000 1422.0800 ;
      RECT 1.1000 1421.1200 5.7000 1422.0200 ;
      RECT 3364.7200 1421.0000 3370.4200 1422.0800 ;
      RECT 3307.6200 1421.0000 3361.1200 1422.0800 ;
      RECT 154.8200 1421.0000 3305.4200 1422.0800 ;
      RECT 9.3000 1421.0000 152.6200 1422.0800 ;
      RECT 0.0000 1421.0000 5.7000 1421.1200 ;
      RECT 0.0000 1419.3600 3370.4200 1421.0000 ;
      RECT 3368.7200 1418.2800 3370.4200 1419.3600 ;
      RECT 3305.0200 1418.2800 3365.1200 1419.3600 ;
      RECT 157.4200 1418.2800 3302.8200 1419.3600 ;
      RECT 5.3000 1418.2800 155.2200 1419.3600 ;
      RECT 0.0000 1418.2800 1.7000 1419.3600 ;
      RECT 0.0000 1416.6400 3370.4200 1418.2800 ;
      RECT 3364.7200 1415.5600 3370.4200 1416.6400 ;
      RECT 3307.6200 1415.5600 3361.1200 1416.6400 ;
      RECT 154.8200 1415.5600 3305.4200 1416.6400 ;
      RECT 9.3000 1415.5600 152.6200 1416.6400 ;
      RECT 0.0000 1415.5600 5.7000 1416.6400 ;
      RECT 0.0000 1413.9200 3370.4200 1415.5600 ;
      RECT 3368.7200 1412.8400 3370.4200 1413.9200 ;
      RECT 3305.0200 1412.8400 3365.1200 1413.9200 ;
      RECT 157.4200 1412.8400 3302.8200 1413.9200 ;
      RECT 5.3000 1412.8400 155.2200 1413.9200 ;
      RECT 0.0000 1412.8400 1.7000 1413.9200 ;
      RECT 0.0000 1411.2000 3370.4200 1412.8400 ;
      RECT 0.0000 1411.0400 5.7000 1411.2000 ;
      RECT 1.1000 1410.1400 5.7000 1411.0400 ;
      RECT 3364.7200 1410.1200 3370.4200 1411.2000 ;
      RECT 3307.6200 1410.1200 3361.1200 1411.2000 ;
      RECT 154.8200 1410.1200 3305.4200 1411.2000 ;
      RECT 9.3000 1410.1200 152.6200 1411.2000 ;
      RECT 0.0000 1410.1200 5.7000 1410.1400 ;
      RECT 0.0000 1408.4800 3370.4200 1410.1200 ;
      RECT 3368.7200 1407.4000 3370.4200 1408.4800 ;
      RECT 3305.0200 1407.4000 3365.1200 1408.4800 ;
      RECT 157.4200 1407.4000 3302.8200 1408.4800 ;
      RECT 5.3000 1407.4000 155.2200 1408.4800 ;
      RECT 0.0000 1407.4000 1.7000 1408.4800 ;
      RECT 0.0000 1405.7600 3370.4200 1407.4000 ;
      RECT 3364.7200 1404.6800 3370.4200 1405.7600 ;
      RECT 3307.6200 1404.6800 3361.1200 1405.7600 ;
      RECT 154.8200 1404.6800 3305.4200 1405.7600 ;
      RECT 9.3000 1404.6800 152.6200 1405.7600 ;
      RECT 0.0000 1404.6800 5.7000 1405.7600 ;
      RECT 0.0000 1403.0400 3370.4200 1404.6800 ;
      RECT 3368.7200 1401.9600 3370.4200 1403.0400 ;
      RECT 3305.0200 1401.9600 3365.1200 1403.0400 ;
      RECT 157.4200 1401.9600 3302.8200 1403.0400 ;
      RECT 5.3000 1401.9600 155.2200 1403.0400 ;
      RECT 0.0000 1401.9600 1.7000 1403.0400 ;
      RECT 0.0000 1400.3200 3370.4200 1401.9600 ;
      RECT 0.0000 1400.0600 5.7000 1400.3200 ;
      RECT 3364.7200 1399.2400 3370.4200 1400.3200 ;
      RECT 3307.6200 1399.2400 3361.1200 1400.3200 ;
      RECT 154.8200 1399.2400 3305.4200 1400.3200 ;
      RECT 9.3000 1399.2400 152.6200 1400.3200 ;
      RECT 1.1000 1399.2400 5.7000 1400.0600 ;
      RECT 1.1000 1399.1600 3370.4200 1399.2400 ;
      RECT 0.0000 1397.6000 3370.4200 1399.1600 ;
      RECT 3368.7200 1396.5200 3370.4200 1397.6000 ;
      RECT 3305.0200 1396.5200 3365.1200 1397.6000 ;
      RECT 157.4200 1396.5200 3302.8200 1397.6000 ;
      RECT 5.3000 1396.5200 155.2200 1397.6000 ;
      RECT 0.0000 1396.5200 1.7000 1397.6000 ;
      RECT 0.0000 1394.8800 3370.4200 1396.5200 ;
      RECT 3364.7200 1393.8000 3370.4200 1394.8800 ;
      RECT 3307.6200 1393.8000 3361.1200 1394.8800 ;
      RECT 154.8200 1393.8000 3305.4200 1394.8800 ;
      RECT 9.3000 1393.8000 152.6200 1394.8800 ;
      RECT 0.0000 1393.8000 5.7000 1394.8800 ;
      RECT 0.0000 1392.1600 3370.4200 1393.8000 ;
      RECT 3368.7200 1391.0800 3370.4200 1392.1600 ;
      RECT 3305.0200 1391.0800 3365.1200 1392.1600 ;
      RECT 157.4200 1391.0800 3302.8200 1392.1600 ;
      RECT 5.3000 1391.0800 155.2200 1392.1600 ;
      RECT 0.0000 1391.0800 1.7000 1392.1600 ;
      RECT 0.0000 1389.6900 3370.4200 1391.0800 ;
      RECT 1.1000 1389.4400 3370.4200 1389.6900 ;
      RECT 1.1000 1388.7900 5.7000 1389.4400 ;
      RECT 3364.7200 1388.3600 3370.4200 1389.4400 ;
      RECT 3307.6200 1388.3600 3361.1200 1389.4400 ;
      RECT 154.8200 1388.3600 3305.4200 1389.4400 ;
      RECT 9.3000 1388.3600 152.6200 1389.4400 ;
      RECT 0.0000 1388.3600 5.7000 1388.7900 ;
      RECT 0.0000 1386.7200 3370.4200 1388.3600 ;
      RECT 3368.7200 1385.6400 3370.4200 1386.7200 ;
      RECT 3305.0200 1385.6400 3365.1200 1386.7200 ;
      RECT 157.4200 1385.6400 3302.8200 1386.7200 ;
      RECT 5.3000 1385.6400 155.2200 1386.7200 ;
      RECT 0.0000 1385.6400 1.7000 1386.7200 ;
      RECT 0.0000 1384.0000 3370.4200 1385.6400 ;
      RECT 3364.7200 1382.9200 3370.4200 1384.0000 ;
      RECT 3307.6200 1382.9200 3361.1200 1384.0000 ;
      RECT 154.8200 1382.9200 3305.4200 1384.0000 ;
      RECT 9.3000 1382.9200 152.6200 1384.0000 ;
      RECT 0.0000 1382.9200 5.7000 1384.0000 ;
      RECT 0.0000 1381.2800 3370.4200 1382.9200 ;
      RECT 3368.7200 1380.2000 3370.4200 1381.2800 ;
      RECT 3305.0200 1380.2000 3365.1200 1381.2800 ;
      RECT 157.4200 1380.2000 3302.8200 1381.2800 ;
      RECT 5.3000 1380.2000 155.2200 1381.2800 ;
      RECT 0.0000 1380.2000 1.7000 1381.2800 ;
      RECT 0.0000 1378.7100 3370.4200 1380.2000 ;
      RECT 1.1000 1378.5600 3370.4200 1378.7100 ;
      RECT 1.1000 1377.8100 5.7000 1378.5600 ;
      RECT 3364.7200 1377.4800 3370.4200 1378.5600 ;
      RECT 3307.6200 1377.4800 3361.1200 1378.5600 ;
      RECT 154.8200 1377.4800 3305.4200 1378.5600 ;
      RECT 9.3000 1377.4800 152.6200 1378.5600 ;
      RECT 0.0000 1377.4800 5.7000 1377.8100 ;
      RECT 0.0000 1375.8400 3370.4200 1377.4800 ;
      RECT 3368.7200 1374.7600 3370.4200 1375.8400 ;
      RECT 3305.0200 1374.7600 3365.1200 1375.8400 ;
      RECT 157.4200 1374.7600 3302.8200 1375.8400 ;
      RECT 5.3000 1374.7600 155.2200 1375.8400 ;
      RECT 0.0000 1374.7600 1.7000 1375.8400 ;
      RECT 0.0000 1373.1200 3370.4200 1374.7600 ;
      RECT 3364.7200 1372.0400 3370.4200 1373.1200 ;
      RECT 3307.6200 1372.0400 3361.1200 1373.1200 ;
      RECT 154.8200 1372.0400 3305.4200 1373.1200 ;
      RECT 9.3000 1372.0400 152.6200 1373.1200 ;
      RECT 0.0000 1372.0400 5.7000 1373.1200 ;
      RECT 0.0000 1370.4000 3370.4200 1372.0400 ;
      RECT 3368.7200 1369.3200 3370.4200 1370.4000 ;
      RECT 3305.0200 1369.3200 3365.1200 1370.4000 ;
      RECT 157.4200 1369.3200 3302.8200 1370.4000 ;
      RECT 5.3000 1369.3200 155.2200 1370.4000 ;
      RECT 0.0000 1369.3200 1.7000 1370.4000 ;
      RECT 0.0000 1367.7300 3370.4200 1369.3200 ;
      RECT 1.1000 1367.6800 3370.4200 1367.7300 ;
      RECT 1.1000 1366.8300 5.7000 1367.6800 ;
      RECT 3364.7200 1366.6000 3370.4200 1367.6800 ;
      RECT 3307.6200 1366.6000 3361.1200 1367.6800 ;
      RECT 154.8200 1366.6000 3305.4200 1367.6800 ;
      RECT 9.3000 1366.6000 152.6200 1367.6800 ;
      RECT 0.0000 1366.6000 5.7000 1366.8300 ;
      RECT 0.0000 1364.9600 3370.4200 1366.6000 ;
      RECT 3368.7200 1363.8800 3370.4200 1364.9600 ;
      RECT 3305.0200 1363.8800 3365.1200 1364.9600 ;
      RECT 157.4200 1363.8800 3302.8200 1364.9600 ;
      RECT 5.3000 1363.8800 155.2200 1364.9600 ;
      RECT 0.0000 1363.8800 1.7000 1364.9600 ;
      RECT 0.0000 1362.2400 3370.4200 1363.8800 ;
      RECT 3364.7200 1361.1600 3370.4200 1362.2400 ;
      RECT 3307.6200 1361.1600 3361.1200 1362.2400 ;
      RECT 154.8200 1361.1600 3305.4200 1362.2400 ;
      RECT 9.3000 1361.1600 152.6200 1362.2400 ;
      RECT 0.0000 1361.1600 5.7000 1362.2400 ;
      RECT 0.0000 1359.5200 3370.4200 1361.1600 ;
      RECT 3368.7200 1358.4400 3370.4200 1359.5200 ;
      RECT 3305.0200 1358.4400 3365.1200 1359.5200 ;
      RECT 157.4200 1358.4400 3302.8200 1359.5200 ;
      RECT 5.3000 1358.4400 155.2200 1359.5200 ;
      RECT 0.0000 1358.4400 1.7000 1359.5200 ;
      RECT 0.0000 1356.8000 3370.4200 1358.4400 ;
      RECT 0.0000 1356.7500 5.7000 1356.8000 ;
      RECT 1.1000 1355.8500 5.7000 1356.7500 ;
      RECT 3364.7200 1355.7200 3370.4200 1356.8000 ;
      RECT 3307.6200 1355.7200 3361.1200 1356.8000 ;
      RECT 154.8200 1355.7200 3305.4200 1356.8000 ;
      RECT 9.3000 1355.7200 152.6200 1356.8000 ;
      RECT 0.0000 1355.7200 5.7000 1355.8500 ;
      RECT 0.0000 1354.0800 3370.4200 1355.7200 ;
      RECT 3368.7200 1353.0000 3370.4200 1354.0800 ;
      RECT 3305.0200 1353.0000 3365.1200 1354.0800 ;
      RECT 157.4200 1353.0000 3302.8200 1354.0800 ;
      RECT 5.3000 1353.0000 155.2200 1354.0800 ;
      RECT 0.0000 1353.0000 1.7000 1354.0800 ;
      RECT 0.0000 1351.3600 3370.4200 1353.0000 ;
      RECT 3364.7200 1350.2800 3370.4200 1351.3600 ;
      RECT 3307.6200 1350.2800 3361.1200 1351.3600 ;
      RECT 154.8200 1350.2800 3305.4200 1351.3600 ;
      RECT 9.3000 1350.2800 152.6200 1351.3600 ;
      RECT 0.0000 1350.2800 5.7000 1351.3600 ;
      RECT 0.0000 1348.6400 3370.4200 1350.2800 ;
      RECT 3368.7200 1347.5600 3370.4200 1348.6400 ;
      RECT 3305.0200 1347.5600 3365.1200 1348.6400 ;
      RECT 157.4200 1347.5600 3302.8200 1348.6400 ;
      RECT 5.3000 1347.5600 155.2200 1348.6400 ;
      RECT 0.0000 1347.5600 1.7000 1348.6400 ;
      RECT 0.0000 1345.9200 3370.4200 1347.5600 ;
      RECT 0.0000 1345.7700 5.7000 1345.9200 ;
      RECT 1.1000 1344.8700 5.7000 1345.7700 ;
      RECT 3364.7200 1344.8400 3370.4200 1345.9200 ;
      RECT 3307.6200 1344.8400 3361.1200 1345.9200 ;
      RECT 154.8200 1344.8400 3305.4200 1345.9200 ;
      RECT 9.3000 1344.8400 152.6200 1345.9200 ;
      RECT 0.0000 1344.8400 5.7000 1344.8700 ;
      RECT 0.0000 1343.2000 3370.4200 1344.8400 ;
      RECT 3368.7200 1342.1200 3370.4200 1343.2000 ;
      RECT 3305.0200 1342.1200 3365.1200 1343.2000 ;
      RECT 157.4200 1342.1200 3302.8200 1343.2000 ;
      RECT 5.3000 1342.1200 155.2200 1343.2000 ;
      RECT 0.0000 1342.1200 1.7000 1343.2000 ;
      RECT 0.0000 1342.0600 3370.4200 1342.1200 ;
      RECT 1017.4800 1341.8000 3370.4200 1342.0600 ;
      RECT 1017.4800 1340.9800 1295.6000 1341.8000 ;
      RECT 0.0000 1340.9800 1015.2800 1342.0600 ;
      RECT 2436.3200 1340.7200 3370.4200 1341.8000 ;
      RECT 2178.6800 1340.7200 2434.1200 1341.8000 ;
      RECT 1738.2400 1340.7200 2176.4800 1341.8000 ;
      RECT 1518.0200 1340.7200 1736.0400 1341.8000 ;
      RECT 1297.8000 1340.7200 1515.8200 1341.8000 ;
      RECT 0.0000 1340.7200 1295.6000 1340.9800 ;
      RECT 0.0000 1340.4800 3370.4200 1340.7200 ;
      RECT 3364.7200 1339.4000 3370.4200 1340.4800 ;
      RECT 3307.6200 1339.4000 3361.1200 1340.4800 ;
      RECT 154.8200 1339.4000 3305.4200 1340.4800 ;
      RECT 9.3000 1339.4000 152.6200 1340.4800 ;
      RECT 0.0000 1339.4000 5.7000 1340.4800 ;
      RECT 0.0000 1338.8900 3370.4200 1339.4000 ;
      RECT 1065.1600 1338.7300 3370.4200 1338.8900 ;
      RECT 2446.4800 1337.7600 3370.4200 1338.7300 ;
      RECT 0.0000 1337.7600 1005.2200 1338.8900 ;
      RECT 1065.1600 1336.6900 1283.0400 1338.7300 ;
      RECT 1011.2200 1336.6900 1059.1600 1338.8900 ;
      RECT 157.4200 1336.6900 1005.2200 1337.7600 ;
      RECT 3368.7200 1336.6800 3370.4200 1337.7600 ;
      RECT 3305.0200 1336.6800 3365.1200 1337.7600 ;
      RECT 2446.4800 1336.6800 3302.8200 1337.7600 ;
      RECT 157.4200 1336.6800 1283.0400 1336.6900 ;
      RECT 5.3000 1336.6800 155.2200 1337.7600 ;
      RECT 0.0000 1336.6800 1.7000 1337.7600 ;
      RECT 2446.4800 1336.5300 3370.4200 1336.6800 ;
      RECT 2392.5400 1336.5300 2440.4800 1338.7300 ;
      RECT 2172.3200 1336.5300 2380.3400 1338.7300 ;
      RECT 1945.9000 1336.5300 2163.9200 1338.7300 ;
      RECT 1731.8800 1336.5300 1939.9000 1338.7300 ;
      RECT 1511.6600 1336.5300 1719.6800 1338.7300 ;
      RECT 1291.4400 1336.5300 1499.4600 1338.7300 ;
      RECT 0.0000 1336.5300 1283.0400 1336.6800 ;
      RECT 0.0000 1336.4900 3370.4200 1336.5300 ;
      RECT 1067.7600 1336.1300 3370.4200 1336.4900 ;
      RECT 0.0000 1335.4000 1002.6200 1336.4900 ;
      RECT 2449.0800 1335.0400 3370.4200 1336.1300 ;
      RECT 1.1000 1335.0400 1002.6200 1335.4000 ;
      RECT 1.1000 1334.5000 5.7000 1335.0400 ;
      RECT 1067.7600 1334.2900 1285.6400 1336.1300 ;
      RECT 1011.2200 1334.2900 1059.1600 1336.4900 ;
      RECT 154.8200 1334.2900 1002.6200 1335.0400 ;
      RECT 3364.7200 1333.9600 3370.4200 1335.0400 ;
      RECT 3307.6200 1333.9600 3361.1200 1335.0400 ;
      RECT 2449.0800 1333.9600 3305.4200 1335.0400 ;
      RECT 154.8200 1333.9600 1285.6400 1334.2900 ;
      RECT 9.3000 1333.9600 152.6200 1335.0400 ;
      RECT 0.0000 1333.9600 5.7000 1334.5000 ;
      RECT 2449.0800 1333.9300 3370.4200 1333.9600 ;
      RECT 2392.5400 1333.9300 2440.4800 1336.1300 ;
      RECT 2172.3200 1333.9300 2380.3400 1336.1300 ;
      RECT 1948.5000 1333.9300 2166.5200 1336.1300 ;
      RECT 1731.8800 1333.9300 1939.9000 1336.1300 ;
      RECT 1511.6600 1333.9300 1719.6800 1336.1300 ;
      RECT 1291.4400 1333.9300 1499.4600 1336.1300 ;
      RECT 0.0000 1333.9300 1285.6400 1333.9600 ;
      RECT 0.0000 1332.3200 3370.4200 1333.9300 ;
      RECT 3368.7200 1331.2400 3370.4200 1332.3200 ;
      RECT 3305.0200 1331.2400 3365.1200 1332.3200 ;
      RECT 157.4200 1331.2400 3302.8200 1332.3200 ;
      RECT 5.3000 1331.2400 155.2200 1332.3200 ;
      RECT 0.0000 1331.2400 1.7000 1332.3200 ;
      RECT 0.0000 1329.7700 3370.4200 1331.2400 ;
      RECT 154.8200 1329.6000 3370.4200 1329.7700 ;
      RECT 154.8200 1328.9600 3305.4200 1329.6000 ;
      RECT 9.3000 1328.9600 152.6200 1329.7700 ;
      RECT 0.0000 1328.9600 5.7000 1329.7700 ;
      RECT 1065.1600 1328.7000 3305.4200 1328.9600 ;
      RECT 3364.7200 1328.5200 3370.4200 1329.6000 ;
      RECT 3307.6200 1328.5200 3361.1200 1329.6000 ;
      RECT 2446.4800 1328.5200 3305.4200 1328.7000 ;
      RECT 2446.4800 1326.8800 3370.4200 1328.5200 ;
      RECT 1065.1600 1326.7600 1283.0400 1328.7000 ;
      RECT 167.4150 1326.7600 953.1450 1328.9600 ;
      RECT 2446.4800 1326.5000 3302.8200 1326.8800 ;
      RECT 1945.9000 1326.5000 2163.9200 1328.7000 ;
      RECT 157.4200 1326.5000 1283.0400 1326.7600 ;
      RECT 157.4200 1326.3600 3302.8200 1326.5000 ;
      RECT 5.3000 1326.3600 155.2200 1326.7600 ;
      RECT 1067.7600 1326.1000 3302.8200 1326.3600 ;
      RECT 3368.7200 1325.8000 3370.4200 1326.8800 ;
      RECT 3305.0200 1325.8000 3365.1200 1326.8800 ;
      RECT 2449.0800 1325.8000 3302.8200 1326.1000 ;
      RECT 5.3000 1325.8000 5.7000 1326.3600 ;
      RECT 0.0000 1325.8000 1.7000 1328.9600 ;
      RECT 0.0000 1324.4200 5.7000 1325.8000 ;
      RECT 2449.0800 1324.1600 3370.4200 1325.8000 ;
      RECT 1067.7600 1324.1600 1285.6400 1326.1000 ;
      RECT 167.4150 1324.1600 953.1450 1326.3600 ;
      RECT 2449.0800 1323.9000 3305.4200 1324.1600 ;
      RECT 1948.5000 1323.9000 2166.5200 1326.1000 ;
      RECT 154.8200 1323.9000 1285.6400 1324.1600 ;
      RECT 1.1000 1323.5200 5.7000 1324.4200 ;
      RECT 3364.7200 1323.0800 3370.4200 1324.1600 ;
      RECT 3307.6200 1323.0800 3361.1200 1324.1600 ;
      RECT 154.8200 1323.0800 3305.4200 1323.9000 ;
      RECT 9.3000 1323.0800 152.6200 1324.1600 ;
      RECT 0.0000 1323.0800 5.7000 1323.5200 ;
      RECT 0.0000 1321.4400 3370.4200 1323.0800 ;
      RECT 3368.7200 1320.3600 3370.4200 1321.4400 ;
      RECT 3305.0200 1320.3600 3365.1200 1321.4400 ;
      RECT 157.4200 1320.3600 3302.8200 1321.4400 ;
      RECT 5.3000 1320.3600 155.2200 1321.4400 ;
      RECT 0.0000 1320.3600 1.7000 1321.4400 ;
      RECT 0.0000 1318.7200 3370.4200 1320.3600 ;
      RECT 154.8200 1318.3500 3305.4200 1318.7200 ;
      RECT 1067.7600 1318.1900 3305.4200 1318.3500 ;
      RECT 3364.7200 1317.6400 3370.4200 1318.7200 ;
      RECT 3307.6200 1317.6400 3361.1200 1318.7200 ;
      RECT 2449.0800 1317.6400 3305.4200 1318.1900 ;
      RECT 154.8200 1317.6400 1002.6200 1318.3500 ;
      RECT 9.3000 1317.6400 152.6200 1318.7200 ;
      RECT 0.0000 1317.6400 5.7000 1318.7200 ;
      RECT 1067.7600 1316.1500 1285.6400 1318.1900 ;
      RECT 1011.2200 1316.1500 1059.1600 1318.3500 ;
      RECT 0.0000 1316.1500 1002.6200 1317.6400 ;
      RECT 2449.0800 1316.0000 3370.4200 1317.6400 ;
      RECT 0.0000 1316.0000 1285.6400 1316.1500 ;
      RECT 2449.0800 1315.9900 3302.8200 1316.0000 ;
      RECT 2392.5400 1315.9900 2440.4800 1318.1900 ;
      RECT 2172.3200 1315.9900 2380.3400 1318.1900 ;
      RECT 1948.5000 1315.9900 2166.5200 1318.1900 ;
      RECT 1731.8800 1315.9900 1939.9000 1318.1900 ;
      RECT 1511.6600 1315.9900 1719.6800 1318.1900 ;
      RECT 1291.4400 1315.9900 1499.4600 1318.1900 ;
      RECT 157.4200 1315.9900 1285.6400 1316.0000 ;
      RECT 157.4200 1315.9500 3302.8200 1315.9900 ;
      RECT 1065.1600 1315.5900 3302.8200 1315.9500 ;
      RECT 3368.7200 1314.9200 3370.4200 1316.0000 ;
      RECT 3305.0200 1314.9200 3365.1200 1316.0000 ;
      RECT 2446.4800 1314.9200 3302.8200 1315.5900 ;
      RECT 157.4200 1314.9200 1005.2200 1315.9500 ;
      RECT 5.3000 1314.9200 155.2200 1316.0000 ;
      RECT 0.0000 1314.9200 1.7000 1316.0000 ;
      RECT 1065.1600 1313.7500 1283.0400 1315.5900 ;
      RECT 1011.2200 1313.7500 1059.1600 1315.9500 ;
      RECT 0.0000 1313.7500 1005.2200 1314.9200 ;
      RECT 0.0000 1313.4400 1283.0400 1313.7500 ;
      RECT 2446.4800 1313.3900 3370.4200 1314.9200 ;
      RECT 2392.5400 1313.3900 2440.4800 1315.5900 ;
      RECT 2172.3200 1313.3900 2380.3400 1315.5900 ;
      RECT 1945.9000 1313.3900 2163.9200 1315.5900 ;
      RECT 1731.8800 1313.3900 1939.9000 1315.5900 ;
      RECT 1511.6600 1313.3900 1719.6800 1315.5900 ;
      RECT 1291.4400 1313.3900 1499.4600 1315.5900 ;
      RECT 1.1000 1313.3900 1283.0400 1313.4400 ;
      RECT 1.1000 1313.2800 3370.4200 1313.3900 ;
      RECT 1.1000 1312.5400 5.7000 1313.2800 ;
      RECT 3364.7200 1312.2000 3370.4200 1313.2800 ;
      RECT 3307.6200 1312.2000 3361.1200 1313.2800 ;
      RECT 154.8200 1312.2000 3305.4200 1313.2800 ;
      RECT 9.3000 1312.2000 152.6200 1313.2800 ;
      RECT 0.0000 1312.2000 5.7000 1312.5400 ;
      RECT 0.0000 1310.9800 3370.4200 1312.2000 ;
      RECT 1015.0800 1310.7200 3370.4200 1310.9800 ;
      RECT 2396.3000 1310.5600 3370.4200 1310.7200 ;
      RECT 0.0000 1310.5600 1012.8800 1310.9800 ;
      RECT 1015.0800 1309.9000 1293.0000 1310.7200 ;
      RECT 157.4200 1309.9000 1012.8800 1310.5600 ;
      RECT 2396.3000 1309.6400 3302.8200 1310.5600 ;
      RECT 2176.0800 1309.6400 2394.1000 1310.7200 ;
      RECT 1735.6400 1309.6400 2173.8800 1310.7200 ;
      RECT 1515.4200 1309.6400 1733.4400 1310.7200 ;
      RECT 1295.2000 1309.6400 1513.2200 1310.7200 ;
      RECT 157.4200 1309.6400 1293.0000 1309.9000 ;
      RECT 3368.7200 1309.4800 3370.4200 1310.5600 ;
      RECT 3305.0200 1309.4800 3365.1200 1310.5600 ;
      RECT 157.4200 1309.4800 3302.8200 1309.6400 ;
      RECT 5.3000 1309.4800 155.2200 1310.5600 ;
      RECT 0.0000 1309.4800 1.7000 1310.5600 ;
      RECT 0.0000 1307.8400 3370.4200 1309.4800 ;
      RECT 3364.7200 1306.7600 3370.4200 1307.8400 ;
      RECT 3307.6200 1306.7600 3361.1200 1307.8400 ;
      RECT 154.8200 1306.7600 3305.4200 1307.8400 ;
      RECT 9.3000 1306.7600 152.6200 1307.8400 ;
      RECT 0.0000 1306.7600 5.7000 1307.8400 ;
      RECT 0.0000 1305.1200 3370.4200 1306.7600 ;
      RECT 3368.7200 1304.0400 3370.4200 1305.1200 ;
      RECT 3305.0200 1304.0400 3365.1200 1305.1200 ;
      RECT 157.4200 1304.0400 3302.8200 1305.1200 ;
      RECT 5.3000 1304.0400 155.2200 1305.1200 ;
      RECT 0.0000 1304.0400 1.7000 1305.1200 ;
      RECT 0.0000 1302.4600 3370.4200 1304.0400 ;
      RECT 1.1000 1302.4000 3370.4200 1302.4600 ;
      RECT 1.1000 1301.5600 5.7000 1302.4000 ;
      RECT 3364.7200 1301.3200 3370.4200 1302.4000 ;
      RECT 3307.6200 1301.3200 3361.1200 1302.4000 ;
      RECT 154.8200 1301.3200 3305.4200 1302.4000 ;
      RECT 9.3000 1301.3200 152.6200 1302.4000 ;
      RECT 0.0000 1301.3200 5.7000 1301.5600 ;
      RECT 0.0000 1299.6800 3370.4200 1301.3200 ;
      RECT 3368.7200 1298.6000 3370.4200 1299.6800 ;
      RECT 3305.0200 1298.6000 3365.1200 1299.6800 ;
      RECT 157.4200 1298.6000 3302.8200 1299.6800 ;
      RECT 5.3000 1298.6000 155.2200 1299.6800 ;
      RECT 0.0000 1298.6000 1.7000 1299.6800 ;
      RECT 0.0000 1296.9600 3370.4200 1298.6000 ;
      RECT 3364.7200 1295.8800 3370.4200 1296.9600 ;
      RECT 3307.6200 1295.8800 3361.1200 1296.9600 ;
      RECT 154.8200 1295.8800 3305.4200 1296.9600 ;
      RECT 9.3000 1295.8800 152.6200 1296.9600 ;
      RECT 0.0000 1295.8800 5.7000 1296.9600 ;
      RECT 0.0000 1294.2400 3370.4200 1295.8800 ;
      RECT 3368.7200 1293.1600 3370.4200 1294.2400 ;
      RECT 3305.0200 1293.1600 3365.1200 1294.2400 ;
      RECT 157.4200 1293.1600 3302.8200 1294.2400 ;
      RECT 5.3000 1293.1600 155.2200 1294.2400 ;
      RECT 0.0000 1293.1600 1.7000 1294.2400 ;
      RECT 0.0000 1291.5200 3370.4200 1293.1600 ;
      RECT 0.0000 1291.4800 5.7000 1291.5200 ;
      RECT 1.1000 1290.5800 5.7000 1291.4800 ;
      RECT 3364.7200 1290.4400 3370.4200 1291.5200 ;
      RECT 3307.6200 1290.4400 3361.1200 1291.5200 ;
      RECT 154.8200 1290.4400 3305.4200 1291.5200 ;
      RECT 9.3000 1290.4400 152.6200 1291.5200 ;
      RECT 0.0000 1290.4400 5.7000 1290.5800 ;
      RECT 0.0000 1288.8000 3370.4200 1290.4400 ;
      RECT 3368.7200 1287.7200 3370.4200 1288.8000 ;
      RECT 3305.0200 1287.7200 3365.1200 1288.8000 ;
      RECT 157.4200 1287.7200 3302.8200 1288.8000 ;
      RECT 5.3000 1287.7200 155.2200 1288.8000 ;
      RECT 0.0000 1287.7200 1.7000 1288.8000 ;
      RECT 0.0000 1286.0800 3370.4200 1287.7200 ;
      RECT 3364.7200 1285.0000 3370.4200 1286.0800 ;
      RECT 3307.6200 1285.0000 3361.1200 1286.0800 ;
      RECT 154.8200 1285.0000 3305.4200 1286.0800 ;
      RECT 9.3000 1285.0000 152.6200 1286.0800 ;
      RECT 0.0000 1285.0000 5.7000 1286.0800 ;
      RECT 0.0000 1283.3600 3370.4200 1285.0000 ;
      RECT 3368.7200 1282.2800 3370.4200 1283.3600 ;
      RECT 3305.0200 1282.2800 3365.1200 1283.3600 ;
      RECT 157.4200 1282.2800 3302.8200 1283.3600 ;
      RECT 5.3000 1282.2800 155.2200 1283.3600 ;
      RECT 0.0000 1282.2800 1.7000 1283.3600 ;
      RECT 0.0000 1281.1100 3370.4200 1282.2800 ;
      RECT 1.1000 1280.6400 3370.4200 1281.1100 ;
      RECT 1.1000 1280.2100 5.7000 1280.6400 ;
      RECT 3364.7200 1279.5600 3370.4200 1280.6400 ;
      RECT 3307.6200 1279.5600 3361.1200 1280.6400 ;
      RECT 154.8200 1279.5600 3305.4200 1280.6400 ;
      RECT 9.3000 1279.5600 152.6200 1280.6400 ;
      RECT 0.0000 1279.5600 5.7000 1280.2100 ;
      RECT 0.0000 1277.9200 3370.4200 1279.5600 ;
      RECT 3368.7200 1276.8400 3370.4200 1277.9200 ;
      RECT 3305.0200 1276.8400 3365.1200 1277.9200 ;
      RECT 157.4200 1276.8400 3302.8200 1277.9200 ;
      RECT 5.3000 1276.8400 155.2200 1277.9200 ;
      RECT 0.0000 1276.8400 1.7000 1277.9200 ;
      RECT 0.0000 1275.2000 3370.4200 1276.8400 ;
      RECT 3364.7200 1274.1200 3370.4200 1275.2000 ;
      RECT 3307.6200 1274.1200 3361.1200 1275.2000 ;
      RECT 154.8200 1274.1200 3305.4200 1275.2000 ;
      RECT 9.3000 1274.1200 152.6200 1275.2000 ;
      RECT 0.0000 1274.1200 5.7000 1275.2000 ;
      RECT 0.0000 1272.4800 3370.4200 1274.1200 ;
      RECT 3368.7200 1271.4000 3370.4200 1272.4800 ;
      RECT 3305.0200 1271.4000 3365.1200 1272.4800 ;
      RECT 157.4200 1271.4000 3302.8200 1272.4800 ;
      RECT 5.3000 1271.4000 155.2200 1272.4800 ;
      RECT 0.0000 1271.4000 1.7000 1272.4800 ;
      RECT 0.0000 1270.1300 3370.4200 1271.4000 ;
      RECT 1.1000 1269.7600 3370.4200 1270.1300 ;
      RECT 1.1000 1269.2300 5.7000 1269.7600 ;
      RECT 3364.7200 1268.6800 3370.4200 1269.7600 ;
      RECT 3307.6200 1268.6800 3361.1200 1269.7600 ;
      RECT 154.8200 1268.6800 3305.4200 1269.7600 ;
      RECT 9.3000 1268.6800 152.6200 1269.7600 ;
      RECT 0.0000 1268.6800 5.7000 1269.2300 ;
      RECT 0.0000 1267.0400 3370.4200 1268.6800 ;
      RECT 3368.7200 1265.9600 3370.4200 1267.0400 ;
      RECT 3305.0200 1265.9600 3365.1200 1267.0400 ;
      RECT 157.4200 1265.9600 3302.8200 1267.0400 ;
      RECT 5.3000 1265.9600 155.2200 1267.0400 ;
      RECT 0.0000 1265.9600 1.7000 1267.0400 ;
      RECT 0.0000 1264.3200 3370.4200 1265.9600 ;
      RECT 3364.7200 1263.2400 3370.4200 1264.3200 ;
      RECT 3307.6200 1263.2400 3361.1200 1264.3200 ;
      RECT 154.8200 1263.2400 3305.4200 1264.3200 ;
      RECT 9.3000 1263.2400 152.6200 1264.3200 ;
      RECT 0.0000 1263.2400 5.7000 1264.3200 ;
      RECT 0.0000 1261.6000 3370.4200 1263.2400 ;
      RECT 3368.7200 1260.5200 3370.4200 1261.6000 ;
      RECT 3305.0200 1260.5200 3365.1200 1261.6000 ;
      RECT 157.4200 1260.5200 3302.8200 1261.6000 ;
      RECT 5.3000 1260.5200 155.2200 1261.6000 ;
      RECT 0.0000 1260.5200 1.7000 1261.6000 ;
      RECT 0.0000 1259.1500 3370.4200 1260.5200 ;
      RECT 1.1000 1258.8800 3370.4200 1259.1500 ;
      RECT 1.1000 1258.2500 5.7000 1258.8800 ;
      RECT 3364.7200 1257.8000 3370.4200 1258.8800 ;
      RECT 3307.6200 1257.8000 3361.1200 1258.8800 ;
      RECT 154.8200 1257.8000 3305.4200 1258.8800 ;
      RECT 9.3000 1257.8000 152.6200 1258.8800 ;
      RECT 0.0000 1257.8000 5.7000 1258.2500 ;
      RECT 0.0000 1256.1600 3370.4200 1257.8000 ;
      RECT 3368.7200 1255.0800 3370.4200 1256.1600 ;
      RECT 3305.0200 1255.0800 3365.1200 1256.1600 ;
      RECT 157.4200 1255.0800 3302.8200 1256.1600 ;
      RECT 5.3000 1255.0800 155.2200 1256.1600 ;
      RECT 0.0000 1255.0800 1.7000 1256.1600 ;
      RECT 0.0000 1253.4400 3370.4200 1255.0800 ;
      RECT 3364.7200 1252.3600 3370.4200 1253.4400 ;
      RECT 3307.6200 1252.3600 3361.1200 1253.4400 ;
      RECT 154.8200 1252.3600 3305.4200 1253.4400 ;
      RECT 9.3000 1252.3600 152.6200 1253.4400 ;
      RECT 0.0000 1252.3600 5.7000 1253.4400 ;
      RECT 0.0000 1250.7200 3370.4200 1252.3600 ;
      RECT 3368.7200 1249.6400 3370.4200 1250.7200 ;
      RECT 3305.0200 1249.6400 3365.1200 1250.7200 ;
      RECT 157.4200 1249.6400 3302.8200 1250.7200 ;
      RECT 5.3000 1249.6400 155.2200 1250.7200 ;
      RECT 0.0000 1249.6400 1.7000 1250.7200 ;
      RECT 0.0000 1248.1700 3370.4200 1249.6400 ;
      RECT 1.1000 1248.0000 3370.4200 1248.1700 ;
      RECT 1.1000 1247.2700 5.7000 1248.0000 ;
      RECT 3364.7200 1246.9200 3370.4200 1248.0000 ;
      RECT 3307.6200 1246.9200 3361.1200 1248.0000 ;
      RECT 154.8200 1246.9200 3305.4200 1248.0000 ;
      RECT 9.3000 1246.9200 152.6200 1248.0000 ;
      RECT 0.0000 1246.9200 5.7000 1247.2700 ;
      RECT 0.0000 1245.2800 3370.4200 1246.9200 ;
      RECT 3368.7200 1244.2000 3370.4200 1245.2800 ;
      RECT 3305.0200 1244.2000 3365.1200 1245.2800 ;
      RECT 157.4200 1244.2000 3302.8200 1245.2800 ;
      RECT 5.3000 1244.2000 155.2200 1245.2800 ;
      RECT 0.0000 1244.2000 1.7000 1245.2800 ;
      RECT 0.0000 1242.5600 3370.4200 1244.2000 ;
      RECT 3364.7200 1241.4800 3370.4200 1242.5600 ;
      RECT 3307.6200 1241.4800 3361.1200 1242.5600 ;
      RECT 154.8200 1241.4800 3305.4200 1242.5600 ;
      RECT 9.3000 1241.4800 152.6200 1242.5600 ;
      RECT 0.0000 1241.4800 5.7000 1242.5600 ;
      RECT 0.0000 1239.8400 3370.4200 1241.4800 ;
      RECT 3368.7200 1238.7600 3370.4200 1239.8400 ;
      RECT 3305.0200 1238.7600 3365.1200 1239.8400 ;
      RECT 157.4200 1238.7600 3302.8200 1239.8400 ;
      RECT 5.3000 1238.7600 155.2200 1239.8400 ;
      RECT 0.0000 1238.7600 1.7000 1239.8400 ;
      RECT 0.0000 1237.1900 3370.4200 1238.7600 ;
      RECT 1.1000 1237.1200 3370.4200 1237.1900 ;
      RECT 1.1000 1236.2900 5.7000 1237.1200 ;
      RECT 3364.7200 1236.0400 3370.4200 1237.1200 ;
      RECT 3307.6200 1236.0400 3361.1200 1237.1200 ;
      RECT 154.8200 1236.0400 3305.4200 1237.1200 ;
      RECT 9.3000 1236.0400 152.6200 1237.1200 ;
      RECT 0.0000 1236.0400 5.7000 1236.2900 ;
      RECT 0.0000 1234.4000 3370.4200 1236.0400 ;
      RECT 3368.7200 1233.3200 3370.4200 1234.4000 ;
      RECT 3305.0200 1233.3200 3365.1200 1234.4000 ;
      RECT 157.4200 1233.3200 3302.8200 1234.4000 ;
      RECT 5.3000 1233.3200 155.2200 1234.4000 ;
      RECT 0.0000 1233.3200 1.7000 1234.4000 ;
      RECT 0.0000 1231.6800 3370.4200 1233.3200 ;
      RECT 3364.7200 1230.6000 3370.4200 1231.6800 ;
      RECT 3307.6200 1230.6000 3361.1200 1231.6800 ;
      RECT 154.8200 1230.6000 3305.4200 1231.6800 ;
      RECT 9.3000 1230.6000 152.6200 1231.6800 ;
      RECT 0.0000 1230.6000 5.7000 1231.6800 ;
      RECT 0.0000 1228.9600 3370.4200 1230.6000 ;
      RECT 3368.7200 1227.8800 3370.4200 1228.9600 ;
      RECT 3305.0200 1227.8800 3365.1200 1228.9600 ;
      RECT 157.4200 1227.8800 3302.8200 1228.9600 ;
      RECT 5.3000 1227.8800 155.2200 1228.9600 ;
      RECT 0.0000 1227.8800 1.7000 1228.9600 ;
      RECT 0.0000 1226.2400 3370.4200 1227.8800 ;
      RECT 0.0000 1226.2100 5.7000 1226.2400 ;
      RECT 1.1000 1225.3100 5.7000 1226.2100 ;
      RECT 3364.7200 1225.1600 3370.4200 1226.2400 ;
      RECT 3307.6200 1225.1600 3361.1200 1226.2400 ;
      RECT 154.8200 1225.1600 3305.4200 1226.2400 ;
      RECT 9.3000 1225.1600 152.6200 1226.2400 ;
      RECT 0.0000 1225.1600 5.7000 1225.3100 ;
      RECT 0.0000 1223.5200 3370.4200 1225.1600 ;
      RECT 3368.7200 1222.4400 3370.4200 1223.5200 ;
      RECT 3305.0200 1222.4400 3365.1200 1223.5200 ;
      RECT 157.4200 1222.4400 3302.8200 1223.5200 ;
      RECT 5.3000 1222.4400 155.2200 1223.5200 ;
      RECT 0.0000 1222.4400 1.7000 1223.5200 ;
      RECT 0.0000 1220.8000 3370.4200 1222.4400 ;
      RECT 3364.7200 1219.7200 3370.4200 1220.8000 ;
      RECT 3307.6200 1219.7200 3361.1200 1220.8000 ;
      RECT 154.8200 1219.7200 3305.4200 1220.8000 ;
      RECT 9.3000 1219.7200 152.6200 1220.8000 ;
      RECT 0.0000 1219.7200 5.7000 1220.8000 ;
      RECT 0.0000 1218.0800 3370.4200 1219.7200 ;
      RECT 3368.7200 1217.0000 3370.4200 1218.0800 ;
      RECT 3305.0200 1217.0000 3365.1200 1218.0800 ;
      RECT 157.4200 1217.0000 3302.8200 1218.0800 ;
      RECT 5.3000 1217.0000 155.2200 1218.0800 ;
      RECT 0.0000 1217.0000 1.7000 1218.0800 ;
      RECT 0.0000 1215.8400 3370.4200 1217.0000 ;
      RECT 1.1000 1215.3600 3370.4200 1215.8400 ;
      RECT 1.1000 1214.9400 5.7000 1215.3600 ;
      RECT 3364.7200 1214.2800 3370.4200 1215.3600 ;
      RECT 3307.6200 1214.2800 3361.1200 1215.3600 ;
      RECT 154.8200 1214.2800 3305.4200 1215.3600 ;
      RECT 9.3000 1214.2800 152.6200 1215.3600 ;
      RECT 0.0000 1214.2800 5.7000 1214.9400 ;
      RECT 0.0000 1212.6400 3370.4200 1214.2800 ;
      RECT 3368.7200 1211.5600 3370.4200 1212.6400 ;
      RECT 3305.0200 1211.5600 3365.1200 1212.6400 ;
      RECT 157.4200 1211.5600 3302.8200 1212.6400 ;
      RECT 5.3000 1211.5600 155.2200 1212.6400 ;
      RECT 0.0000 1211.5600 1.7000 1212.6400 ;
      RECT 0.0000 1209.9200 3370.4200 1211.5600 ;
      RECT 3364.7200 1208.8400 3370.4200 1209.9200 ;
      RECT 3307.6200 1208.8400 3361.1200 1209.9200 ;
      RECT 154.8200 1208.8400 3305.4200 1209.9200 ;
      RECT 9.3000 1208.8400 152.6200 1209.9200 ;
      RECT 0.0000 1208.8400 5.7000 1209.9200 ;
      RECT 0.0000 1207.2000 3370.4200 1208.8400 ;
      RECT 3368.7200 1206.1200 3370.4200 1207.2000 ;
      RECT 3305.0200 1206.1200 3365.1200 1207.2000 ;
      RECT 157.4200 1206.1200 3302.8200 1207.2000 ;
      RECT 5.3000 1206.1200 155.2200 1207.2000 ;
      RECT 0.0000 1206.1200 1.7000 1207.2000 ;
      RECT 0.0000 1204.8600 3370.4200 1206.1200 ;
      RECT 1.1000 1204.4800 3370.4200 1204.8600 ;
      RECT 1.1000 1203.9600 5.7000 1204.4800 ;
      RECT 3364.7200 1203.4000 3370.4200 1204.4800 ;
      RECT 3307.6200 1203.4000 3361.1200 1204.4800 ;
      RECT 154.8200 1203.4000 3305.4200 1204.4800 ;
      RECT 9.3000 1203.4000 152.6200 1204.4800 ;
      RECT 0.0000 1203.4000 5.7000 1203.9600 ;
      RECT 0.0000 1201.7600 3370.4200 1203.4000 ;
      RECT 3368.7200 1200.6800 3370.4200 1201.7600 ;
      RECT 3305.0200 1200.6800 3365.1200 1201.7600 ;
      RECT 157.4200 1200.6800 3302.8200 1201.7600 ;
      RECT 5.3000 1200.6800 155.2200 1201.7600 ;
      RECT 0.0000 1200.6800 1.7000 1201.7600 ;
      RECT 0.0000 1199.0400 3370.4200 1200.6800 ;
      RECT 3364.7200 1197.9600 3370.4200 1199.0400 ;
      RECT 3307.6200 1197.9600 3361.1200 1199.0400 ;
      RECT 154.8200 1197.9600 3305.4200 1199.0400 ;
      RECT 9.3000 1197.9600 152.6200 1199.0400 ;
      RECT 0.0000 1197.9600 5.7000 1199.0400 ;
      RECT 0.0000 1196.3200 3370.4200 1197.9600 ;
      RECT 3368.7200 1195.2400 3370.4200 1196.3200 ;
      RECT 3305.0200 1195.2400 3365.1200 1196.3200 ;
      RECT 157.4200 1195.2400 3302.8200 1196.3200 ;
      RECT 5.3000 1195.2400 155.2200 1196.3200 ;
      RECT 0.0000 1195.2400 1.7000 1196.3200 ;
      RECT 0.0000 1193.8800 3370.4200 1195.2400 ;
      RECT 1.1000 1193.6000 3370.4200 1193.8800 ;
      RECT 1.1000 1192.9800 5.7000 1193.6000 ;
      RECT 3364.7200 1192.5200 3370.4200 1193.6000 ;
      RECT 3307.6200 1192.5200 3361.1200 1193.6000 ;
      RECT 154.8200 1192.5200 3305.4200 1193.6000 ;
      RECT 9.3000 1192.5200 152.6200 1193.6000 ;
      RECT 0.0000 1192.5200 5.7000 1192.9800 ;
      RECT 0.0000 1190.8800 3370.4200 1192.5200 ;
      RECT 3368.7200 1189.8000 3370.4200 1190.8800 ;
      RECT 3305.0200 1189.8000 3365.1200 1190.8800 ;
      RECT 157.4200 1189.8000 3302.8200 1190.8800 ;
      RECT 5.3000 1189.8000 155.2200 1190.8800 ;
      RECT 0.0000 1189.8000 1.7000 1190.8800 ;
      RECT 0.0000 1188.1600 3370.4200 1189.8000 ;
      RECT 3364.7200 1187.0800 3370.4200 1188.1600 ;
      RECT 3307.6200 1187.0800 3361.1200 1188.1600 ;
      RECT 154.8200 1187.0800 3305.4200 1188.1600 ;
      RECT 9.3000 1187.0800 152.6200 1188.1600 ;
      RECT 0.0000 1187.0800 5.7000 1188.1600 ;
      RECT 0.0000 1185.4400 3370.4200 1187.0800 ;
      RECT 3368.7200 1184.3600 3370.4200 1185.4400 ;
      RECT 3305.0200 1184.3600 3365.1200 1185.4400 ;
      RECT 157.4200 1184.3600 3302.8200 1185.4400 ;
      RECT 5.3000 1184.3600 155.2200 1185.4400 ;
      RECT 0.0000 1184.3600 1.7000 1185.4400 ;
      RECT 0.0000 1182.9000 3370.4200 1184.3600 ;
      RECT 1.1000 1182.7200 3370.4200 1182.9000 ;
      RECT 1.1000 1182.0000 5.7000 1182.7200 ;
      RECT 3364.7200 1181.6400 3370.4200 1182.7200 ;
      RECT 3307.6200 1181.6400 3361.1200 1182.7200 ;
      RECT 154.8200 1181.6400 3305.4200 1182.7200 ;
      RECT 9.3000 1181.6400 152.6200 1182.7200 ;
      RECT 0.0000 1181.6400 5.7000 1182.0000 ;
      RECT 0.0000 1180.0000 3370.4200 1181.6400 ;
      RECT 3368.7200 1178.9200 3370.4200 1180.0000 ;
      RECT 3305.0200 1178.9200 3365.1200 1180.0000 ;
      RECT 157.4200 1178.9200 3302.8200 1180.0000 ;
      RECT 5.3000 1178.9200 155.2200 1180.0000 ;
      RECT 0.0000 1178.9200 1.7000 1180.0000 ;
      RECT 0.0000 1177.2800 3370.4200 1178.9200 ;
      RECT 3364.7200 1176.2000 3370.4200 1177.2800 ;
      RECT 3307.6200 1176.2000 3361.1200 1177.2800 ;
      RECT 154.8200 1176.2000 3305.4200 1177.2800 ;
      RECT 9.3000 1176.2000 152.6200 1177.2800 ;
      RECT 0.0000 1176.2000 5.7000 1177.2800 ;
      RECT 0.0000 1174.5600 3370.4200 1176.2000 ;
      RECT 3368.7200 1173.4800 3370.4200 1174.5600 ;
      RECT 3305.0200 1173.4800 3365.1200 1174.5600 ;
      RECT 157.4200 1173.4800 3302.8200 1174.5600 ;
      RECT 5.3000 1173.4800 155.2200 1174.5600 ;
      RECT 0.0000 1173.4800 1.7000 1174.5600 ;
      RECT 0.0000 1171.9200 3370.4200 1173.4800 ;
      RECT 1.1000 1171.8400 3370.4200 1171.9200 ;
      RECT 1.1000 1171.0200 5.7000 1171.8400 ;
      RECT 3364.7200 1170.7600 3370.4200 1171.8400 ;
      RECT 3307.6200 1170.7600 3361.1200 1171.8400 ;
      RECT 154.8200 1170.7600 3305.4200 1171.8400 ;
      RECT 9.3000 1170.7600 152.6200 1171.8400 ;
      RECT 0.0000 1170.7600 5.7000 1171.0200 ;
      RECT 0.0000 1169.1200 3370.4200 1170.7600 ;
      RECT 3368.7200 1168.0400 3370.4200 1169.1200 ;
      RECT 3305.0200 1168.0400 3365.1200 1169.1200 ;
      RECT 157.4200 1168.0400 3302.8200 1169.1200 ;
      RECT 5.3000 1168.0400 155.2200 1169.1200 ;
      RECT 0.0000 1168.0400 1.7000 1169.1200 ;
      RECT 0.0000 1166.4000 3370.4200 1168.0400 ;
      RECT 3364.7200 1165.3200 3370.4200 1166.4000 ;
      RECT 3307.6200 1165.3200 3361.1200 1166.4000 ;
      RECT 154.8200 1165.3200 3305.4200 1166.4000 ;
      RECT 9.3000 1165.3200 152.6200 1166.4000 ;
      RECT 0.0000 1165.3200 5.7000 1166.4000 ;
      RECT 0.0000 1163.6800 3370.4200 1165.3200 ;
      RECT 3368.7200 1162.6000 3370.4200 1163.6800 ;
      RECT 3305.0200 1162.6000 3365.1200 1163.6800 ;
      RECT 157.4200 1162.6000 3302.8200 1163.6800 ;
      RECT 5.3000 1162.6000 155.2200 1163.6800 ;
      RECT 0.0000 1162.6000 1.7000 1163.6800 ;
      RECT 0.0000 1161.5500 3370.4200 1162.6000 ;
      RECT 1.1000 1160.9600 3370.4200 1161.5500 ;
      RECT 1.1000 1160.6500 5.7000 1160.9600 ;
      RECT 3364.7200 1159.8800 3370.4200 1160.9600 ;
      RECT 3307.6200 1159.8800 3361.1200 1160.9600 ;
      RECT 154.8200 1159.8800 3305.4200 1160.9600 ;
      RECT 9.3000 1159.8800 152.6200 1160.9600 ;
      RECT 0.0000 1159.8800 5.7000 1160.6500 ;
      RECT 0.0000 1158.2400 3370.4200 1159.8800 ;
      RECT 3368.7200 1157.1600 3370.4200 1158.2400 ;
      RECT 3305.0200 1157.1600 3365.1200 1158.2400 ;
      RECT 157.4200 1157.1600 3302.8200 1158.2400 ;
      RECT 5.3000 1157.1600 155.2200 1158.2400 ;
      RECT 0.0000 1157.1600 1.7000 1158.2400 ;
      RECT 0.0000 1155.5200 3370.4200 1157.1600 ;
      RECT 3364.7200 1154.4400 3370.4200 1155.5200 ;
      RECT 3307.6200 1154.4400 3361.1200 1155.5200 ;
      RECT 154.8200 1154.4400 3305.4200 1155.5200 ;
      RECT 9.3000 1154.4400 152.6200 1155.5200 ;
      RECT 0.0000 1154.4400 5.7000 1155.5200 ;
      RECT 0.0000 1152.8000 3370.4200 1154.4400 ;
      RECT 3368.7200 1151.7200 3370.4200 1152.8000 ;
      RECT 3305.0200 1151.7200 3365.1200 1152.8000 ;
      RECT 157.4200 1151.7200 3302.8200 1152.8000 ;
      RECT 5.3000 1151.7200 155.2200 1152.8000 ;
      RECT 0.0000 1151.7200 1.7000 1152.8000 ;
      RECT 0.0000 1150.5700 3370.4200 1151.7200 ;
      RECT 1.1000 1150.0800 3370.4200 1150.5700 ;
      RECT 1.1000 1149.6700 5.7000 1150.0800 ;
      RECT 3364.7200 1149.0000 3370.4200 1150.0800 ;
      RECT 3307.6200 1149.0000 3361.1200 1150.0800 ;
      RECT 154.8200 1149.0000 3305.4200 1150.0800 ;
      RECT 9.3000 1149.0000 152.6200 1150.0800 ;
      RECT 0.0000 1149.0000 5.7000 1149.6700 ;
      RECT 0.0000 1147.3600 3370.4200 1149.0000 ;
      RECT 3368.7200 1146.2800 3370.4200 1147.3600 ;
      RECT 3305.0200 1146.2800 3365.1200 1147.3600 ;
      RECT 157.4200 1146.2800 3302.8200 1147.3600 ;
      RECT 5.3000 1146.2800 155.2200 1147.3600 ;
      RECT 0.0000 1146.2800 1.7000 1147.3600 ;
      RECT 0.0000 1144.6400 3370.4200 1146.2800 ;
      RECT 3364.7200 1143.5600 3370.4200 1144.6400 ;
      RECT 3307.6200 1143.5600 3361.1200 1144.6400 ;
      RECT 154.8200 1143.5600 3305.4200 1144.6400 ;
      RECT 9.3000 1143.5600 152.6200 1144.6400 ;
      RECT 0.0000 1143.5600 5.7000 1144.6400 ;
      RECT 0.0000 1141.9200 3370.4200 1143.5600 ;
      RECT 3368.7200 1140.8400 3370.4200 1141.9200 ;
      RECT 3305.0200 1140.8400 3365.1200 1141.9200 ;
      RECT 157.4200 1140.8400 3302.8200 1141.9200 ;
      RECT 5.3000 1140.8400 155.2200 1141.9200 ;
      RECT 0.0000 1140.8400 1.7000 1141.9200 ;
      RECT 0.0000 1139.5900 3370.4200 1140.8400 ;
      RECT 1.1000 1139.2000 3370.4200 1139.5900 ;
      RECT 1.1000 1138.6900 5.7000 1139.2000 ;
      RECT 3364.7200 1138.1200 3370.4200 1139.2000 ;
      RECT 3307.6200 1138.1200 3361.1200 1139.2000 ;
      RECT 154.8200 1138.1200 3305.4200 1139.2000 ;
      RECT 9.3000 1138.1200 152.6200 1139.2000 ;
      RECT 0.0000 1138.1200 5.7000 1138.6900 ;
      RECT 0.0000 1136.4800 3370.4200 1138.1200 ;
      RECT 3368.7200 1135.4000 3370.4200 1136.4800 ;
      RECT 3305.0200 1135.4000 3365.1200 1136.4800 ;
      RECT 157.4200 1135.4000 3302.8200 1136.4800 ;
      RECT 5.3000 1135.4000 155.2200 1136.4800 ;
      RECT 0.0000 1135.4000 1.7000 1136.4800 ;
      RECT 0.0000 1133.7600 3370.4200 1135.4000 ;
      RECT 3364.7200 1132.6800 3370.4200 1133.7600 ;
      RECT 3307.6200 1132.6800 3361.1200 1133.7600 ;
      RECT 154.8200 1132.6800 3305.4200 1133.7600 ;
      RECT 9.3000 1132.6800 152.6200 1133.7600 ;
      RECT 0.0000 1132.6800 5.7000 1133.7600 ;
      RECT 0.0000 1131.0400 3370.4200 1132.6800 ;
      RECT 3368.7200 1129.9600 3370.4200 1131.0400 ;
      RECT 3305.0200 1129.9600 3365.1200 1131.0400 ;
      RECT 157.4200 1129.9600 3302.8200 1131.0400 ;
      RECT 5.3000 1129.9600 155.2200 1131.0400 ;
      RECT 0.0000 1129.9600 1.7000 1131.0400 ;
      RECT 0.0000 1128.6100 3370.4200 1129.9600 ;
      RECT 1.1000 1128.3200 3370.4200 1128.6100 ;
      RECT 1.1000 1127.7100 5.7000 1128.3200 ;
      RECT 3364.7200 1127.2400 3370.4200 1128.3200 ;
      RECT 3307.6200 1127.2400 3361.1200 1128.3200 ;
      RECT 154.8200 1127.2400 3305.4200 1128.3200 ;
      RECT 9.3000 1127.2400 152.6200 1128.3200 ;
      RECT 0.0000 1127.2400 5.7000 1127.7100 ;
      RECT 0.0000 1125.6000 3370.4200 1127.2400 ;
      RECT 3368.7200 1124.5200 3370.4200 1125.6000 ;
      RECT 3305.0200 1124.5200 3365.1200 1125.6000 ;
      RECT 157.4200 1124.5200 3302.8200 1125.6000 ;
      RECT 5.3000 1124.5200 155.2200 1125.6000 ;
      RECT 0.0000 1124.5200 1.7000 1125.6000 ;
      RECT 0.0000 1122.8800 3370.4200 1124.5200 ;
      RECT 3364.7200 1121.8000 3370.4200 1122.8800 ;
      RECT 3307.6200 1121.8000 3361.1200 1122.8800 ;
      RECT 154.8200 1121.8000 3305.4200 1122.8800 ;
      RECT 9.3000 1121.8000 152.6200 1122.8800 ;
      RECT 0.0000 1121.8000 5.7000 1122.8800 ;
      RECT 0.0000 1120.1600 3370.4200 1121.8000 ;
      RECT 3368.7200 1119.0800 3370.4200 1120.1600 ;
      RECT 3305.0200 1119.0800 3365.1200 1120.1600 ;
      RECT 157.4200 1119.0800 3302.8200 1120.1600 ;
      RECT 5.3000 1119.0800 155.2200 1120.1600 ;
      RECT 0.0000 1119.0800 1.7000 1120.1600 ;
      RECT 0.0000 1117.6300 3370.4200 1119.0800 ;
      RECT 1.1000 1117.4400 3370.4200 1117.6300 ;
      RECT 1.1000 1116.7300 5.7000 1117.4400 ;
      RECT 3364.7200 1116.3600 3370.4200 1117.4400 ;
      RECT 3307.6200 1116.3600 3361.1200 1117.4400 ;
      RECT 154.8200 1116.3600 3305.4200 1117.4400 ;
      RECT 9.3000 1116.3600 152.6200 1117.4400 ;
      RECT 0.0000 1116.3600 5.7000 1116.7300 ;
      RECT 0.0000 1114.7200 3370.4200 1116.3600 ;
      RECT 3368.7200 1113.6400 3370.4200 1114.7200 ;
      RECT 3305.0200 1113.6400 3365.1200 1114.7200 ;
      RECT 157.4200 1113.6400 3302.8200 1114.7200 ;
      RECT 5.3000 1113.6400 155.2200 1114.7200 ;
      RECT 0.0000 1113.6400 1.7000 1114.7200 ;
      RECT 0.0000 1112.4200 3370.4200 1113.6400 ;
      RECT 1077.7200 1112.1600 3370.4200 1112.4200 ;
      RECT 2436.3200 1112.0000 3370.4200 1112.1600 ;
      RECT 0.0000 1112.0000 1015.2800 1112.4200 ;
      RECT 1077.7200 1111.3400 1295.6000 1112.1600 ;
      RECT 1017.4800 1111.3400 1075.5200 1112.4200 ;
      RECT 154.8200 1111.3400 1015.2800 1112.0000 ;
      RECT 2436.3200 1111.0800 3305.4200 1112.0000 ;
      RECT 2178.6800 1111.0800 2434.1200 1112.1600 ;
      RECT 1958.4600 1111.0800 2176.4800 1112.1600 ;
      RECT 1738.2400 1111.0800 1956.2600 1112.1600 ;
      RECT 1518.0200 1111.0800 1736.0400 1112.1600 ;
      RECT 1297.8000 1111.0800 1515.8200 1112.1600 ;
      RECT 154.8200 1111.0800 1295.6000 1111.3400 ;
      RECT 3364.7200 1110.9200 3370.4200 1112.0000 ;
      RECT 3307.6200 1110.9200 3361.1200 1112.0000 ;
      RECT 154.8200 1110.9200 3305.4200 1111.0800 ;
      RECT 9.3000 1110.9200 152.6200 1112.0000 ;
      RECT 0.0000 1110.9200 5.7000 1112.0000 ;
      RECT 0.0000 1109.3500 3370.4200 1110.9200 ;
      RECT 1285.3800 1109.2800 3370.4200 1109.3500 ;
      RECT 0.0000 1109.2800 1062.9600 1109.3500 ;
      RECT 157.4200 1109.2500 1062.9600 1109.2800 ;
      RECT 1285.3800 1109.0900 3302.8200 1109.2800 ;
      RECT 3368.7200 1108.2000 3370.4200 1109.2800 ;
      RECT 3305.0200 1108.2000 3365.1200 1109.2800 ;
      RECT 2446.4800 1108.2000 3302.8200 1109.0900 ;
      RECT 157.4200 1108.2000 1005.2200 1109.2500 ;
      RECT 5.3000 1108.2000 155.2200 1109.2800 ;
      RECT 0.0000 1108.2000 1.7000 1109.2800 ;
      RECT 0.0000 1107.2600 1005.2200 1108.2000 ;
      RECT 1071.3600 1107.1500 1279.3800 1109.3500 ;
      RECT 1065.1600 1107.0500 1283.0400 1107.1500 ;
      RECT 1011.2200 1107.0500 1059.1600 1109.2500 ;
      RECT 1.1000 1107.0500 1005.2200 1107.2600 ;
      RECT 2446.4800 1106.8900 3370.4200 1108.2000 ;
      RECT 2392.5400 1106.8900 2440.4800 1109.0900 ;
      RECT 2172.3200 1106.8900 2380.3400 1109.0900 ;
      RECT 1952.1000 1106.8900 2160.1200 1109.0900 ;
      RECT 1731.8800 1106.8900 1939.9000 1109.0900 ;
      RECT 1511.6600 1106.8900 1719.6800 1109.0900 ;
      RECT 1291.4400 1106.8900 1499.4600 1109.0900 ;
      RECT 1.1000 1106.8900 1283.0400 1107.0500 ;
      RECT 1.1000 1106.8500 3370.4200 1106.8900 ;
      RECT 1067.7600 1106.7500 3370.4200 1106.8500 ;
      RECT 1287.9800 1106.5600 3370.4200 1106.7500 ;
      RECT 1.1000 1106.5600 1002.6200 1106.8500 ;
      RECT 1287.9800 1106.4900 3305.4200 1106.5600 ;
      RECT 1.1000 1106.3600 5.7000 1106.5600 ;
      RECT 3364.7200 1105.4800 3370.4200 1106.5600 ;
      RECT 3307.6200 1105.4800 3361.1200 1106.5600 ;
      RECT 2449.0800 1105.4800 3305.4200 1106.4900 ;
      RECT 154.8200 1105.4800 1002.6200 1106.5600 ;
      RECT 9.3000 1105.4800 152.6200 1106.5600 ;
      RECT 0.0000 1105.4800 5.7000 1106.3600 ;
      RECT 1011.2200 1104.6500 1059.1600 1106.8500 ;
      RECT 0.0000 1104.6500 1002.6200 1105.4800 ;
      RECT 1071.3600 1104.5500 1279.3800 1106.7500 ;
      RECT 0.0000 1104.5500 1065.5600 1104.6500 ;
      RECT 2449.0800 1104.2900 3370.4200 1105.4800 ;
      RECT 2392.5400 1104.2900 2440.4800 1106.4900 ;
      RECT 2172.3200 1104.2900 2380.3400 1106.4900 ;
      RECT 1952.1000 1104.2900 2166.5200 1106.4900 ;
      RECT 1731.8800 1104.2900 1939.9000 1106.4900 ;
      RECT 1511.6600 1104.2900 1719.6800 1106.4900 ;
      RECT 1291.4400 1104.2900 1505.8600 1106.4900 ;
      RECT 0.0000 1104.2900 1285.6400 1104.5500 ;
      RECT 0.0000 1103.8400 3370.4200 1104.2900 ;
      RECT 3368.7200 1102.7600 3370.4200 1103.8400 ;
      RECT 3305.0200 1102.7600 3365.1200 1103.8400 ;
      RECT 157.4200 1102.7600 3302.8200 1103.8400 ;
      RECT 5.3000 1102.7600 155.2200 1103.8400 ;
      RECT 0.0000 1102.7600 1.7000 1103.8400 ;
      RECT 0.0000 1101.1200 3370.4200 1102.7600 ;
      RECT 3364.7200 1100.0400 3370.4200 1101.1200 ;
      RECT 3307.6200 1100.0400 3361.1200 1101.1200 ;
      RECT 154.8200 1100.0400 3305.4200 1101.1200 ;
      RECT 9.3000 1100.0400 152.6200 1101.1200 ;
      RECT 0.0000 1100.0400 5.7000 1101.1200 ;
      RECT 0.0000 1099.3200 3370.4200 1100.0400 ;
      RECT 1285.3800 1099.0600 3370.4200 1099.3200 ;
      RECT 2446.4800 1098.4000 3370.4200 1099.0600 ;
      RECT 3368.7200 1097.3200 3370.4200 1098.4000 ;
      RECT 3305.0200 1097.3200 3365.1200 1098.4000 ;
      RECT 2446.4800 1097.3200 3302.8200 1098.4000 ;
      RECT 167.4150 1097.1200 953.1450 1099.3200 ;
      RECT 0.0000 1097.1200 1.7000 1099.3200 ;
      RECT 2446.4800 1096.8600 3370.4200 1097.3200 ;
      RECT 0.0000 1096.8600 1283.0400 1097.1200 ;
      RECT 0.0000 1096.8200 3370.4200 1096.8600 ;
      RECT 1065.0600 1096.7200 3370.4200 1096.8200 ;
      RECT 0.0000 1096.7200 1062.6600 1096.8200 ;
      RECT 1287.9800 1096.5600 3370.4200 1096.7200 ;
      RECT 1945.8000 1096.4600 3370.4200 1096.5600 ;
      RECT 1287.9800 1096.4600 1943.4000 1096.5600 ;
      RECT 0.0000 1096.2800 5.7000 1096.7200 ;
      RECT 2449.0800 1095.6800 3370.4200 1096.4600 ;
      RECT 1.1000 1095.3800 5.7000 1096.2800 ;
      RECT 3364.7200 1094.6000 3370.4200 1095.6800 ;
      RECT 3307.6200 1094.6000 3361.1200 1095.6800 ;
      RECT 2449.0800 1094.6000 3305.4200 1095.6800 ;
      RECT 167.4150 1094.5200 953.1450 1096.7200 ;
      RECT 0.0000 1094.5200 5.7000 1095.3800 ;
      RECT 2449.0800 1094.2600 3370.4200 1094.6000 ;
      RECT 1065.0600 1094.2600 1285.6400 1094.5200 ;
      RECT 1945.8000 1092.9600 3370.4200 1094.2600 ;
      RECT 0.0000 1092.9600 1062.6600 1094.5200 ;
      RECT 1065.0600 1092.8200 1943.4000 1094.2600 ;
      RECT 157.4200 1092.8200 1062.6600 1092.9600 ;
      RECT 1945.8000 1092.5600 3302.8200 1092.9600 ;
      RECT 157.4200 1092.5600 1943.4000 1092.8200 ;
      RECT 3368.7200 1091.8800 3370.4200 1092.9600 ;
      RECT 3305.0200 1091.8800 3365.1200 1092.9600 ;
      RECT 157.4200 1091.8800 3302.8200 1092.5600 ;
      RECT 5.3000 1091.8800 155.2200 1092.9600 ;
      RECT 0.0000 1091.8800 1.7000 1092.9600 ;
      RECT 0.0000 1090.2400 3370.4200 1091.8800 ;
      RECT 154.8200 1089.8600 3305.4200 1090.2400 ;
      RECT 1287.9800 1089.6000 3305.4200 1089.8600 ;
      RECT 3364.7200 1089.1600 3370.4200 1090.2400 ;
      RECT 3307.6200 1089.1600 3361.1200 1090.2400 ;
      RECT 2168.7200 1089.1600 3305.4200 1089.6000 ;
      RECT 154.8200 1089.1600 1065.5600 1089.8600 ;
      RECT 9.3000 1089.1600 152.6200 1090.2400 ;
      RECT 0.0000 1089.1600 5.7000 1090.2400 ;
      RECT 0.0000 1088.7100 1065.5600 1089.1600 ;
      RECT 2168.7200 1088.5500 3370.4200 1089.1600 ;
      RECT 1287.9800 1088.5500 1946.3000 1089.6000 ;
      RECT 1071.3600 1087.6600 1279.3800 1089.8600 ;
      RECT 1062.4600 1087.6600 1065.5600 1088.7100 ;
      RECT 2449.0800 1087.5200 3370.4200 1088.5500 ;
      RECT 0.0000 1087.5200 1002.6200 1088.7100 ;
      RECT 1952.1000 1087.4000 2160.1200 1089.6000 ;
      RECT 1943.2000 1087.4000 1946.3000 1088.5500 ;
      RECT 1062.4600 1087.2600 1285.6400 1087.6600 ;
      RECT 1943.2000 1087.0000 2166.5200 1087.4000 ;
      RECT 1062.4600 1086.5100 1062.9600 1087.2600 ;
      RECT 1011.2200 1086.5100 1059.1600 1088.7100 ;
      RECT 157.4200 1086.5100 1002.6200 1087.5200 ;
      RECT 3368.7200 1086.4400 3370.4200 1087.5200 ;
      RECT 3305.0200 1086.4400 3365.1200 1087.5200 ;
      RECT 2449.0800 1086.4400 3302.8200 1087.5200 ;
      RECT 157.4200 1086.4400 1062.9600 1086.5100 ;
      RECT 5.3000 1086.4400 155.2200 1087.5200 ;
      RECT 0.0000 1086.4400 1.7000 1087.5200 ;
      RECT 2449.0800 1086.3500 3370.4200 1086.4400 ;
      RECT 2392.5400 1086.3500 2440.4800 1088.5500 ;
      RECT 2172.3200 1086.3500 2380.3400 1088.5500 ;
      RECT 2166.1200 1086.3500 2166.5200 1087.0000 ;
      RECT 1943.2000 1086.3500 1943.7000 1087.0000 ;
      RECT 1731.8800 1086.3500 1939.9000 1088.5500 ;
      RECT 1511.6600 1086.3500 1719.6800 1088.5500 ;
      RECT 1291.4400 1086.3500 1499.4600 1088.5500 ;
      RECT 1285.3800 1086.3500 1285.6400 1087.2600 ;
      RECT 0.0000 1086.3100 1062.9600 1086.4400 ;
      RECT 2166.1200 1085.9500 3370.4200 1086.3500 ;
      RECT 1285.3800 1085.9500 1943.7000 1086.3500 ;
      RECT 0.0000 1085.3000 1005.2200 1086.3100 ;
      RECT 1071.3600 1085.0600 1279.3800 1087.2600 ;
      RECT 2446.4800 1084.8000 3370.4200 1085.9500 ;
      RECT 1952.1000 1084.8000 2160.1200 1087.0000 ;
      RECT 1.1000 1084.8000 1005.2200 1085.3000 ;
      RECT 1.1000 1084.4000 5.7000 1084.8000 ;
      RECT 1065.1600 1084.1100 1283.0400 1085.0600 ;
      RECT 1011.2200 1084.1100 1059.1600 1086.3100 ;
      RECT 154.8200 1084.1100 1005.2200 1084.8000 ;
      RECT 2446.4800 1083.7500 3305.4200 1084.8000 ;
      RECT 2392.5400 1083.7500 2440.4800 1085.9500 ;
      RECT 2172.3200 1083.7500 2380.3400 1085.9500 ;
      RECT 1945.9000 1083.7500 2163.9200 1084.8000 ;
      RECT 1731.8800 1083.7500 1939.9000 1085.9500 ;
      RECT 1511.6600 1083.7500 1719.6800 1085.9500 ;
      RECT 1291.4400 1083.7500 1499.4600 1085.9500 ;
      RECT 154.8200 1083.7500 1283.0400 1084.1100 ;
      RECT 3364.7200 1083.7200 3370.4200 1084.8000 ;
      RECT 3307.6200 1083.7200 3361.1200 1084.8000 ;
      RECT 154.8200 1083.7200 3305.4200 1083.7500 ;
      RECT 9.3000 1083.7200 152.6200 1084.8000 ;
      RECT 0.0000 1083.7200 5.7000 1084.4000 ;
      RECT 0.0000 1082.0800 3370.4200 1083.7200 ;
      RECT 157.4200 1081.3400 3302.8200 1082.0800 ;
      RECT 1057.5000 1081.0800 3302.8200 1081.3400 ;
      RECT 3368.7200 1081.0000 3370.4200 1082.0800 ;
      RECT 3305.0200 1081.0000 3365.1200 1082.0800 ;
      RECT 2396.3000 1081.0000 3302.8200 1081.0800 ;
      RECT 157.4200 1081.0000 1055.3000 1081.3400 ;
      RECT 5.3000 1081.0000 155.2200 1082.0800 ;
      RECT 0.0000 1081.0000 1.7000 1082.0800 ;
      RECT 1057.5000 1080.2600 1293.0000 1081.0800 ;
      RECT 0.0000 1080.2600 1055.3000 1081.0000 ;
      RECT 0.0000 1080.1800 1293.0000 1080.2600 ;
      RECT 2396.3000 1080.0000 3370.4200 1081.0000 ;
      RECT 2176.0800 1080.0000 2394.1000 1081.0800 ;
      RECT 1735.6400 1080.0000 2173.8800 1081.0800 ;
      RECT 1515.4200 1080.0000 1733.4400 1081.0800 ;
      RECT 1295.2000 1080.0000 1513.2200 1081.0800 ;
      RECT 1075.1200 1080.0000 1293.0000 1080.1800 ;
      RECT 1075.1200 1079.9200 3370.4200 1080.0000 ;
      RECT 1955.8600 1079.3600 3370.4200 1079.9200 ;
      RECT 0.0000 1079.3600 1072.9200 1080.1800 ;
      RECT 1075.1200 1079.1000 1953.6600 1079.9200 ;
      RECT 154.8200 1079.1000 1072.9200 1079.3600 ;
      RECT 1955.8600 1078.8400 3305.4200 1079.3600 ;
      RECT 154.8200 1078.8400 1953.6600 1079.1000 ;
      RECT 3364.7200 1078.2800 3370.4200 1079.3600 ;
      RECT 3307.6200 1078.2800 3361.1200 1079.3600 ;
      RECT 154.8200 1078.2800 3305.4200 1078.8400 ;
      RECT 9.3000 1078.2800 152.6200 1079.3600 ;
      RECT 0.0000 1078.2800 5.7000 1079.3600 ;
      RECT 0.0000 1076.6400 3370.4200 1078.2800 ;
      RECT 3368.7200 1075.5600 3370.4200 1076.6400 ;
      RECT 3305.0200 1075.5600 3365.1200 1076.6400 ;
      RECT 157.4200 1075.5600 3302.8200 1076.6400 ;
      RECT 5.3000 1075.5600 155.2200 1076.6400 ;
      RECT 0.0000 1075.5600 1.7000 1076.6400 ;
      RECT 0.0000 1074.3200 3370.4200 1075.5600 ;
      RECT 1.1000 1073.9200 3370.4200 1074.3200 ;
      RECT 1.1000 1073.4200 5.7000 1073.9200 ;
      RECT 3364.7200 1072.8400 3370.4200 1073.9200 ;
      RECT 3307.6200 1072.8400 3361.1200 1073.9200 ;
      RECT 154.8200 1072.8400 3305.4200 1073.9200 ;
      RECT 9.3000 1072.8400 152.6200 1073.9200 ;
      RECT 0.0000 1072.8400 5.7000 1073.4200 ;
      RECT 0.0000 1071.2000 3370.4200 1072.8400 ;
      RECT 3368.7200 1070.1200 3370.4200 1071.2000 ;
      RECT 3305.0200 1070.1200 3365.1200 1071.2000 ;
      RECT 157.4200 1070.1200 3302.8200 1071.2000 ;
      RECT 5.3000 1070.1200 155.2200 1071.2000 ;
      RECT 0.0000 1070.1200 1.7000 1071.2000 ;
      RECT 0.0000 1068.4800 3370.4200 1070.1200 ;
      RECT 3364.7200 1067.4000 3370.4200 1068.4800 ;
      RECT 3307.6200 1067.4000 3361.1200 1068.4800 ;
      RECT 154.8200 1067.4000 3305.4200 1068.4800 ;
      RECT 9.3000 1067.4000 152.6200 1068.4800 ;
      RECT 0.0000 1067.4000 5.7000 1068.4800 ;
      RECT 0.0000 1065.7600 3370.4200 1067.4000 ;
      RECT 3368.7200 1064.6800 3370.4200 1065.7600 ;
      RECT 3305.0200 1064.6800 3365.1200 1065.7600 ;
      RECT 157.4200 1064.6800 3302.8200 1065.7600 ;
      RECT 5.3000 1064.6800 155.2200 1065.7600 ;
      RECT 0.0000 1064.6800 1.7000 1065.7600 ;
      RECT 0.0000 1063.3400 3370.4200 1064.6800 ;
      RECT 1.1000 1063.0400 3370.4200 1063.3400 ;
      RECT 1.1000 1062.4400 5.7000 1063.0400 ;
      RECT 3364.7200 1061.9600 3370.4200 1063.0400 ;
      RECT 3307.6200 1061.9600 3361.1200 1063.0400 ;
      RECT 154.8200 1061.9600 3305.4200 1063.0400 ;
      RECT 9.3000 1061.9600 152.6200 1063.0400 ;
      RECT 0.0000 1061.9600 5.7000 1062.4400 ;
      RECT 0.0000 1060.3200 3370.4200 1061.9600 ;
      RECT 3368.7200 1059.2400 3370.4200 1060.3200 ;
      RECT 3305.0200 1059.2400 3365.1200 1060.3200 ;
      RECT 157.4200 1059.2400 3302.8200 1060.3200 ;
      RECT 5.3000 1059.2400 155.2200 1060.3200 ;
      RECT 0.0000 1059.2400 1.7000 1060.3200 ;
      RECT 0.0000 1057.6000 3370.4200 1059.2400 ;
      RECT 3364.7200 1056.5200 3370.4200 1057.6000 ;
      RECT 3307.6200 1056.5200 3361.1200 1057.6000 ;
      RECT 154.8200 1056.5200 3305.4200 1057.6000 ;
      RECT 9.3000 1056.5200 152.6200 1057.6000 ;
      RECT 0.0000 1056.5200 5.7000 1057.6000 ;
      RECT 0.0000 1054.8800 3370.4200 1056.5200 ;
      RECT 3368.7200 1053.8000 3370.4200 1054.8800 ;
      RECT 3305.0200 1053.8000 3365.1200 1054.8800 ;
      RECT 157.4200 1053.8000 3302.8200 1054.8800 ;
      RECT 5.3000 1053.8000 155.2200 1054.8800 ;
      RECT 0.0000 1053.8000 1.7000 1054.8800 ;
      RECT 0.0000 1052.9700 3370.4200 1053.8000 ;
      RECT 1.1000 1052.1600 3370.4200 1052.9700 ;
      RECT 1.1000 1052.0700 5.7000 1052.1600 ;
      RECT 3364.7200 1051.0800 3370.4200 1052.1600 ;
      RECT 3307.6200 1051.0800 3361.1200 1052.1600 ;
      RECT 154.8200 1051.0800 3305.4200 1052.1600 ;
      RECT 9.3000 1051.0800 152.6200 1052.1600 ;
      RECT 0.0000 1051.0800 5.7000 1052.0700 ;
      RECT 0.0000 1049.4400 3370.4200 1051.0800 ;
      RECT 3368.7200 1048.3600 3370.4200 1049.4400 ;
      RECT 3305.0200 1048.3600 3365.1200 1049.4400 ;
      RECT 157.4200 1048.3600 3302.8200 1049.4400 ;
      RECT 5.3000 1048.3600 155.2200 1049.4400 ;
      RECT 0.0000 1048.3600 1.7000 1049.4400 ;
      RECT 0.0000 1046.7200 3370.4200 1048.3600 ;
      RECT 3364.7200 1045.6400 3370.4200 1046.7200 ;
      RECT 3307.6200 1045.6400 3361.1200 1046.7200 ;
      RECT 154.8200 1045.6400 3305.4200 1046.7200 ;
      RECT 9.3000 1045.6400 152.6200 1046.7200 ;
      RECT 0.0000 1045.6400 5.7000 1046.7200 ;
      RECT 0.0000 1044.0000 3370.4200 1045.6400 ;
      RECT 3368.7200 1042.9200 3370.4200 1044.0000 ;
      RECT 3305.0200 1042.9200 3365.1200 1044.0000 ;
      RECT 157.4200 1042.9200 3302.8200 1044.0000 ;
      RECT 5.3000 1042.9200 155.2200 1044.0000 ;
      RECT 0.0000 1042.9200 1.7000 1044.0000 ;
      RECT 0.0000 1041.9900 3370.4200 1042.9200 ;
      RECT 1.1000 1041.2800 3370.4200 1041.9900 ;
      RECT 1.1000 1041.0900 5.7000 1041.2800 ;
      RECT 3364.7200 1040.2000 3370.4200 1041.2800 ;
      RECT 3307.6200 1040.2000 3361.1200 1041.2800 ;
      RECT 154.8200 1040.2000 3305.4200 1041.2800 ;
      RECT 9.3000 1040.2000 152.6200 1041.2800 ;
      RECT 0.0000 1040.2000 5.7000 1041.0900 ;
      RECT 0.0000 1038.5600 3370.4200 1040.2000 ;
      RECT 3368.7200 1037.4800 3370.4200 1038.5600 ;
      RECT 3305.0200 1037.4800 3365.1200 1038.5600 ;
      RECT 157.4200 1037.4800 3302.8200 1038.5600 ;
      RECT 5.3000 1037.4800 155.2200 1038.5600 ;
      RECT 0.0000 1037.4800 1.7000 1038.5600 ;
      RECT 0.0000 1035.8400 3370.4200 1037.4800 ;
      RECT 3364.7200 1034.7600 3370.4200 1035.8400 ;
      RECT 3307.6200 1034.7600 3361.1200 1035.8400 ;
      RECT 154.8200 1034.7600 3305.4200 1035.8400 ;
      RECT 9.3000 1034.7600 152.6200 1035.8400 ;
      RECT 0.0000 1034.7600 5.7000 1035.8400 ;
      RECT 0.0000 1033.1200 3370.4200 1034.7600 ;
      RECT 3368.7200 1032.0400 3370.4200 1033.1200 ;
      RECT 3305.0200 1032.0400 3365.1200 1033.1200 ;
      RECT 157.4200 1032.0400 3302.8200 1033.1200 ;
      RECT 5.3000 1032.0400 155.2200 1033.1200 ;
      RECT 0.0000 1032.0400 1.7000 1033.1200 ;
      RECT 0.0000 1031.0100 3370.4200 1032.0400 ;
      RECT 1.1000 1030.4000 3370.4200 1031.0100 ;
      RECT 1.1000 1030.1100 5.7000 1030.4000 ;
      RECT 3364.7200 1029.3200 3370.4200 1030.4000 ;
      RECT 3307.6200 1029.3200 3361.1200 1030.4000 ;
      RECT 154.8200 1029.3200 3305.4200 1030.4000 ;
      RECT 9.3000 1029.3200 152.6200 1030.4000 ;
      RECT 0.0000 1029.3200 5.7000 1030.1100 ;
      RECT 0.0000 1027.6800 3370.4200 1029.3200 ;
      RECT 3368.7200 1026.6000 3370.4200 1027.6800 ;
      RECT 3305.0200 1026.6000 3365.1200 1027.6800 ;
      RECT 157.4200 1026.6000 3302.8200 1027.6800 ;
      RECT 5.3000 1026.6000 155.2200 1027.6800 ;
      RECT 0.0000 1026.6000 1.7000 1027.6800 ;
      RECT 0.0000 1024.9600 3370.4200 1026.6000 ;
      RECT 3364.7200 1023.8800 3370.4200 1024.9600 ;
      RECT 3307.6200 1023.8800 3361.1200 1024.9600 ;
      RECT 154.8200 1023.8800 3305.4200 1024.9600 ;
      RECT 9.3000 1023.8800 152.6200 1024.9600 ;
      RECT 0.0000 1023.8800 5.7000 1024.9600 ;
      RECT 0.0000 1022.2400 3370.4200 1023.8800 ;
      RECT 3368.7200 1021.1600 3370.4200 1022.2400 ;
      RECT 3305.0200 1021.1600 3365.1200 1022.2400 ;
      RECT 157.4200 1021.1600 3302.8200 1022.2400 ;
      RECT 5.3000 1021.1600 155.2200 1022.2400 ;
      RECT 0.0000 1021.1600 1.7000 1022.2400 ;
      RECT 0.0000 1020.0300 3370.4200 1021.1600 ;
      RECT 1.1000 1019.5200 3370.4200 1020.0300 ;
      RECT 1.1000 1019.1300 5.7000 1019.5200 ;
      RECT 3364.7200 1018.4400 3370.4200 1019.5200 ;
      RECT 3307.6200 1018.4400 3361.1200 1019.5200 ;
      RECT 154.8200 1018.4400 3305.4200 1019.5200 ;
      RECT 9.3000 1018.4400 152.6200 1019.5200 ;
      RECT 0.0000 1018.4400 5.7000 1019.1300 ;
      RECT 0.0000 1016.8000 3370.4200 1018.4400 ;
      RECT 3368.7200 1015.7200 3370.4200 1016.8000 ;
      RECT 3305.0200 1015.7200 3365.1200 1016.8000 ;
      RECT 157.4200 1015.7200 3302.8200 1016.8000 ;
      RECT 5.3000 1015.7200 155.2200 1016.8000 ;
      RECT 0.0000 1015.7200 1.7000 1016.8000 ;
      RECT 0.0000 1014.0800 3370.4200 1015.7200 ;
      RECT 3364.7200 1013.0000 3370.4200 1014.0800 ;
      RECT 3307.6200 1013.0000 3361.1200 1014.0800 ;
      RECT 154.8200 1013.0000 3305.4200 1014.0800 ;
      RECT 9.3000 1013.0000 152.6200 1014.0800 ;
      RECT 0.0000 1013.0000 5.7000 1014.0800 ;
      RECT 0.0000 1011.3600 3370.4200 1013.0000 ;
      RECT 3368.7200 1010.2800 3370.4200 1011.3600 ;
      RECT 3305.0200 1010.2800 3365.1200 1011.3600 ;
      RECT 157.4200 1010.2800 3302.8200 1011.3600 ;
      RECT 5.3000 1010.2800 155.2200 1011.3600 ;
      RECT 0.0000 1010.2800 1.7000 1011.3600 ;
      RECT 0.0000 1009.0500 3370.4200 1010.2800 ;
      RECT 1.1000 1008.6400 3370.4200 1009.0500 ;
      RECT 1.1000 1008.1500 5.7000 1008.6400 ;
      RECT 3364.7200 1007.5600 3370.4200 1008.6400 ;
      RECT 3307.6200 1007.5600 3361.1200 1008.6400 ;
      RECT 154.8200 1007.5600 3305.4200 1008.6400 ;
      RECT 9.3000 1007.5600 152.6200 1008.6400 ;
      RECT 0.0000 1007.5600 5.7000 1008.1500 ;
      RECT 0.0000 1005.9200 3370.4200 1007.5600 ;
      RECT 3368.7200 1004.8400 3370.4200 1005.9200 ;
      RECT 3305.0200 1004.8400 3365.1200 1005.9200 ;
      RECT 157.4200 1004.8400 3302.8200 1005.9200 ;
      RECT 5.3000 1004.8400 155.2200 1005.9200 ;
      RECT 0.0000 1004.8400 1.7000 1005.9200 ;
      RECT 0.0000 1003.2000 3370.4200 1004.8400 ;
      RECT 3364.7200 1002.1200 3370.4200 1003.2000 ;
      RECT 3307.6200 1002.1200 3361.1200 1003.2000 ;
      RECT 154.8200 1002.1200 3305.4200 1003.2000 ;
      RECT 9.3000 1002.1200 152.6200 1003.2000 ;
      RECT 0.0000 1002.1200 5.7000 1003.2000 ;
      RECT 0.0000 1000.4800 3370.4200 1002.1200 ;
      RECT 3368.7200 999.4000 3370.4200 1000.4800 ;
      RECT 3305.0200 999.4000 3365.1200 1000.4800 ;
      RECT 157.4200 999.4000 3302.8200 1000.4800 ;
      RECT 5.3000 999.4000 155.2200 1000.4800 ;
      RECT 0.0000 999.4000 1.7000 1000.4800 ;
      RECT 0.0000 998.6800 3370.4200 999.4000 ;
      RECT 1.1000 997.7800 3370.4200 998.6800 ;
      RECT 0.0000 997.7600 3370.4200 997.7800 ;
      RECT 3364.7200 996.6800 3370.4200 997.7600 ;
      RECT 3307.6200 996.6800 3361.1200 997.7600 ;
      RECT 154.8200 996.6800 3305.4200 997.7600 ;
      RECT 9.3000 996.6800 152.6200 997.7600 ;
      RECT 0.0000 996.6800 5.7000 997.7600 ;
      RECT 0.0000 995.0400 3370.4200 996.6800 ;
      RECT 3368.7200 993.9600 3370.4200 995.0400 ;
      RECT 3305.0200 993.9600 3365.1200 995.0400 ;
      RECT 157.4200 993.9600 3302.8200 995.0400 ;
      RECT 5.3000 993.9600 155.2200 995.0400 ;
      RECT 0.0000 993.9600 1.7000 995.0400 ;
      RECT 0.0000 992.3200 3370.4200 993.9600 ;
      RECT 3364.7200 991.2400 3370.4200 992.3200 ;
      RECT 3307.6200 991.2400 3361.1200 992.3200 ;
      RECT 154.8200 991.2400 3305.4200 992.3200 ;
      RECT 9.3000 991.2400 152.6200 992.3200 ;
      RECT 0.0000 991.2400 5.7000 992.3200 ;
      RECT 0.0000 989.6000 3370.4200 991.2400 ;
      RECT 3368.7200 988.5200 3370.4200 989.6000 ;
      RECT 3305.0200 988.5200 3365.1200 989.6000 ;
      RECT 157.4200 988.5200 3302.8200 989.6000 ;
      RECT 5.3000 988.5200 155.2200 989.6000 ;
      RECT 0.0000 988.5200 1.7000 989.6000 ;
      RECT 0.0000 987.7000 3370.4200 988.5200 ;
      RECT 1.1000 986.8800 3370.4200 987.7000 ;
      RECT 1.1000 986.8000 5.7000 986.8800 ;
      RECT 3364.7200 985.8000 3370.4200 986.8800 ;
      RECT 3307.6200 985.8000 3361.1200 986.8800 ;
      RECT 154.8200 985.8000 3305.4200 986.8800 ;
      RECT 9.3000 985.8000 152.6200 986.8800 ;
      RECT 0.0000 985.8000 5.7000 986.8000 ;
      RECT 0.0000 984.1600 3370.4200 985.8000 ;
      RECT 3368.7200 983.0800 3370.4200 984.1600 ;
      RECT 3305.0200 983.0800 3365.1200 984.1600 ;
      RECT 157.4200 983.0800 3302.8200 984.1600 ;
      RECT 5.3000 983.0800 155.2200 984.1600 ;
      RECT 0.0000 983.0800 1.7000 984.1600 ;
      RECT 0.0000 981.4400 3370.4200 983.0800 ;
      RECT 3364.7200 980.3600 3370.4200 981.4400 ;
      RECT 3307.6200 980.3600 3361.1200 981.4400 ;
      RECT 154.8200 980.3600 3305.4200 981.4400 ;
      RECT 9.3000 980.3600 152.6200 981.4400 ;
      RECT 0.0000 980.3600 5.7000 981.4400 ;
      RECT 0.0000 978.7200 3370.4200 980.3600 ;
      RECT 3368.7200 977.6400 3370.4200 978.7200 ;
      RECT 3305.0200 977.6400 3365.1200 978.7200 ;
      RECT 157.4200 977.6400 3302.8200 978.7200 ;
      RECT 5.3000 977.6400 155.2200 978.7200 ;
      RECT 0.0000 977.6400 1.7000 978.7200 ;
      RECT 0.0000 976.7200 3370.4200 977.6400 ;
      RECT 1.1000 976.0000 3370.4200 976.7200 ;
      RECT 1.1000 975.8200 5.7000 976.0000 ;
      RECT 3364.7200 974.9200 3370.4200 976.0000 ;
      RECT 3307.6200 974.9200 3361.1200 976.0000 ;
      RECT 154.8200 974.9200 3305.4200 976.0000 ;
      RECT 9.3000 974.9200 152.6200 976.0000 ;
      RECT 0.0000 974.9200 5.7000 975.8200 ;
      RECT 0.0000 973.2800 3370.4200 974.9200 ;
      RECT 3368.7200 972.2000 3370.4200 973.2800 ;
      RECT 3305.0200 972.2000 3365.1200 973.2800 ;
      RECT 157.4200 972.2000 3302.8200 973.2800 ;
      RECT 5.3000 972.2000 155.2200 973.2800 ;
      RECT 0.0000 972.2000 1.7000 973.2800 ;
      RECT 0.0000 970.5600 3370.4200 972.2000 ;
      RECT 3364.7200 969.4800 3370.4200 970.5600 ;
      RECT 3307.6200 969.4800 3361.1200 970.5600 ;
      RECT 154.8200 969.4800 3305.4200 970.5600 ;
      RECT 9.3000 969.4800 152.6200 970.5600 ;
      RECT 0.0000 969.4800 5.7000 970.5600 ;
      RECT 0.0000 967.8400 3370.4200 969.4800 ;
      RECT 3368.7200 966.7600 3370.4200 967.8400 ;
      RECT 3305.0200 966.7600 3365.1200 967.8400 ;
      RECT 157.4200 966.7600 3302.8200 967.8400 ;
      RECT 5.3000 966.7600 155.2200 967.8400 ;
      RECT 0.0000 966.7600 1.7000 967.8400 ;
      RECT 0.0000 965.7400 3370.4200 966.7600 ;
      RECT 1.1000 965.1200 3370.4200 965.7400 ;
      RECT 1.1000 964.8400 5.7000 965.1200 ;
      RECT 3364.7200 964.0400 3370.4200 965.1200 ;
      RECT 3307.6200 964.0400 3361.1200 965.1200 ;
      RECT 154.8200 964.0400 3305.4200 965.1200 ;
      RECT 9.3000 964.0400 152.6200 965.1200 ;
      RECT 0.0000 964.0400 5.7000 964.8400 ;
      RECT 0.0000 962.4000 3370.4200 964.0400 ;
      RECT 3368.7200 961.3200 3370.4200 962.4000 ;
      RECT 3305.0200 961.3200 3365.1200 962.4000 ;
      RECT 157.4200 961.3200 3302.8200 962.4000 ;
      RECT 5.3000 961.3200 155.2200 962.4000 ;
      RECT 0.0000 961.3200 1.7000 962.4000 ;
      RECT 0.0000 959.6800 3370.4200 961.3200 ;
      RECT 3364.7200 958.6000 3370.4200 959.6800 ;
      RECT 3307.6200 958.6000 3361.1200 959.6800 ;
      RECT 154.8200 958.6000 3305.4200 959.6800 ;
      RECT 9.3000 958.6000 152.6200 959.6800 ;
      RECT 0.0000 958.6000 5.7000 959.6800 ;
      RECT 0.0000 956.9600 3370.4200 958.6000 ;
      RECT 3368.7200 955.8800 3370.4200 956.9600 ;
      RECT 3305.0200 955.8800 3365.1200 956.9600 ;
      RECT 157.4200 955.8800 3302.8200 956.9600 ;
      RECT 5.3000 955.8800 155.2200 956.9600 ;
      RECT 0.0000 955.8800 1.7000 956.9600 ;
      RECT 0.0000 954.7600 3370.4200 955.8800 ;
      RECT 1.1000 954.2400 3370.4200 954.7600 ;
      RECT 1.1000 953.8600 5.7000 954.2400 ;
      RECT 3364.7200 953.1600 3370.4200 954.2400 ;
      RECT 3307.6200 953.1600 3361.1200 954.2400 ;
      RECT 154.8200 953.1600 3305.4200 954.2400 ;
      RECT 9.3000 953.1600 152.6200 954.2400 ;
      RECT 0.0000 953.1600 5.7000 953.8600 ;
      RECT 0.0000 951.5200 3370.4200 953.1600 ;
      RECT 3368.7200 950.4400 3370.4200 951.5200 ;
      RECT 3305.0200 950.4400 3365.1200 951.5200 ;
      RECT 157.4200 950.4400 3302.8200 951.5200 ;
      RECT 5.3000 950.4400 155.2200 951.5200 ;
      RECT 0.0000 950.4400 1.7000 951.5200 ;
      RECT 0.0000 948.8000 3370.4200 950.4400 ;
      RECT 3364.7200 947.7200 3370.4200 948.8000 ;
      RECT 3307.6200 947.7200 3361.1200 948.8000 ;
      RECT 154.8200 947.7200 3305.4200 948.8000 ;
      RECT 9.3000 947.7200 152.6200 948.8000 ;
      RECT 0.0000 947.7200 5.7000 948.8000 ;
      RECT 0.0000 946.0800 3370.4200 947.7200 ;
      RECT 3368.7200 945.0000 3370.4200 946.0800 ;
      RECT 3305.0200 945.0000 3365.1200 946.0800 ;
      RECT 157.4200 945.0000 3302.8200 946.0800 ;
      RECT 5.3000 945.0000 155.2200 946.0800 ;
      RECT 0.0000 945.0000 1.7000 946.0800 ;
      RECT 0.0000 944.3900 3370.4200 945.0000 ;
      RECT 1.1000 943.4900 3370.4200 944.3900 ;
      RECT 0.0000 943.3600 3370.4200 943.4900 ;
      RECT 3364.7200 942.2800 3370.4200 943.3600 ;
      RECT 3307.6200 942.2800 3361.1200 943.3600 ;
      RECT 154.8200 942.2800 3305.4200 943.3600 ;
      RECT 9.3000 942.2800 152.6200 943.3600 ;
      RECT 0.0000 942.2800 5.7000 943.3600 ;
      RECT 0.0000 940.6400 3370.4200 942.2800 ;
      RECT 3368.7200 939.5600 3370.4200 940.6400 ;
      RECT 3305.0200 939.5600 3365.1200 940.6400 ;
      RECT 157.4200 939.5600 3302.8200 940.6400 ;
      RECT 5.3000 939.5600 155.2200 940.6400 ;
      RECT 0.0000 939.5600 1.7000 940.6400 ;
      RECT 0.0000 937.9200 3370.4200 939.5600 ;
      RECT 3364.7200 936.8400 3370.4200 937.9200 ;
      RECT 3307.6200 936.8400 3361.1200 937.9200 ;
      RECT 154.8200 936.8400 3305.4200 937.9200 ;
      RECT 9.3000 936.8400 152.6200 937.9200 ;
      RECT 0.0000 936.8400 5.7000 937.9200 ;
      RECT 0.0000 935.2000 3370.4200 936.8400 ;
      RECT 3368.7200 934.1200 3370.4200 935.2000 ;
      RECT 3305.0200 934.1200 3365.1200 935.2000 ;
      RECT 157.4200 934.1200 3302.8200 935.2000 ;
      RECT 5.3000 934.1200 155.2200 935.2000 ;
      RECT 0.0000 934.1200 1.7000 935.2000 ;
      RECT 0.0000 933.4100 3370.4200 934.1200 ;
      RECT 1.1000 932.5100 3370.4200 933.4100 ;
      RECT 0.0000 932.4800 3370.4200 932.5100 ;
      RECT 3364.7200 931.4000 3370.4200 932.4800 ;
      RECT 3307.6200 931.4000 3361.1200 932.4800 ;
      RECT 154.8200 931.4000 3305.4200 932.4800 ;
      RECT 9.3000 931.4000 152.6200 932.4800 ;
      RECT 0.0000 931.4000 5.7000 932.4800 ;
      RECT 0.0000 929.7600 3370.4200 931.4000 ;
      RECT 3368.7200 928.6800 3370.4200 929.7600 ;
      RECT 3305.0200 928.6800 3365.1200 929.7600 ;
      RECT 157.4200 928.6800 3302.8200 929.7600 ;
      RECT 5.3000 928.6800 155.2200 929.7600 ;
      RECT 0.0000 928.6800 1.7000 929.7600 ;
      RECT 0.0000 927.0400 3370.4200 928.6800 ;
      RECT 3364.7200 925.9600 3370.4200 927.0400 ;
      RECT 3307.6200 925.9600 3361.1200 927.0400 ;
      RECT 154.8200 925.9600 3305.4200 927.0400 ;
      RECT 9.3000 925.9600 152.6200 927.0400 ;
      RECT 0.0000 925.9600 5.7000 927.0400 ;
      RECT 0.0000 924.3200 3370.4200 925.9600 ;
      RECT 3368.7200 923.2400 3370.4200 924.3200 ;
      RECT 3305.0200 923.2400 3365.1200 924.3200 ;
      RECT 157.4200 923.2400 3302.8200 924.3200 ;
      RECT 5.3000 923.2400 155.2200 924.3200 ;
      RECT 0.0000 923.2400 1.7000 924.3200 ;
      RECT 0.0000 922.4300 3370.4200 923.2400 ;
      RECT 1.1000 921.6000 3370.4200 922.4300 ;
      RECT 1.1000 921.5300 5.7000 921.6000 ;
      RECT 3364.7200 920.5200 3370.4200 921.6000 ;
      RECT 3307.6200 920.5200 3361.1200 921.6000 ;
      RECT 154.8200 920.5200 3305.4200 921.6000 ;
      RECT 9.3000 920.5200 152.6200 921.6000 ;
      RECT 0.0000 920.5200 5.7000 921.5300 ;
      RECT 0.0000 918.8800 3370.4200 920.5200 ;
      RECT 3368.7200 917.8000 3370.4200 918.8800 ;
      RECT 3305.0200 917.8000 3365.1200 918.8800 ;
      RECT 157.4200 917.8000 3302.8200 918.8800 ;
      RECT 5.3000 917.8000 155.2200 918.8800 ;
      RECT 0.0000 917.8000 1.7000 918.8800 ;
      RECT 0.0000 916.1600 3370.4200 917.8000 ;
      RECT 3364.7200 915.0800 3370.4200 916.1600 ;
      RECT 3307.6200 915.0800 3361.1200 916.1600 ;
      RECT 154.8200 915.0800 3305.4200 916.1600 ;
      RECT 9.3000 915.0800 152.6200 916.1600 ;
      RECT 0.0000 915.0800 5.7000 916.1600 ;
      RECT 0.0000 913.4400 3370.4200 915.0800 ;
      RECT 3368.7200 912.3600 3370.4200 913.4400 ;
      RECT 3305.0200 912.3600 3365.1200 913.4400 ;
      RECT 157.4200 912.3600 3302.8200 913.4400 ;
      RECT 5.3000 912.3600 155.2200 913.4400 ;
      RECT 0.0000 912.3600 1.7000 913.4400 ;
      RECT 0.0000 911.4500 3370.4200 912.3600 ;
      RECT 1.1000 910.7200 3370.4200 911.4500 ;
      RECT 1.1000 910.5500 5.7000 910.7200 ;
      RECT 3364.7200 909.6400 3370.4200 910.7200 ;
      RECT 3307.6200 909.6400 3361.1200 910.7200 ;
      RECT 154.8200 909.6400 3305.4200 910.7200 ;
      RECT 9.3000 909.6400 152.6200 910.7200 ;
      RECT 0.0000 909.6400 5.7000 910.5500 ;
      RECT 0.0000 908.0000 3370.4200 909.6400 ;
      RECT 3368.7200 906.9200 3370.4200 908.0000 ;
      RECT 3305.0200 906.9200 3365.1200 908.0000 ;
      RECT 157.4200 906.9200 3302.8200 908.0000 ;
      RECT 5.3000 906.9200 155.2200 908.0000 ;
      RECT 0.0000 906.9200 1.7000 908.0000 ;
      RECT 0.0000 905.2800 3370.4200 906.9200 ;
      RECT 3364.7200 904.2000 3370.4200 905.2800 ;
      RECT 3307.6200 904.2000 3361.1200 905.2800 ;
      RECT 154.8200 904.2000 3305.4200 905.2800 ;
      RECT 9.3000 904.2000 152.6200 905.2800 ;
      RECT 0.0000 904.2000 5.7000 905.2800 ;
      RECT 0.0000 902.5600 3370.4200 904.2000 ;
      RECT 3368.7200 901.4800 3370.4200 902.5600 ;
      RECT 3305.0200 901.4800 3365.1200 902.5600 ;
      RECT 157.4200 901.4800 3302.8200 902.5600 ;
      RECT 5.3000 901.4800 155.2200 902.5600 ;
      RECT 0.0000 901.4800 1.7000 902.5600 ;
      RECT 0.0000 900.4700 3370.4200 901.4800 ;
      RECT 1.1000 899.8400 3370.4200 900.4700 ;
      RECT 1.1000 899.5700 5.7000 899.8400 ;
      RECT 3364.7200 898.7600 3370.4200 899.8400 ;
      RECT 3307.6200 898.7600 3361.1200 899.8400 ;
      RECT 154.8200 898.7600 3305.4200 899.8400 ;
      RECT 9.3000 898.7600 152.6200 899.8400 ;
      RECT 0.0000 898.7600 5.7000 899.5700 ;
      RECT 0.0000 897.1200 3370.4200 898.7600 ;
      RECT 3368.7200 896.0400 3370.4200 897.1200 ;
      RECT 3305.0200 896.0400 3365.1200 897.1200 ;
      RECT 157.4200 896.0400 3302.8200 897.1200 ;
      RECT 5.3000 896.0400 155.2200 897.1200 ;
      RECT 0.0000 896.0400 1.7000 897.1200 ;
      RECT 0.0000 894.4000 3370.4200 896.0400 ;
      RECT 3364.7200 893.3200 3370.4200 894.4000 ;
      RECT 3307.6200 893.3200 3361.1200 894.4000 ;
      RECT 154.8200 893.3200 3305.4200 894.4000 ;
      RECT 9.3000 893.3200 152.6200 894.4000 ;
      RECT 0.0000 893.3200 5.7000 894.4000 ;
      RECT 0.0000 891.6800 3370.4200 893.3200 ;
      RECT 3368.7200 890.6000 3370.4200 891.6800 ;
      RECT 3305.0200 890.6000 3365.1200 891.6800 ;
      RECT 157.4200 890.6000 3302.8200 891.6800 ;
      RECT 5.3000 890.6000 155.2200 891.6800 ;
      RECT 0.0000 890.6000 1.7000 891.6800 ;
      RECT 0.0000 890.1000 3370.4200 890.6000 ;
      RECT 1.1000 889.2000 3370.4200 890.1000 ;
      RECT 0.0000 888.9600 3370.4200 889.2000 ;
      RECT 3364.7200 887.8800 3370.4200 888.9600 ;
      RECT 3307.6200 887.8800 3361.1200 888.9600 ;
      RECT 154.8200 887.8800 3305.4200 888.9600 ;
      RECT 9.3000 887.8800 152.6200 888.9600 ;
      RECT 0.0000 887.8800 5.7000 888.9600 ;
      RECT 0.0000 886.2400 3370.4200 887.8800 ;
      RECT 3368.7200 885.1600 3370.4200 886.2400 ;
      RECT 3305.0200 885.1600 3365.1200 886.2400 ;
      RECT 157.4200 885.1600 3302.8200 886.2400 ;
      RECT 5.3000 885.1600 155.2200 886.2400 ;
      RECT 0.0000 885.1600 1.7000 886.2400 ;
      RECT 0.0000 883.5200 3370.4200 885.1600 ;
      RECT 154.8200 882.7800 3305.4200 883.5200 ;
      RECT 1017.4800 882.5200 3305.4200 882.7800 ;
      RECT 3364.7200 882.4400 3370.4200 883.5200 ;
      RECT 3307.6200 882.4400 3361.1200 883.5200 ;
      RECT 2436.3200 882.4400 3305.4200 882.5200 ;
      RECT 154.8200 882.4400 1015.2800 882.7800 ;
      RECT 9.3000 882.4400 152.6200 883.5200 ;
      RECT 0.0000 882.4400 5.7000 883.5200 ;
      RECT 1017.4800 881.7000 1295.6000 882.5200 ;
      RECT 0.0000 881.7000 1015.2800 882.4400 ;
      RECT 2436.3200 881.4400 3370.4200 882.4400 ;
      RECT 2178.6800 881.4400 2434.1200 882.5200 ;
      RECT 1738.2400 881.4400 2176.4800 882.5200 ;
      RECT 1518.0200 881.4400 1736.0400 882.5200 ;
      RECT 1297.8000 881.4400 1515.8200 882.5200 ;
      RECT 0.0000 881.4400 1295.6000 881.7000 ;
      RECT 0.0000 880.8000 3370.4200 881.4400 ;
      RECT 3368.7200 879.7200 3370.4200 880.8000 ;
      RECT 3305.0200 879.7200 3365.1200 880.8000 ;
      RECT 157.4200 879.7200 3302.8200 880.8000 ;
      RECT 5.3000 879.7200 155.2200 880.8000 ;
      RECT 0.0000 879.7200 1.7000 880.8000 ;
      RECT 0.0000 879.6100 3370.4200 879.7200 ;
      RECT 1065.1600 879.4500 3370.4200 879.6100 ;
      RECT 0.0000 879.1200 1005.2200 879.6100 ;
      RECT 1.1000 878.2200 1005.2200 879.1200 ;
      RECT 2446.4800 878.0800 3370.4200 879.4500 ;
      RECT 0.0000 878.0800 1005.2200 878.2200 ;
      RECT 1065.1600 877.4100 1283.0400 879.4500 ;
      RECT 1011.2200 877.4100 1059.1600 879.6100 ;
      RECT 154.8200 877.4100 1005.2200 878.0800 ;
      RECT 2446.4800 877.2500 3305.4200 878.0800 ;
      RECT 2392.5400 877.2500 2440.4800 879.4500 ;
      RECT 2172.3200 877.2500 2380.3400 879.4500 ;
      RECT 1945.9000 877.2500 2163.9200 879.4500 ;
      RECT 1731.8800 877.2500 1939.9000 879.4500 ;
      RECT 1511.6600 877.2500 1719.6800 879.4500 ;
      RECT 1291.4400 877.2500 1499.4600 879.4500 ;
      RECT 154.8200 877.2500 1283.0400 877.4100 ;
      RECT 154.8200 877.2100 3305.4200 877.2500 ;
      RECT 3364.7200 877.0000 3370.4200 878.0800 ;
      RECT 3307.6200 877.0000 3361.1200 878.0800 ;
      RECT 1067.7600 877.0000 3305.4200 877.2100 ;
      RECT 154.8200 877.0000 1002.6200 877.2100 ;
      RECT 9.3000 877.0000 152.6200 878.0800 ;
      RECT 0.0000 877.0000 5.7000 878.0800 ;
      RECT 1067.7600 876.8500 3370.4200 877.0000 ;
      RECT 2449.0800 875.3600 3370.4200 876.8500 ;
      RECT 0.0000 875.3600 1002.6200 877.0000 ;
      RECT 1067.7600 875.0100 1285.6400 876.8500 ;
      RECT 1011.2200 875.0100 1059.1600 877.2100 ;
      RECT 157.4200 875.0100 1002.6200 875.3600 ;
      RECT 2449.0800 874.6500 3302.8200 875.3600 ;
      RECT 2392.5400 874.6500 2440.4800 876.8500 ;
      RECT 2172.3200 874.6500 2380.3400 876.8500 ;
      RECT 1948.5000 874.6500 2166.5200 876.8500 ;
      RECT 1731.8800 874.6500 1939.9000 876.8500 ;
      RECT 1511.6600 874.6500 1719.6800 876.8500 ;
      RECT 1291.4400 874.6500 1499.4600 876.8500 ;
      RECT 157.4200 874.6500 1285.6400 875.0100 ;
      RECT 3368.7200 874.2800 3370.4200 875.3600 ;
      RECT 3305.0200 874.2800 3365.1200 875.3600 ;
      RECT 157.4200 874.2800 3302.8200 874.6500 ;
      RECT 5.3000 874.2800 155.2200 875.3600 ;
      RECT 0.0000 874.2800 1.7000 875.3600 ;
      RECT 0.0000 872.6400 3370.4200 874.2800 ;
      RECT 3364.7200 871.5600 3370.4200 872.6400 ;
      RECT 3307.6200 871.5600 3361.1200 872.6400 ;
      RECT 154.8200 871.5600 3305.4200 872.6400 ;
      RECT 9.3000 871.5600 152.6200 872.6400 ;
      RECT 0.0000 871.5600 5.7000 872.6400 ;
      RECT 0.0000 869.9200 3370.4200 871.5600 ;
      RECT 157.4200 869.6800 3302.8200 869.9200 ;
      RECT 5.3000 869.6800 155.2200 869.9200 ;
      RECT 1065.1600 869.4200 3302.8200 869.6800 ;
      RECT 3368.7200 868.8400 3370.4200 869.9200 ;
      RECT 3305.0200 868.8400 3365.1200 869.9200 ;
      RECT 2446.4800 868.8400 3302.8200 869.4200 ;
      RECT 0.0000 868.1400 1.7000 869.9200 ;
      RECT 1065.1600 867.4800 1283.0400 869.4200 ;
      RECT 167.4150 867.4800 953.1450 869.6800 ;
      RECT 1.1000 867.4800 1.7000 868.1400 ;
      RECT 1.1000 867.2400 1283.0400 867.4800 ;
      RECT 2446.4800 867.2200 3370.4200 868.8400 ;
      RECT 1945.9000 867.2200 2163.9200 869.4200 ;
      RECT 0.0000 867.2200 1283.0400 867.2400 ;
      RECT 0.0000 867.2000 3370.4200 867.2200 ;
      RECT 154.8200 867.0800 3305.4200 867.2000 ;
      RECT 9.3000 867.0800 152.6200 867.2000 ;
      RECT 1067.7600 866.8200 3305.4200 867.0800 ;
      RECT 3364.7200 866.1200 3370.4200 867.2000 ;
      RECT 3307.6200 866.1200 3361.1200 867.2000 ;
      RECT 2449.0800 866.1200 3305.4200 866.8200 ;
      RECT 1067.7600 864.8800 1285.6400 866.8200 ;
      RECT 167.4150 864.8800 953.1450 867.0800 ;
      RECT 0.0000 864.8800 5.7000 867.2000 ;
      RECT 2449.0800 864.6200 3370.4200 866.1200 ;
      RECT 1948.5000 864.6200 2166.5200 866.8200 ;
      RECT 0.0000 864.6200 1285.6400 864.8800 ;
      RECT 0.0000 864.4800 3370.4200 864.6200 ;
      RECT 3368.7200 863.4000 3370.4200 864.4800 ;
      RECT 3305.0200 863.4000 3365.1200 864.4800 ;
      RECT 157.4200 863.4000 3302.8200 864.4800 ;
      RECT 5.3000 863.4000 155.2200 864.4800 ;
      RECT 0.0000 863.4000 1.7000 864.4800 ;
      RECT 0.0000 861.7600 3370.4200 863.4000 ;
      RECT 3364.7200 860.6800 3370.4200 861.7600 ;
      RECT 3307.6200 860.6800 3361.1200 861.7600 ;
      RECT 154.8200 860.6800 3305.4200 861.7600 ;
      RECT 9.3000 860.6800 152.6200 861.7600 ;
      RECT 0.0000 860.6800 5.7000 861.7600 ;
      RECT 0.0000 859.0700 3370.4200 860.6800 ;
      RECT 1067.7600 859.0400 3370.4200 859.0700 ;
      RECT 0.0000 859.0400 1002.6200 859.0700 ;
      RECT 1067.7600 858.9100 3302.8200 859.0400 ;
      RECT 3368.7200 857.9600 3370.4200 859.0400 ;
      RECT 3305.0200 857.9600 3365.1200 859.0400 ;
      RECT 2449.0800 857.9600 3302.8200 858.9100 ;
      RECT 157.4200 857.9600 1002.6200 859.0400 ;
      RECT 5.3000 857.9600 155.2200 859.0400 ;
      RECT 0.0000 857.9600 1.7000 859.0400 ;
      RECT 0.0000 857.1600 1002.6200 857.9600 ;
      RECT 1067.7600 856.8700 1285.6400 858.9100 ;
      RECT 1011.2200 856.8700 1059.1600 859.0700 ;
      RECT 1.1000 856.8700 1002.6200 857.1600 ;
      RECT 2449.0800 856.7100 3370.4200 857.9600 ;
      RECT 2392.5400 856.7100 2440.4800 858.9100 ;
      RECT 2172.3200 856.7100 2380.3400 858.9100 ;
      RECT 1948.5000 856.7100 2166.5200 858.9100 ;
      RECT 1731.8800 856.7100 1939.9000 858.9100 ;
      RECT 1511.6600 856.7100 1719.6800 858.9100 ;
      RECT 1291.4400 856.7100 1499.4600 858.9100 ;
      RECT 1.1000 856.7100 1285.6400 856.8700 ;
      RECT 1.1000 856.6700 3370.4200 856.7100 ;
      RECT 1065.1600 856.3200 3370.4200 856.6700 ;
      RECT 1.1000 856.3200 1005.2200 856.6700 ;
      RECT 1065.1600 856.3100 3305.4200 856.3200 ;
      RECT 1.1000 856.2600 5.7000 856.3200 ;
      RECT 3364.7200 855.2400 3370.4200 856.3200 ;
      RECT 3307.6200 855.2400 3361.1200 856.3200 ;
      RECT 2446.4800 855.2400 3305.4200 856.3100 ;
      RECT 154.8200 855.2400 1005.2200 856.3200 ;
      RECT 9.3000 855.2400 152.6200 856.3200 ;
      RECT 0.0000 855.2400 5.7000 856.2600 ;
      RECT 1065.1600 854.4700 1283.0400 856.3100 ;
      RECT 1011.2200 854.4700 1059.1600 856.6700 ;
      RECT 0.0000 854.4700 1005.2200 855.2400 ;
      RECT 2446.4800 854.1100 3370.4200 855.2400 ;
      RECT 2392.5400 854.1100 2440.4800 856.3100 ;
      RECT 2172.3200 854.1100 2380.3400 856.3100 ;
      RECT 1945.9000 854.1100 2163.9200 856.3100 ;
      RECT 1731.8800 854.1100 1939.9000 856.3100 ;
      RECT 1511.6600 854.1100 1719.6800 856.3100 ;
      RECT 1291.4400 854.1100 1499.4600 856.3100 ;
      RECT 0.0000 854.1100 1283.0400 854.4700 ;
      RECT 0.0000 853.6000 3370.4200 854.1100 ;
      RECT 3368.7200 852.5200 3370.4200 853.6000 ;
      RECT 3305.0200 852.5200 3365.1200 853.6000 ;
      RECT 157.4200 852.5200 3302.8200 853.6000 ;
      RECT 5.3000 852.5200 155.2200 853.6000 ;
      RECT 0.0000 852.5200 1.7000 853.6000 ;
      RECT 0.0000 851.7000 3370.4200 852.5200 ;
      RECT 1015.0800 851.4400 3370.4200 851.7000 ;
      RECT 2396.3000 850.8800 3370.4200 851.4400 ;
      RECT 0.0000 850.8800 1012.8800 851.7000 ;
      RECT 1015.0800 850.6200 1293.0000 851.4400 ;
      RECT 154.8200 850.6200 1012.8800 850.8800 ;
      RECT 2396.3000 850.3600 3305.4200 850.8800 ;
      RECT 2176.0800 850.3600 2394.1000 851.4400 ;
      RECT 1735.6400 850.3600 2173.8800 851.4400 ;
      RECT 1515.4200 850.3600 1733.4400 851.4400 ;
      RECT 1295.2000 850.3600 1513.2200 851.4400 ;
      RECT 154.8200 850.3600 1293.0000 850.6200 ;
      RECT 3364.7200 849.8000 3370.4200 850.8800 ;
      RECT 3307.6200 849.8000 3361.1200 850.8800 ;
      RECT 154.8200 849.8000 3305.4200 850.3600 ;
      RECT 9.3000 849.8000 152.6200 850.8800 ;
      RECT 0.0000 849.8000 5.7000 850.8800 ;
      RECT 0.0000 848.1600 3370.4200 849.8000 ;
      RECT 3368.7200 847.0800 3370.4200 848.1600 ;
      RECT 3305.0200 847.0800 3365.1200 848.1600 ;
      RECT 157.4200 847.0800 3302.8200 848.1600 ;
      RECT 5.3000 847.0800 155.2200 848.1600 ;
      RECT 0.0000 847.0800 1.7000 848.1600 ;
      RECT 0.0000 846.1800 3370.4200 847.0800 ;
      RECT 1.1000 845.4400 3370.4200 846.1800 ;
      RECT 1.1000 845.2800 5.7000 845.4400 ;
      RECT 3364.7200 844.3600 3370.4200 845.4400 ;
      RECT 3307.6200 844.3600 3361.1200 845.4400 ;
      RECT 154.8200 844.3600 3305.4200 845.4400 ;
      RECT 9.3000 844.3600 152.6200 845.4400 ;
      RECT 0.0000 844.3600 5.7000 845.2800 ;
      RECT 0.0000 842.7200 3370.4200 844.3600 ;
      RECT 3368.7200 841.6400 3370.4200 842.7200 ;
      RECT 3305.0200 841.6400 3365.1200 842.7200 ;
      RECT 157.4200 841.6400 3302.8200 842.7200 ;
      RECT 5.3000 841.6400 155.2200 842.7200 ;
      RECT 0.0000 841.6400 1.7000 842.7200 ;
      RECT 0.0000 840.0000 3370.4200 841.6400 ;
      RECT 3364.7200 838.9200 3370.4200 840.0000 ;
      RECT 3307.6200 838.9200 3361.1200 840.0000 ;
      RECT 154.8200 838.9200 3305.4200 840.0000 ;
      RECT 9.3000 838.9200 152.6200 840.0000 ;
      RECT 0.0000 838.9200 5.7000 840.0000 ;
      RECT 0.0000 837.2800 3370.4200 838.9200 ;
      RECT 3368.7200 836.2000 3370.4200 837.2800 ;
      RECT 3305.0200 836.2000 3365.1200 837.2800 ;
      RECT 157.4200 836.2000 3302.8200 837.2800 ;
      RECT 5.3000 836.2000 155.2200 837.2800 ;
      RECT 0.0000 836.2000 1.7000 837.2800 ;
      RECT 0.0000 835.8100 3370.4200 836.2000 ;
      RECT 1.1000 834.9100 3370.4200 835.8100 ;
      RECT 0.0000 834.5600 3370.4200 834.9100 ;
      RECT 3364.7200 833.4800 3370.4200 834.5600 ;
      RECT 3307.6200 833.4800 3361.1200 834.5600 ;
      RECT 154.8200 833.4800 3305.4200 834.5600 ;
      RECT 9.3000 833.4800 152.6200 834.5600 ;
      RECT 0.0000 833.4800 5.7000 834.5600 ;
      RECT 0.0000 831.8400 3370.4200 833.4800 ;
      RECT 3368.7200 830.7600 3370.4200 831.8400 ;
      RECT 3305.0200 830.7600 3365.1200 831.8400 ;
      RECT 157.4200 830.7600 3302.8200 831.8400 ;
      RECT 5.3000 830.7600 155.2200 831.8400 ;
      RECT 0.0000 830.7600 1.7000 831.8400 ;
      RECT 0.0000 829.1200 3370.4200 830.7600 ;
      RECT 3364.7200 828.0400 3370.4200 829.1200 ;
      RECT 3307.6200 828.0400 3361.1200 829.1200 ;
      RECT 154.8200 828.0400 3305.4200 829.1200 ;
      RECT 9.3000 828.0400 152.6200 829.1200 ;
      RECT 0.0000 828.0400 5.7000 829.1200 ;
      RECT 0.0000 826.4000 3370.4200 828.0400 ;
      RECT 3368.7200 825.3200 3370.4200 826.4000 ;
      RECT 3305.0200 825.3200 3365.1200 826.4000 ;
      RECT 157.4200 825.3200 3302.8200 826.4000 ;
      RECT 5.3000 825.3200 155.2200 826.4000 ;
      RECT 0.0000 825.3200 1.7000 826.4000 ;
      RECT 0.0000 824.8300 3370.4200 825.3200 ;
      RECT 1.1000 823.9300 3370.4200 824.8300 ;
      RECT 0.0000 823.6800 3370.4200 823.9300 ;
      RECT 3364.7200 822.6000 3370.4200 823.6800 ;
      RECT 3307.6200 822.6000 3361.1200 823.6800 ;
      RECT 154.8200 822.6000 3305.4200 823.6800 ;
      RECT 9.3000 822.6000 152.6200 823.6800 ;
      RECT 0.0000 822.6000 5.7000 823.6800 ;
      RECT 0.0000 820.9600 3370.4200 822.6000 ;
      RECT 3368.7200 819.8800 3370.4200 820.9600 ;
      RECT 3305.0200 819.8800 3365.1200 820.9600 ;
      RECT 157.4200 819.8800 3302.8200 820.9600 ;
      RECT 5.3000 819.8800 155.2200 820.9600 ;
      RECT 0.0000 819.8800 1.7000 820.9600 ;
      RECT 0.0000 818.2400 3370.4200 819.8800 ;
      RECT 3364.7200 817.1600 3370.4200 818.2400 ;
      RECT 3307.6200 817.1600 3361.1200 818.2400 ;
      RECT 154.8200 817.1600 3305.4200 818.2400 ;
      RECT 9.3000 817.1600 152.6200 818.2400 ;
      RECT 0.0000 817.1600 5.7000 818.2400 ;
      RECT 0.0000 815.5200 3370.4200 817.1600 ;
      RECT 3368.7200 814.4400 3370.4200 815.5200 ;
      RECT 3305.0200 814.4400 3365.1200 815.5200 ;
      RECT 157.4200 814.4400 3302.8200 815.5200 ;
      RECT 5.3000 814.4400 155.2200 815.5200 ;
      RECT 0.0000 814.4400 1.7000 815.5200 ;
      RECT 0.0000 813.8500 3370.4200 814.4400 ;
      RECT 1.1000 812.9500 3370.4200 813.8500 ;
      RECT 0.0000 812.8000 3370.4200 812.9500 ;
      RECT 3364.7200 811.7200 3370.4200 812.8000 ;
      RECT 3307.6200 811.7200 3361.1200 812.8000 ;
      RECT 154.8200 811.7200 3305.4200 812.8000 ;
      RECT 9.3000 811.7200 152.6200 812.8000 ;
      RECT 0.0000 811.7200 5.7000 812.8000 ;
      RECT 0.0000 810.0800 3370.4200 811.7200 ;
      RECT 3368.7200 809.0000 3370.4200 810.0800 ;
      RECT 3305.0200 809.0000 3365.1200 810.0800 ;
      RECT 157.4200 809.0000 3302.8200 810.0800 ;
      RECT 5.3000 809.0000 155.2200 810.0800 ;
      RECT 0.0000 809.0000 1.7000 810.0800 ;
      RECT 0.0000 807.3600 3370.4200 809.0000 ;
      RECT 3364.7200 806.2800 3370.4200 807.3600 ;
      RECT 3307.6200 806.2800 3361.1200 807.3600 ;
      RECT 154.8200 806.2800 3305.4200 807.3600 ;
      RECT 9.3000 806.2800 152.6200 807.3600 ;
      RECT 0.0000 806.2800 5.7000 807.3600 ;
      RECT 0.0000 804.6400 3370.4200 806.2800 ;
      RECT 3368.7200 803.5600 3370.4200 804.6400 ;
      RECT 3305.0200 803.5600 3365.1200 804.6400 ;
      RECT 157.4200 803.5600 3302.8200 804.6400 ;
      RECT 5.3000 803.5600 155.2200 804.6400 ;
      RECT 0.0000 803.5600 1.7000 804.6400 ;
      RECT 0.0000 802.8700 3370.4200 803.5600 ;
      RECT 1.1000 801.9700 3370.4200 802.8700 ;
      RECT 0.0000 801.9200 3370.4200 801.9700 ;
      RECT 3364.7200 800.8400 3370.4200 801.9200 ;
      RECT 3307.6200 800.8400 3361.1200 801.9200 ;
      RECT 154.8200 800.8400 3305.4200 801.9200 ;
      RECT 9.3000 800.8400 152.6200 801.9200 ;
      RECT 0.0000 800.8400 5.7000 801.9200 ;
      RECT 0.0000 799.2000 3370.4200 800.8400 ;
      RECT 3368.7200 798.1200 3370.4200 799.2000 ;
      RECT 3305.0200 798.1200 3365.1200 799.2000 ;
      RECT 157.4200 798.1200 3302.8200 799.2000 ;
      RECT 5.3000 798.1200 155.2200 799.2000 ;
      RECT 0.0000 798.1200 1.7000 799.2000 ;
      RECT 0.0000 796.4800 3370.4200 798.1200 ;
      RECT 3364.7200 795.4000 3370.4200 796.4800 ;
      RECT 3307.6200 795.4000 3361.1200 796.4800 ;
      RECT 154.8200 795.4000 3305.4200 796.4800 ;
      RECT 9.3000 795.4000 152.6200 796.4800 ;
      RECT 0.0000 795.4000 5.7000 796.4800 ;
      RECT 0.0000 793.7600 3370.4200 795.4000 ;
      RECT 3368.7200 792.6800 3370.4200 793.7600 ;
      RECT 3305.0200 792.6800 3365.1200 793.7600 ;
      RECT 157.4200 792.6800 3302.8200 793.7600 ;
      RECT 5.3000 792.6800 155.2200 793.7600 ;
      RECT 0.0000 792.6800 1.7000 793.7600 ;
      RECT 0.0000 791.8900 3370.4200 792.6800 ;
      RECT 1.1000 791.0400 3370.4200 791.8900 ;
      RECT 1.1000 790.9900 5.7000 791.0400 ;
      RECT 3364.7200 789.9600 3370.4200 791.0400 ;
      RECT 3307.6200 789.9600 3361.1200 791.0400 ;
      RECT 154.8200 789.9600 3305.4200 791.0400 ;
      RECT 9.3000 789.9600 152.6200 791.0400 ;
      RECT 0.0000 789.9600 5.7000 790.9900 ;
      RECT 0.0000 788.3200 3370.4200 789.9600 ;
      RECT 3368.7200 787.2400 3370.4200 788.3200 ;
      RECT 3305.0200 787.2400 3365.1200 788.3200 ;
      RECT 157.4200 787.2400 3302.8200 788.3200 ;
      RECT 5.3000 787.2400 155.2200 788.3200 ;
      RECT 0.0000 787.2400 1.7000 788.3200 ;
      RECT 0.0000 785.6000 3370.4200 787.2400 ;
      RECT 3364.7200 784.5200 3370.4200 785.6000 ;
      RECT 3307.6200 784.5200 3361.1200 785.6000 ;
      RECT 154.8200 784.5200 3305.4200 785.6000 ;
      RECT 9.3000 784.5200 152.6200 785.6000 ;
      RECT 0.0000 784.5200 5.7000 785.6000 ;
      RECT 0.0000 782.8800 3370.4200 784.5200 ;
      RECT 3368.7200 781.8000 3370.4200 782.8800 ;
      RECT 3305.0200 781.8000 3365.1200 782.8800 ;
      RECT 157.4200 781.8000 3302.8200 782.8800 ;
      RECT 5.3000 781.8000 155.2200 782.8800 ;
      RECT 0.0000 781.8000 1.7000 782.8800 ;
      RECT 0.0000 781.5200 3370.4200 781.8000 ;
      RECT 1.1000 780.6200 3370.4200 781.5200 ;
      RECT 0.0000 780.1600 3370.4200 780.6200 ;
      RECT 3364.7200 779.0800 3370.4200 780.1600 ;
      RECT 3307.6200 779.0800 3361.1200 780.1600 ;
      RECT 154.8200 779.0800 3305.4200 780.1600 ;
      RECT 9.3000 779.0800 152.6200 780.1600 ;
      RECT 0.0000 779.0800 5.7000 780.1600 ;
      RECT 0.0000 777.4400 3370.4200 779.0800 ;
      RECT 3368.7200 776.3600 3370.4200 777.4400 ;
      RECT 3305.0200 776.3600 3365.1200 777.4400 ;
      RECT 157.4200 776.3600 3302.8200 777.4400 ;
      RECT 5.3000 776.3600 155.2200 777.4400 ;
      RECT 0.0000 776.3600 1.7000 777.4400 ;
      RECT 0.0000 774.7200 3370.4200 776.3600 ;
      RECT 3364.7200 773.6400 3370.4200 774.7200 ;
      RECT 3307.6200 773.6400 3361.1200 774.7200 ;
      RECT 154.8200 773.6400 3305.4200 774.7200 ;
      RECT 9.3000 773.6400 152.6200 774.7200 ;
      RECT 0.0000 773.6400 5.7000 774.7200 ;
      RECT 0.0000 772.0000 3370.4200 773.6400 ;
      RECT 3368.7200 770.9200 3370.4200 772.0000 ;
      RECT 3305.0200 770.9200 3365.1200 772.0000 ;
      RECT 157.4200 770.9200 3302.8200 772.0000 ;
      RECT 5.3000 770.9200 155.2200 772.0000 ;
      RECT 0.0000 770.9200 1.7000 772.0000 ;
      RECT 0.0000 770.5400 3370.4200 770.9200 ;
      RECT 1.1000 769.6400 3370.4200 770.5400 ;
      RECT 0.0000 769.2800 3370.4200 769.6400 ;
      RECT 3364.7200 768.2000 3370.4200 769.2800 ;
      RECT 3307.6200 768.2000 3361.1200 769.2800 ;
      RECT 154.8200 768.2000 3305.4200 769.2800 ;
      RECT 9.3000 768.2000 152.6200 769.2800 ;
      RECT 0.0000 768.2000 5.7000 769.2800 ;
      RECT 0.0000 766.5600 3370.4200 768.2000 ;
      RECT 3368.7200 765.4800 3370.4200 766.5600 ;
      RECT 3305.0200 765.4800 3365.1200 766.5600 ;
      RECT 157.4200 765.4800 3302.8200 766.5600 ;
      RECT 5.3000 765.4800 155.2200 766.5600 ;
      RECT 0.0000 765.4800 1.7000 766.5600 ;
      RECT 0.0000 763.8400 3370.4200 765.4800 ;
      RECT 3364.7200 762.7600 3370.4200 763.8400 ;
      RECT 3307.6200 762.7600 3361.1200 763.8400 ;
      RECT 154.8200 762.7600 3305.4200 763.8400 ;
      RECT 9.3000 762.7600 152.6200 763.8400 ;
      RECT 0.0000 762.7600 5.7000 763.8400 ;
      RECT 0.0000 761.1200 3370.4200 762.7600 ;
      RECT 3368.7200 760.0400 3370.4200 761.1200 ;
      RECT 3305.0200 760.0400 3365.1200 761.1200 ;
      RECT 157.4200 760.0400 3302.8200 761.1200 ;
      RECT 5.3000 760.0400 155.2200 761.1200 ;
      RECT 0.0000 760.0400 1.7000 761.1200 ;
      RECT 0.0000 759.5600 3370.4200 760.0400 ;
      RECT 1.1000 758.6600 3370.4200 759.5600 ;
      RECT 0.0000 758.4000 3370.4200 758.6600 ;
      RECT 3364.7200 757.3200 3370.4200 758.4000 ;
      RECT 3307.6200 757.3200 3361.1200 758.4000 ;
      RECT 154.8200 757.3200 3305.4200 758.4000 ;
      RECT 9.3000 757.3200 152.6200 758.4000 ;
      RECT 0.0000 757.3200 5.7000 758.4000 ;
      RECT 0.0000 755.6800 3370.4200 757.3200 ;
      RECT 3368.7200 754.6000 3370.4200 755.6800 ;
      RECT 3305.0200 754.6000 3365.1200 755.6800 ;
      RECT 157.4200 754.6000 3302.8200 755.6800 ;
      RECT 5.3000 754.6000 155.2200 755.6800 ;
      RECT 0.0000 754.6000 1.7000 755.6800 ;
      RECT 0.0000 752.9600 3370.4200 754.6000 ;
      RECT 3364.7200 751.8800 3370.4200 752.9600 ;
      RECT 3307.6200 751.8800 3361.1200 752.9600 ;
      RECT 154.8200 751.8800 3305.4200 752.9600 ;
      RECT 9.3000 751.8800 152.6200 752.9600 ;
      RECT 0.0000 751.8800 5.7000 752.9600 ;
      RECT 0.0000 750.2400 3370.4200 751.8800 ;
      RECT 3368.7200 749.1600 3370.4200 750.2400 ;
      RECT 3305.0200 749.1600 3365.1200 750.2400 ;
      RECT 2497.4200 749.1600 3302.8200 750.2400 ;
      RECT 2446.4800 749.1600 2495.2200 750.2400 ;
      RECT 1007.4200 749.1600 2444.2800 750.2400 ;
      RECT 965.0200 749.1600 1005.2200 750.2400 ;
      RECT 157.4200 749.1600 962.8200 750.2400 ;
      RECT 5.3000 749.1600 155.2200 750.2400 ;
      RECT 0.0000 749.1600 1.7000 750.2400 ;
      RECT 0.0000 748.5800 3370.4200 749.1600 ;
      RECT 1.1000 747.6800 3370.4200 748.5800 ;
      RECT 0.0000 747.5200 3370.4200 747.6800 ;
      RECT 3364.7200 746.4400 3370.4200 747.5200 ;
      RECT 3307.6200 746.4400 3361.1200 747.5200 ;
      RECT 2494.8200 746.4400 3305.4200 747.5200 ;
      RECT 2449.0800 746.4400 2492.6200 747.5200 ;
      RECT 1004.8200 746.4400 2446.8800 747.5200 ;
      RECT 967.6200 746.4400 1002.6200 747.5200 ;
      RECT 154.8200 746.4400 965.4200 747.5200 ;
      RECT 9.3000 746.4400 152.6200 747.5200 ;
      RECT 0.0000 746.4400 5.7000 747.5200 ;
      RECT 0.0000 744.8000 3370.4200 746.4400 ;
      RECT 3368.7200 743.7200 3370.4200 744.8000 ;
      RECT 3305.0200 743.7200 3365.1200 744.8000 ;
      RECT 2497.4200 743.7200 3302.8200 744.8000 ;
      RECT 2446.4800 743.7200 2495.2200 744.8000 ;
      RECT 1007.4200 743.7200 2444.2800 744.8000 ;
      RECT 965.0200 743.7200 1005.2200 744.8000 ;
      RECT 157.4200 743.7200 962.8200 744.8000 ;
      RECT 5.3000 743.7200 155.2200 744.8000 ;
      RECT 0.0000 743.7200 1.7000 744.8000 ;
      RECT 0.0000 742.0800 3370.4200 743.7200 ;
      RECT 3364.7200 741.0000 3370.4200 742.0800 ;
      RECT 3307.6200 741.0000 3361.1200 742.0800 ;
      RECT 2494.8200 741.0000 3305.4200 742.0800 ;
      RECT 2449.0800 741.0000 2492.6200 742.0800 ;
      RECT 1004.8200 741.0000 2446.8800 742.0800 ;
      RECT 967.6200 741.0000 1002.6200 742.0800 ;
      RECT 154.8200 741.0000 965.4200 742.0800 ;
      RECT 9.3000 741.0000 152.6200 742.0800 ;
      RECT 0.0000 741.0000 5.7000 742.0800 ;
      RECT 0.0000 739.3600 3370.4200 741.0000 ;
      RECT 3368.7200 738.2800 3370.4200 739.3600 ;
      RECT 3305.0200 738.2800 3365.1200 739.3600 ;
      RECT 2497.4200 738.2800 3302.8200 739.3600 ;
      RECT 2446.4800 738.2800 2495.2200 739.3600 ;
      RECT 1007.4200 738.2800 2444.2800 739.3600 ;
      RECT 965.0200 738.2800 1005.2200 739.3600 ;
      RECT 157.4200 738.2800 962.8200 739.3600 ;
      RECT 5.3000 738.2800 155.2200 739.3600 ;
      RECT 0.0000 738.2800 1.7000 739.3600 ;
      RECT 0.0000 737.6000 3370.4200 738.2800 ;
      RECT 1.1000 736.7000 3370.4200 737.6000 ;
      RECT 0.0000 736.6400 3370.4200 736.7000 ;
      RECT 3364.7200 735.5600 3370.4200 736.6400 ;
      RECT 3307.6200 735.5600 3361.1200 736.6400 ;
      RECT 2494.8200 735.5600 3305.4200 736.6400 ;
      RECT 2449.0800 735.5600 2492.6200 736.6400 ;
      RECT 1004.8200 735.5600 2446.8800 736.6400 ;
      RECT 967.6200 735.5600 1002.6200 736.6400 ;
      RECT 154.8200 735.5600 965.4200 736.6400 ;
      RECT 9.3000 735.5600 152.6200 736.6400 ;
      RECT 0.0000 735.5600 5.7000 736.6400 ;
      RECT 0.0000 733.9200 3370.4200 735.5600 ;
      RECT 3368.7200 732.8400 3370.4200 733.9200 ;
      RECT 3305.0200 732.8400 3365.1200 733.9200 ;
      RECT 2497.4200 732.8400 3302.8200 733.9200 ;
      RECT 2446.4800 732.8400 2495.2200 733.9200 ;
      RECT 1007.4200 732.8400 2444.2800 733.9200 ;
      RECT 965.0200 732.8400 1005.2200 733.9200 ;
      RECT 157.4200 732.8400 962.8200 733.9200 ;
      RECT 5.3000 732.8400 155.2200 733.9200 ;
      RECT 0.0000 732.8400 1.7000 733.9200 ;
      RECT 0.0000 731.2000 3370.4200 732.8400 ;
      RECT 3364.7200 730.1200 3370.4200 731.2000 ;
      RECT 3307.6200 730.1200 3361.1200 731.2000 ;
      RECT 2494.8200 730.1200 3305.4200 731.2000 ;
      RECT 2449.0800 730.1200 2492.6200 731.2000 ;
      RECT 1004.8200 730.1200 2446.8800 731.2000 ;
      RECT 967.6200 730.1200 1002.6200 731.2000 ;
      RECT 154.8200 730.1200 965.4200 731.2000 ;
      RECT 9.3000 730.1200 152.6200 731.2000 ;
      RECT 0.0000 730.1200 5.7000 731.2000 ;
      RECT 0.0000 728.4800 3370.4200 730.1200 ;
      RECT 3368.7200 727.4000 3370.4200 728.4800 ;
      RECT 3305.0200 727.4000 3365.1200 728.4800 ;
      RECT 2497.4200 727.4000 3302.8200 728.4800 ;
      RECT 2446.4800 727.4000 2495.2200 728.4800 ;
      RECT 1007.4200 727.4000 2444.2800 728.4800 ;
      RECT 965.0200 727.4000 1005.2200 728.4800 ;
      RECT 157.4200 727.4000 962.8200 728.4800 ;
      RECT 5.3000 727.4000 155.2200 728.4800 ;
      RECT 0.0000 727.4000 1.7000 728.4800 ;
      RECT 0.0000 727.2300 3370.4200 727.4000 ;
      RECT 1.1000 726.3300 3370.4200 727.2300 ;
      RECT 0.0000 725.7600 3370.4200 726.3300 ;
      RECT 3364.7200 724.6800 3370.4200 725.7600 ;
      RECT 3307.6200 724.6800 3361.1200 725.7600 ;
      RECT 2494.8200 724.6800 3305.4200 725.7600 ;
      RECT 2449.0800 724.6800 2492.6200 725.7600 ;
      RECT 1004.8200 724.6800 2446.8800 725.7600 ;
      RECT 967.6200 724.6800 1002.6200 725.7600 ;
      RECT 154.8200 724.6800 965.4200 725.7600 ;
      RECT 9.3000 724.6800 152.6200 725.7600 ;
      RECT 0.0000 724.6800 5.7000 725.7600 ;
      RECT 0.0000 723.0400 3370.4200 724.6800 ;
      RECT 3368.7200 721.9600 3370.4200 723.0400 ;
      RECT 3305.0200 721.9600 3365.1200 723.0400 ;
      RECT 2497.4200 721.9600 3302.8200 723.0400 ;
      RECT 2446.4800 721.9600 2495.2200 723.0400 ;
      RECT 1007.4200 721.9600 2444.2800 723.0400 ;
      RECT 965.0200 721.9600 1005.2200 723.0400 ;
      RECT 157.4200 721.9600 962.8200 723.0400 ;
      RECT 5.3000 721.9600 155.2200 723.0400 ;
      RECT 0.0000 721.9600 1.7000 723.0400 ;
      RECT 0.0000 720.3200 3370.4200 721.9600 ;
      RECT 3364.7200 719.2400 3370.4200 720.3200 ;
      RECT 3307.6200 719.2400 3361.1200 720.3200 ;
      RECT 2494.8200 719.2400 3305.4200 720.3200 ;
      RECT 2449.0800 719.2400 2492.6200 720.3200 ;
      RECT 1004.8200 719.2400 2446.8800 720.3200 ;
      RECT 967.6200 719.2400 1002.6200 720.3200 ;
      RECT 154.8200 719.2400 965.4200 720.3200 ;
      RECT 9.3000 719.2400 152.6200 720.3200 ;
      RECT 0.0000 719.2400 5.7000 720.3200 ;
      RECT 0.0000 717.6000 3370.4200 719.2400 ;
      RECT 3368.7200 716.5200 3370.4200 717.6000 ;
      RECT 3305.0200 716.5200 3365.1200 717.6000 ;
      RECT 2497.4200 716.5200 3302.8200 717.6000 ;
      RECT 2446.4800 716.5200 2495.2200 717.6000 ;
      RECT 1007.4200 716.5200 2444.2800 717.6000 ;
      RECT 965.0200 716.5200 1005.2200 717.6000 ;
      RECT 157.4200 716.5200 962.8200 717.6000 ;
      RECT 5.3000 716.5200 155.2200 717.6000 ;
      RECT 0.0000 716.5200 1.7000 717.6000 ;
      RECT 0.0000 716.2500 3370.4200 716.5200 ;
      RECT 1.1000 715.3500 3370.4200 716.2500 ;
      RECT 0.0000 714.8800 3370.4200 715.3500 ;
      RECT 3364.7200 713.8000 3370.4200 714.8800 ;
      RECT 3307.6200 713.8000 3361.1200 714.8800 ;
      RECT 2494.8200 713.8000 3305.4200 714.8800 ;
      RECT 2449.0800 713.8000 2492.6200 714.8800 ;
      RECT 1004.8200 713.8000 2446.8800 714.8800 ;
      RECT 967.6200 713.8000 1002.6200 714.8800 ;
      RECT 154.8200 713.8000 965.4200 714.8800 ;
      RECT 9.3000 713.8000 152.6200 714.8800 ;
      RECT 0.0000 713.8000 5.7000 714.8800 ;
      RECT 0.0000 712.1600 3370.4200 713.8000 ;
      RECT 3368.7200 711.0800 3370.4200 712.1600 ;
      RECT 3305.0200 711.0800 3365.1200 712.1600 ;
      RECT 2497.4200 711.0800 3302.8200 712.1600 ;
      RECT 2446.4800 711.0800 2495.2200 712.1600 ;
      RECT 1007.4200 711.0800 2444.2800 712.1600 ;
      RECT 965.0200 711.0800 1005.2200 712.1600 ;
      RECT 157.4200 711.0800 962.8200 712.1600 ;
      RECT 5.3000 711.0800 155.2200 712.1600 ;
      RECT 0.0000 711.0800 1.7000 712.1600 ;
      RECT 0.0000 709.4400 3370.4200 711.0800 ;
      RECT 3364.7200 708.3600 3370.4200 709.4400 ;
      RECT 3307.6200 708.3600 3361.1200 709.4400 ;
      RECT 2494.8200 708.3600 3305.4200 709.4400 ;
      RECT 2449.0800 708.3600 2492.6200 709.4400 ;
      RECT 1004.8200 708.3600 2446.8800 709.4400 ;
      RECT 967.6200 708.3600 1002.6200 709.4400 ;
      RECT 154.8200 708.3600 965.4200 709.4400 ;
      RECT 9.3000 708.3600 152.6200 709.4400 ;
      RECT 0.0000 708.3600 5.7000 709.4400 ;
      RECT 0.0000 706.7200 3370.4200 708.3600 ;
      RECT 3368.7200 705.6400 3370.4200 706.7200 ;
      RECT 3305.0200 705.6400 3365.1200 706.7200 ;
      RECT 2497.4200 705.6400 3302.8200 706.7200 ;
      RECT 2446.4800 705.6400 2495.2200 706.7200 ;
      RECT 1007.4200 705.6400 2444.2800 706.7200 ;
      RECT 965.0200 705.6400 1005.2200 706.7200 ;
      RECT 157.4200 705.6400 962.8200 706.7200 ;
      RECT 5.3000 705.6400 155.2200 706.7200 ;
      RECT 0.0000 705.6400 1.7000 706.7200 ;
      RECT 0.0000 705.2700 3370.4200 705.6400 ;
      RECT 1.1000 704.3700 3370.4200 705.2700 ;
      RECT 0.0000 704.0000 3370.4200 704.3700 ;
      RECT 3364.7200 702.9200 3370.4200 704.0000 ;
      RECT 3307.6200 702.9200 3361.1200 704.0000 ;
      RECT 2494.8200 702.9200 3305.4200 704.0000 ;
      RECT 2449.0800 702.9200 2492.6200 704.0000 ;
      RECT 1004.8200 702.9200 2446.8800 704.0000 ;
      RECT 967.6200 702.9200 1002.6200 704.0000 ;
      RECT 154.8200 702.9200 965.4200 704.0000 ;
      RECT 9.3000 702.9200 152.6200 704.0000 ;
      RECT 0.0000 702.9200 5.7000 704.0000 ;
      RECT 0.0000 701.2800 3370.4200 702.9200 ;
      RECT 3368.7200 700.2000 3370.4200 701.2800 ;
      RECT 3305.0200 700.2000 3365.1200 701.2800 ;
      RECT 2497.4200 700.2000 3302.8200 701.2800 ;
      RECT 2446.4800 700.2000 2495.2200 701.2800 ;
      RECT 1007.4200 700.2000 2444.2800 701.2800 ;
      RECT 965.0200 700.2000 1005.2200 701.2800 ;
      RECT 157.4200 700.2000 962.8200 701.2800 ;
      RECT 5.3000 700.2000 155.2200 701.2800 ;
      RECT 0.0000 700.2000 1.7000 701.2800 ;
      RECT 0.0000 698.5600 3370.4200 700.2000 ;
      RECT 3364.7200 697.4800 3370.4200 698.5600 ;
      RECT 3307.6200 697.4800 3361.1200 698.5600 ;
      RECT 2494.8200 697.4800 3305.4200 698.5600 ;
      RECT 2449.0800 697.4800 2492.6200 698.5600 ;
      RECT 1004.8200 697.4800 2446.8800 698.5600 ;
      RECT 967.6200 697.4800 1002.6200 698.5600 ;
      RECT 154.8200 697.4800 965.4200 698.5600 ;
      RECT 9.3000 697.4800 152.6200 698.5600 ;
      RECT 0.0000 697.4800 5.7000 698.5600 ;
      RECT 0.0000 695.8400 3370.4200 697.4800 ;
      RECT 3368.7200 694.7600 3370.4200 695.8400 ;
      RECT 3305.0200 694.7600 3365.1200 695.8400 ;
      RECT 2497.4200 694.7600 3302.8200 695.8400 ;
      RECT 2446.4800 694.7600 2495.2200 695.8400 ;
      RECT 1007.4200 694.7600 2444.2800 695.8400 ;
      RECT 965.0200 694.7600 1005.2200 695.8400 ;
      RECT 157.4200 694.7600 962.8200 695.8400 ;
      RECT 5.3000 694.7600 155.2200 695.8400 ;
      RECT 0.0000 694.7600 1.7000 695.8400 ;
      RECT 0.0000 694.2900 3370.4200 694.7600 ;
      RECT 1.1000 693.3900 3370.4200 694.2900 ;
      RECT 0.0000 693.1200 3370.4200 693.3900 ;
      RECT 3364.7200 692.0400 3370.4200 693.1200 ;
      RECT 3307.6200 692.0400 3361.1200 693.1200 ;
      RECT 2494.8200 692.0400 3305.4200 693.1200 ;
      RECT 2449.0800 692.0400 2492.6200 693.1200 ;
      RECT 1004.8200 692.0400 2446.8800 693.1200 ;
      RECT 967.6200 692.0400 1002.6200 693.1200 ;
      RECT 154.8200 692.0400 965.4200 693.1200 ;
      RECT 9.3000 692.0400 152.6200 693.1200 ;
      RECT 0.0000 692.0400 5.7000 693.1200 ;
      RECT 0.0000 690.4000 3370.4200 692.0400 ;
      RECT 3368.7200 689.3200 3370.4200 690.4000 ;
      RECT 3305.0200 689.3200 3365.1200 690.4000 ;
      RECT 2497.4200 689.3200 3302.8200 690.4000 ;
      RECT 2446.4800 689.3200 2495.2200 690.4000 ;
      RECT 1007.4200 689.3200 2444.2800 690.4000 ;
      RECT 965.0200 689.3200 1005.2200 690.4000 ;
      RECT 157.4200 689.3200 962.8200 690.4000 ;
      RECT 5.3000 689.3200 155.2200 690.4000 ;
      RECT 0.0000 689.3200 1.7000 690.4000 ;
      RECT 0.0000 687.6800 3370.4200 689.3200 ;
      RECT 3364.7200 686.6000 3370.4200 687.6800 ;
      RECT 3307.6200 686.6000 3361.1200 687.6800 ;
      RECT 2494.8200 686.6000 3305.4200 687.6800 ;
      RECT 2449.0800 686.6000 2492.6200 687.6800 ;
      RECT 1004.8200 686.6000 2446.8800 687.6800 ;
      RECT 967.6200 686.6000 1002.6200 687.6800 ;
      RECT 154.8200 686.6000 965.4200 687.6800 ;
      RECT 9.3000 686.6000 152.6200 687.6800 ;
      RECT 0.0000 686.6000 5.7000 687.6800 ;
      RECT 0.0000 684.9600 3370.4200 686.6000 ;
      RECT 3368.7200 683.8800 3370.4200 684.9600 ;
      RECT 3305.0200 683.8800 3365.1200 684.9600 ;
      RECT 2497.4200 683.8800 3302.8200 684.9600 ;
      RECT 2446.4800 683.8800 2495.2200 684.9600 ;
      RECT 1007.4200 683.8800 2444.2800 684.9600 ;
      RECT 965.0200 683.8800 1005.2200 684.9600 ;
      RECT 157.4200 683.8800 962.8200 684.9600 ;
      RECT 5.3000 683.8800 155.2200 684.9600 ;
      RECT 0.0000 683.8800 1.7000 684.9600 ;
      RECT 0.0000 683.3100 3370.4200 683.8800 ;
      RECT 1.1000 682.4100 3370.4200 683.3100 ;
      RECT 0.0000 682.2400 3370.4200 682.4100 ;
      RECT 3364.7200 681.1600 3370.4200 682.2400 ;
      RECT 3307.6200 681.1600 3361.1200 682.2400 ;
      RECT 2494.8200 681.1600 3305.4200 682.2400 ;
      RECT 2449.0800 681.1600 2492.6200 682.2400 ;
      RECT 1004.8200 681.1600 2446.8800 682.2400 ;
      RECT 967.6200 681.1600 1002.6200 682.2400 ;
      RECT 154.8200 681.1600 965.4200 682.2400 ;
      RECT 9.3000 681.1600 152.6200 682.2400 ;
      RECT 0.0000 681.1600 5.7000 682.2400 ;
      RECT 0.0000 679.5200 3370.4200 681.1600 ;
      RECT 3368.7200 678.4400 3370.4200 679.5200 ;
      RECT 3305.0200 678.4400 3365.1200 679.5200 ;
      RECT 2497.4200 678.4400 3302.8200 679.5200 ;
      RECT 2446.4800 678.4400 2495.2200 679.5200 ;
      RECT 1007.4200 678.4400 2444.2800 679.5200 ;
      RECT 965.0200 678.4400 1005.2200 679.5200 ;
      RECT 157.4200 678.4400 962.8200 679.5200 ;
      RECT 5.3000 678.4400 155.2200 679.5200 ;
      RECT 0.0000 678.4400 1.7000 679.5200 ;
      RECT 0.0000 676.8000 3370.4200 678.4400 ;
      RECT 3364.7200 675.7200 3370.4200 676.8000 ;
      RECT 3307.6200 675.7200 3361.1200 676.8000 ;
      RECT 2494.8200 675.7200 3305.4200 676.8000 ;
      RECT 2449.0800 675.7200 2492.6200 676.8000 ;
      RECT 1004.8200 675.7200 2446.8800 676.8000 ;
      RECT 967.6200 675.7200 1002.6200 676.8000 ;
      RECT 154.8200 675.7200 965.4200 676.8000 ;
      RECT 9.3000 675.7200 152.6200 676.8000 ;
      RECT 0.0000 675.7200 5.7000 676.8000 ;
      RECT 0.0000 674.0800 3370.4200 675.7200 ;
      RECT 3368.7200 673.0000 3370.4200 674.0800 ;
      RECT 3305.0200 673.0000 3365.1200 674.0800 ;
      RECT 2497.4200 673.0000 3302.8200 674.0800 ;
      RECT 2446.4800 673.0000 2495.2200 674.0800 ;
      RECT 1007.4200 673.0000 2444.2800 674.0800 ;
      RECT 965.0200 673.0000 1005.2200 674.0800 ;
      RECT 157.4200 673.0000 962.8200 674.0800 ;
      RECT 5.3000 673.0000 155.2200 674.0800 ;
      RECT 0.0000 673.0000 1.7000 674.0800 ;
      RECT 0.0000 672.9400 3370.4200 673.0000 ;
      RECT 1.1000 672.0400 3370.4200 672.9400 ;
      RECT 0.0000 671.3600 3370.4200 672.0400 ;
      RECT 3364.7200 670.2800 3370.4200 671.3600 ;
      RECT 3307.6200 670.2800 3361.1200 671.3600 ;
      RECT 2494.8200 670.2800 3305.4200 671.3600 ;
      RECT 2449.0800 670.2800 2492.6200 671.3600 ;
      RECT 1004.8200 670.2800 2446.8800 671.3600 ;
      RECT 967.6200 670.2800 1002.6200 671.3600 ;
      RECT 154.8200 670.2800 965.4200 671.3600 ;
      RECT 9.3000 670.2800 152.6200 671.3600 ;
      RECT 0.0000 670.2800 5.7000 671.3600 ;
      RECT 0.0000 668.6400 3370.4200 670.2800 ;
      RECT 3368.7200 667.5600 3370.4200 668.6400 ;
      RECT 3305.0200 667.5600 3365.1200 668.6400 ;
      RECT 2497.4200 667.5600 3302.8200 668.6400 ;
      RECT 2446.4800 667.5600 2495.2200 668.6400 ;
      RECT 1007.4200 667.5600 2444.2800 668.6400 ;
      RECT 965.0200 667.5600 1005.2200 668.6400 ;
      RECT 157.4200 667.5600 962.8200 668.6400 ;
      RECT 5.3000 667.5600 155.2200 668.6400 ;
      RECT 0.0000 667.5600 1.7000 668.6400 ;
      RECT 0.0000 665.9200 3370.4200 667.5600 ;
      RECT 3364.7200 664.8400 3370.4200 665.9200 ;
      RECT 3307.6200 664.8400 3361.1200 665.9200 ;
      RECT 2494.8200 664.8400 3305.4200 665.9200 ;
      RECT 2449.0800 664.8400 2492.6200 665.9200 ;
      RECT 1004.8200 664.8400 2446.8800 665.9200 ;
      RECT 967.6200 664.8400 1002.6200 665.9200 ;
      RECT 154.8200 664.8400 965.4200 665.9200 ;
      RECT 9.3000 664.8400 152.6200 665.9200 ;
      RECT 0.0000 664.8400 5.7000 665.9200 ;
      RECT 0.0000 663.2000 3370.4200 664.8400 ;
      RECT 3368.7200 662.1200 3370.4200 663.2000 ;
      RECT 3305.0200 662.1200 3365.1200 663.2000 ;
      RECT 2497.4200 662.1200 3302.8200 663.2000 ;
      RECT 2446.4800 662.1200 2495.2200 663.2000 ;
      RECT 1007.4200 662.1200 2444.2800 663.2000 ;
      RECT 965.0200 662.1200 1005.2200 663.2000 ;
      RECT 157.4200 662.1200 962.8200 663.2000 ;
      RECT 5.3000 662.1200 155.2200 663.2000 ;
      RECT 0.0000 662.1200 1.7000 663.2000 ;
      RECT 0.0000 661.9600 3370.4200 662.1200 ;
      RECT 1.1000 661.0600 3370.4200 661.9600 ;
      RECT 0.0000 660.4800 3370.4200 661.0600 ;
      RECT 3364.7200 659.4000 3370.4200 660.4800 ;
      RECT 3307.6200 659.4000 3361.1200 660.4800 ;
      RECT 2494.8200 659.4000 3305.4200 660.4800 ;
      RECT 2449.0800 659.4000 2492.6200 660.4800 ;
      RECT 1004.8200 659.4000 2446.8800 660.4800 ;
      RECT 967.6200 659.4000 1002.6200 660.4800 ;
      RECT 154.8200 659.4000 965.4200 660.4800 ;
      RECT 9.3000 659.4000 152.6200 660.4800 ;
      RECT 0.0000 659.4000 5.7000 660.4800 ;
      RECT 0.0000 657.7600 3370.4200 659.4000 ;
      RECT 3368.7200 656.6800 3370.4200 657.7600 ;
      RECT 3305.0200 656.6800 3365.1200 657.7600 ;
      RECT 2497.4200 656.6800 3302.8200 657.7600 ;
      RECT 2446.4800 656.6800 2495.2200 657.7600 ;
      RECT 1007.4200 656.6800 2444.2800 657.7600 ;
      RECT 965.0200 656.6800 1005.2200 657.7600 ;
      RECT 157.4200 656.6800 962.8200 657.7600 ;
      RECT 5.3000 656.6800 155.2200 657.7600 ;
      RECT 0.0000 656.6800 1.7000 657.7600 ;
      RECT 0.0000 655.0400 3370.4200 656.6800 ;
      RECT 3364.7200 653.9600 3370.4200 655.0400 ;
      RECT 3307.6200 653.9600 3361.1200 655.0400 ;
      RECT 2494.8200 653.9600 3305.4200 655.0400 ;
      RECT 2449.0800 653.9600 2492.6200 655.0400 ;
      RECT 1004.8200 653.9600 2446.8800 655.0400 ;
      RECT 967.6200 653.9600 1002.6200 655.0400 ;
      RECT 154.8200 653.9600 965.4200 655.0400 ;
      RECT 9.3000 653.9600 152.6200 655.0400 ;
      RECT 0.0000 653.9600 5.7000 655.0400 ;
      RECT 0.0000 653.1400 3370.4200 653.9600 ;
      RECT 1077.7200 652.8800 3370.4200 653.1400 ;
      RECT 2436.3200 652.3200 3370.4200 652.8800 ;
      RECT 0.0000 652.3200 1015.2800 653.1400 ;
      RECT 1077.7200 652.0600 1295.6000 652.8800 ;
      RECT 1017.4800 652.0600 1075.5200 653.1400 ;
      RECT 1007.4200 652.0600 1015.2800 652.3200 ;
      RECT 2436.3200 651.8000 2444.2800 652.3200 ;
      RECT 2178.6800 651.8000 2434.1200 652.8800 ;
      RECT 1958.4600 651.8000 2176.4800 652.8800 ;
      RECT 1738.2400 651.8000 1956.2600 652.8800 ;
      RECT 1518.0200 651.8000 1736.0400 652.8800 ;
      RECT 1297.8000 651.8000 1515.8200 652.8800 ;
      RECT 1007.4200 651.8000 1295.6000 652.0600 ;
      RECT 3368.7200 651.2400 3370.4200 652.3200 ;
      RECT 3305.0200 651.2400 3365.1200 652.3200 ;
      RECT 2497.4200 651.2400 3302.8200 652.3200 ;
      RECT 2446.4800 651.2400 2495.2200 652.3200 ;
      RECT 1007.4200 651.2400 2444.2800 651.8000 ;
      RECT 965.0200 651.2400 1005.2200 652.3200 ;
      RECT 157.4200 651.2400 962.8200 652.3200 ;
      RECT 5.3000 651.2400 155.2200 652.3200 ;
      RECT 0.0000 651.2400 1.7000 652.3200 ;
      RECT 0.0000 650.9800 3370.4200 651.2400 ;
      RECT 1.1000 650.0800 3370.4200 650.9800 ;
      RECT 0.0000 650.0700 3370.4200 650.0800 ;
      RECT 0.0000 649.9700 1062.9600 650.0700 ;
      RECT 1285.3800 649.8100 3370.4200 650.0700 ;
      RECT 2446.4800 649.6000 3370.4200 649.8100 ;
      RECT 0.0000 649.6000 1005.2200 649.9700 ;
      RECT 3364.7200 648.5200 3370.4200 649.6000 ;
      RECT 3307.6200 648.5200 3361.1200 649.6000 ;
      RECT 2494.8200 648.5200 3305.4200 649.6000 ;
      RECT 2449.0800 648.5200 2492.6200 649.6000 ;
      RECT 2446.4800 648.5200 2446.8800 649.6000 ;
      RECT 1004.8200 648.5200 1005.2200 649.6000 ;
      RECT 967.6200 648.5200 1002.6200 649.6000 ;
      RECT 154.8200 648.5200 965.4200 649.6000 ;
      RECT 9.3000 648.5200 152.6200 649.6000 ;
      RECT 0.0000 648.5200 5.7000 649.6000 ;
      RECT 1071.3600 647.8700 1279.3800 650.0700 ;
      RECT 1065.1600 647.7700 1283.0400 647.8700 ;
      RECT 1011.2200 647.7700 1059.1600 649.9700 ;
      RECT 0.0000 647.7700 1005.2200 648.5200 ;
      RECT 2392.5400 647.6100 2440.4800 649.8100 ;
      RECT 2172.3200 647.6100 2380.3400 649.8100 ;
      RECT 1952.1000 647.6100 2160.1200 649.8100 ;
      RECT 1731.8800 647.6100 1939.9000 649.8100 ;
      RECT 1511.6600 647.6100 1719.6800 649.8100 ;
      RECT 1291.4400 647.6100 1499.4600 649.8100 ;
      RECT 0.0000 647.6100 1283.0400 647.7700 ;
      RECT 0.0000 647.5700 2444.2800 647.6100 ;
      RECT 1067.7600 647.4700 2444.2800 647.5700 ;
      RECT 2446.4800 647.3300 3370.4200 648.5200 ;
      RECT 1287.9800 647.3300 2444.2800 647.4700 ;
      RECT 1287.9800 647.2100 3370.4200 647.3300 ;
      RECT 2449.0800 646.8800 3370.4200 647.2100 ;
      RECT 0.0000 646.8800 1002.6200 647.5700 ;
      RECT 3368.7200 645.8000 3370.4200 646.8800 ;
      RECT 3305.0200 645.8000 3365.1200 646.8800 ;
      RECT 2497.4200 645.8000 3302.8200 646.8800 ;
      RECT 2449.0800 645.8000 2495.2200 646.8800 ;
      RECT 965.0200 645.8000 1002.6200 646.8800 ;
      RECT 157.4200 645.8000 962.8200 646.8800 ;
      RECT 5.3000 645.8000 155.2200 646.8800 ;
      RECT 0.0000 645.8000 1.7000 646.8800 ;
      RECT 1011.2200 645.3700 1059.1600 647.5700 ;
      RECT 0.0000 645.3700 1002.6200 645.8000 ;
      RECT 1071.3600 645.2700 1279.3800 647.4700 ;
      RECT 1007.4200 645.2700 1065.5600 645.3700 ;
      RECT 2449.0800 645.0100 3370.4200 645.8000 ;
      RECT 2392.5400 645.0100 2440.4800 647.2100 ;
      RECT 2172.3200 645.0100 2380.3400 647.2100 ;
      RECT 1952.1000 645.0100 2166.5200 647.2100 ;
      RECT 1731.8800 645.0100 1939.9000 647.2100 ;
      RECT 1511.6600 645.0100 1719.6800 647.2100 ;
      RECT 1291.4400 645.0100 1499.4600 647.2100 ;
      RECT 1007.4200 645.0100 1285.6400 645.2700 ;
      RECT 1007.4200 644.5000 3370.4200 645.0100 ;
      RECT 0.0000 644.5000 1005.2200 645.3700 ;
      RECT 0.0000 644.1600 3370.4200 644.5000 ;
      RECT 3364.7200 643.0800 3370.4200 644.1600 ;
      RECT 3307.6200 643.0800 3361.1200 644.1600 ;
      RECT 2494.8200 643.0800 3305.4200 644.1600 ;
      RECT 2449.0800 643.0800 2492.6200 644.1600 ;
      RECT 1004.8200 643.0800 2446.8800 644.1600 ;
      RECT 967.6200 643.0800 1002.6200 644.1600 ;
      RECT 154.8200 643.0800 965.4200 644.1600 ;
      RECT 9.3000 643.0800 152.6200 644.1600 ;
      RECT 0.0000 643.0800 5.7000 644.1600 ;
      RECT 0.0000 641.4400 3370.4200 643.0800 ;
      RECT 3368.7200 640.3600 3370.4200 641.4400 ;
      RECT 3305.0200 640.3600 3365.1200 641.4400 ;
      RECT 2497.4200 640.3600 3302.8200 641.4400 ;
      RECT 2446.4800 640.3600 2495.2200 641.4400 ;
      RECT 1007.4200 640.3600 2444.2800 641.4400 ;
      RECT 965.0200 640.3600 1005.2200 641.4400 ;
      RECT 157.4200 640.3600 962.8200 641.4400 ;
      RECT 5.3000 640.3600 155.2200 641.4400 ;
      RECT 0.0000 640.3600 1.7000 641.4400 ;
      RECT 0.0000 640.0400 3370.4200 640.3600 ;
      RECT 0.0000 640.0000 1.7000 640.0400 ;
      RECT 1285.3800 639.7800 3370.4200 640.0400 ;
      RECT 1.1000 639.1000 1.7000 640.0000 ;
      RECT 2446.4800 638.7200 3370.4200 639.7800 ;
      RECT 0.0000 637.8400 1.7000 639.1000 ;
      RECT 3364.7200 637.6400 3370.4200 638.7200 ;
      RECT 3307.6200 637.6400 3361.1200 638.7200 ;
      RECT 2494.8200 637.6400 3305.4200 638.7200 ;
      RECT 2449.0800 637.6400 2492.6200 638.7200 ;
      RECT 2446.4800 637.6400 2446.8800 638.7200 ;
      RECT 2446.4800 637.5800 3370.4200 637.6400 ;
      RECT 1004.8200 637.5800 1283.0400 637.8400 ;
      RECT 1004.8200 637.5400 3370.4200 637.5800 ;
      RECT 1065.0600 637.4400 3370.4200 637.5400 ;
      RECT 1004.8200 637.4400 1062.6600 637.5400 ;
      RECT 9.3000 637.4400 1002.6200 637.8400 ;
      RECT 1287.9800 637.2800 3370.4200 637.4400 ;
      RECT 1945.8000 637.1800 3370.4200 637.2800 ;
      RECT 1287.9800 637.1800 1943.4000 637.2800 ;
      RECT 2449.0800 636.0000 3370.4200 637.1800 ;
      RECT 0.0000 636.0000 5.7000 637.8400 ;
      RECT 5.3000 635.2400 5.7000 636.0000 ;
      RECT 2449.0800 634.9800 2495.2200 636.0000 ;
      RECT 1065.0600 634.9800 1285.6400 635.2400 ;
      RECT 3368.7200 634.9200 3370.4200 636.0000 ;
      RECT 3305.0200 634.9200 3365.1200 636.0000 ;
      RECT 2497.4200 634.9200 3302.8200 636.0000 ;
      RECT 2446.4800 634.9200 2495.2200 634.9800 ;
      RECT 5.3000 634.9200 1005.2200 635.2400 ;
      RECT 0.0000 634.9200 1.7000 636.0000 ;
      RECT 1007.4200 634.4100 1062.6600 635.2400 ;
      RECT 0.0000 634.4100 1005.2200 634.9200 ;
      RECT 2446.4800 634.1300 3370.4200 634.9200 ;
      RECT 1945.8000 634.1300 2444.2800 634.9800 ;
      RECT 1065.0600 633.5400 1943.4000 634.9800 ;
      RECT 0.0000 633.5400 1062.6600 634.4100 ;
      RECT 1945.8000 633.2800 3370.4200 634.1300 ;
      RECT 0.0000 633.2800 1943.4000 633.5400 ;
      RECT 3364.7200 632.2000 3370.4200 633.2800 ;
      RECT 3307.6200 632.2000 3361.1200 633.2800 ;
      RECT 2494.8200 632.2000 3305.4200 633.2800 ;
      RECT 2449.0800 632.2000 2492.6200 633.2800 ;
      RECT 1004.8200 632.2000 2446.8800 633.2800 ;
      RECT 667.6200 632.2000 1002.6200 633.2800 ;
      RECT 504.8200 632.2000 665.4200 633.2800 ;
      RECT 9.3000 632.2000 502.6200 633.2800 ;
      RECT 0.0000 632.2000 5.7000 633.2800 ;
      RECT 0.0000 630.5800 3370.4200 632.2000 ;
      RECT 1287.9800 630.5600 3370.4200 630.5800 ;
      RECT 0.0000 630.5600 1065.5600 630.5800 ;
      RECT 1287.9800 630.3200 2444.2800 630.5600 ;
      RECT 3368.7200 629.4800 3370.4200 630.5600 ;
      RECT 3305.0200 629.4800 3365.1200 630.5600 ;
      RECT 2497.4200 629.4800 3302.8200 630.5600 ;
      RECT 2446.4800 629.4800 2495.2200 630.5600 ;
      RECT 2168.7200 629.4800 2444.2800 630.3200 ;
      RECT 1007.4200 629.4800 1065.5600 630.5600 ;
      RECT 665.0200 629.4800 1005.2200 630.5600 ;
      RECT 507.4200 629.4800 662.8200 630.5600 ;
      RECT 5.3000 629.4800 505.2200 630.5600 ;
      RECT 0.0000 629.4800 1.7000 630.5600 ;
      RECT 0.0000 629.4300 1065.5600 629.4800 ;
      RECT 2168.7200 629.2700 3370.4200 629.4800 ;
      RECT 1287.9800 629.2700 1946.3000 630.3200 ;
      RECT 0.0000 629.0200 1002.6200 629.4300 ;
      RECT 1071.3600 628.3800 1279.3800 630.5800 ;
      RECT 1062.4600 628.3800 1065.5600 629.4300 ;
      RECT 1952.1000 628.1200 2160.1200 630.3200 ;
      RECT 1943.2000 628.1200 1946.3000 629.2700 ;
      RECT 1.1000 628.1200 1002.6200 629.0200 ;
      RECT 1062.4600 627.9800 1285.6400 628.3800 ;
      RECT 2449.0800 627.8400 3370.4200 629.2700 ;
      RECT 0.0000 627.8400 1002.6200 628.1200 ;
      RECT 1943.2000 627.7200 2166.5200 628.1200 ;
      RECT 1062.4600 627.2300 1062.9600 627.9800 ;
      RECT 1011.2200 627.2300 1059.1600 629.4300 ;
      RECT 2392.5400 627.0700 2440.4800 629.2700 ;
      RECT 2172.3200 627.0700 2380.3400 629.2700 ;
      RECT 2166.1200 627.0700 2166.5200 627.7200 ;
      RECT 1943.2000 627.0700 1943.7000 627.7200 ;
      RECT 1731.8800 627.0700 1939.9000 629.2700 ;
      RECT 1511.6600 627.0700 1719.6800 629.2700 ;
      RECT 1291.4400 627.0700 1499.4600 629.2700 ;
      RECT 1285.3800 627.0700 1285.6400 627.9800 ;
      RECT 1004.8200 627.0300 1062.9600 627.2300 ;
      RECT 3364.7200 626.7600 3370.4200 627.8400 ;
      RECT 3307.6200 626.7600 3361.1200 627.8400 ;
      RECT 2494.8200 626.7600 3305.4200 627.8400 ;
      RECT 2449.0800 626.7600 2492.6200 627.8400 ;
      RECT 2166.1200 626.7600 2446.8800 627.0700 ;
      RECT 1004.8200 626.7600 1005.2200 627.0300 ;
      RECT 667.6200 626.7600 1002.6200 627.8400 ;
      RECT 504.8200 626.7600 665.4200 627.8400 ;
      RECT 9.3000 626.7600 502.6200 627.8400 ;
      RECT 0.0000 626.7600 5.7000 627.8400 ;
      RECT 2166.1200 626.6700 3370.4200 626.7600 ;
      RECT 1285.3800 626.6700 1943.7000 627.0700 ;
      RECT 1071.3600 625.7800 1279.3800 627.9800 ;
      RECT 1952.1000 625.5200 2160.1200 627.7200 ;
      RECT 2446.4800 625.1200 3370.4200 626.6700 ;
      RECT 0.0000 625.1200 1005.2200 626.7600 ;
      RECT 1065.1600 624.8300 1283.0400 625.7800 ;
      RECT 1011.2200 624.8300 1059.1600 627.0300 ;
      RECT 2392.5400 624.4700 2440.4800 626.6700 ;
      RECT 2172.3200 624.4700 2380.3400 626.6700 ;
      RECT 1945.9000 624.4700 2163.9200 625.5200 ;
      RECT 1731.8800 624.4700 1939.9000 626.6700 ;
      RECT 1511.6600 624.4700 1719.6800 626.6700 ;
      RECT 1291.4400 624.4700 1499.4600 626.6700 ;
      RECT 1007.4200 624.4700 1283.0400 624.8300 ;
      RECT 3368.7200 624.0400 3370.4200 625.1200 ;
      RECT 3305.0200 624.0400 3365.1200 625.1200 ;
      RECT 2497.4200 624.0400 3302.8200 625.1200 ;
      RECT 2446.4800 624.0400 2495.2200 625.1200 ;
      RECT 1007.4200 624.0400 2444.2800 624.4700 ;
      RECT 665.0200 624.0400 1005.2200 625.1200 ;
      RECT 507.4200 624.0400 662.8200 625.1200 ;
      RECT 5.3000 624.0400 505.2200 625.1200 ;
      RECT 0.0000 624.0400 1.7000 625.1200 ;
      RECT 0.0000 622.4000 3370.4200 624.0400 ;
      RECT 1004.8200 622.0600 2446.8800 622.4000 ;
      RECT 1057.5000 621.8000 2446.8800 622.0600 ;
      RECT 3364.7200 621.3200 3370.4200 622.4000 ;
      RECT 3307.6200 621.3200 3361.1200 622.4000 ;
      RECT 2494.8200 621.3200 3305.4200 622.4000 ;
      RECT 2449.0800 621.3200 2492.6200 622.4000 ;
      RECT 2396.3000 621.3200 2446.8800 621.8000 ;
      RECT 1004.8200 621.3200 1055.3000 622.0600 ;
      RECT 667.6200 621.3200 1002.6200 622.4000 ;
      RECT 504.8200 621.3200 665.4200 622.4000 ;
      RECT 9.3000 621.3200 502.6200 622.4000 ;
      RECT 0.0000 621.3200 5.7000 622.4000 ;
      RECT 1057.5000 620.9800 1293.0000 621.8000 ;
      RECT 0.0000 620.9800 1055.3000 621.3200 ;
      RECT 0.0000 620.9000 1293.0000 620.9800 ;
      RECT 2396.3000 620.7200 3370.4200 621.3200 ;
      RECT 2176.0800 620.7200 2394.1000 621.8000 ;
      RECT 1735.6400 620.7200 2173.8800 621.8000 ;
      RECT 1515.4200 620.7200 1733.4400 621.8000 ;
      RECT 1295.2000 620.7200 1513.2200 621.8000 ;
      RECT 1075.1200 620.7200 1293.0000 620.9000 ;
      RECT 1075.1200 620.6400 3370.4200 620.7200 ;
      RECT 1075.1200 619.8200 1953.6600 620.6400 ;
      RECT 0.0000 619.8200 1072.9200 620.9000 ;
      RECT 1955.8600 619.6800 3370.4200 620.6400 ;
      RECT 0.0000 619.6800 1953.6600 619.8200 ;
      RECT 1955.8600 619.5600 2444.2800 619.6800 ;
      RECT 1007.4200 619.5600 1953.6600 619.6800 ;
      RECT 0.0000 618.6500 1.7000 619.6800 ;
      RECT 3368.7200 618.6000 3370.4200 619.6800 ;
      RECT 3305.0200 618.6000 3365.1200 619.6800 ;
      RECT 2497.4200 618.6000 3302.8200 619.6800 ;
      RECT 2446.4800 618.6000 2495.2200 619.6800 ;
      RECT 1007.4200 618.6000 2444.2800 619.5600 ;
      RECT 665.0200 618.6000 1005.2200 619.6800 ;
      RECT 507.4200 618.6000 662.8200 619.6800 ;
      RECT 5.3000 618.6000 505.2200 619.6800 ;
      RECT 1.1000 618.6000 1.7000 618.6500 ;
      RECT 1.1000 617.7500 3370.4200 618.6000 ;
      RECT 0.0000 616.9600 3370.4200 617.7500 ;
      RECT 3364.7200 615.8800 3370.4200 616.9600 ;
      RECT 3307.6200 615.8800 3361.1200 616.9600 ;
      RECT 2494.8200 615.8800 3305.4200 616.9600 ;
      RECT 2449.0800 615.8800 2492.6200 616.9600 ;
      RECT 1004.8200 615.8800 2446.8800 616.9600 ;
      RECT 667.6200 615.8800 1002.6200 616.9600 ;
      RECT 504.8200 615.8800 665.4200 616.9600 ;
      RECT 9.3000 615.8800 502.6200 616.9600 ;
      RECT 0.0000 615.8800 5.7000 616.9600 ;
      RECT 0.0000 614.2400 3370.4200 615.8800 ;
      RECT 3368.7200 613.1600 3370.4200 614.2400 ;
      RECT 3305.0200 613.1600 3365.1200 614.2400 ;
      RECT 2497.4200 613.1600 3302.8200 614.2400 ;
      RECT 2446.4800 613.1600 2495.2200 614.2400 ;
      RECT 1007.4200 613.1600 2444.2800 614.2400 ;
      RECT 665.0200 613.1600 1005.2200 614.2400 ;
      RECT 507.4200 613.1600 662.8200 614.2400 ;
      RECT 5.3000 613.1600 505.2200 614.2400 ;
      RECT 0.0000 613.1600 1.7000 614.2400 ;
      RECT 0.0000 611.5200 3370.4200 613.1600 ;
      RECT 3364.7200 610.4400 3370.4200 611.5200 ;
      RECT 3307.6200 610.4400 3361.1200 611.5200 ;
      RECT 2494.8200 610.4400 3305.4200 611.5200 ;
      RECT 2449.0800 610.4400 2492.6200 611.5200 ;
      RECT 1004.8200 610.4400 2446.8800 611.5200 ;
      RECT 667.6200 610.4400 1002.6200 611.5200 ;
      RECT 504.8200 610.4400 665.4200 611.5200 ;
      RECT 9.3000 610.4400 502.6200 611.5200 ;
      RECT 0.0000 610.4400 5.7000 611.5200 ;
      RECT 0.0000 608.8000 3370.4200 610.4400 ;
      RECT 3368.7200 607.7200 3370.4200 608.8000 ;
      RECT 3305.0200 607.7200 3365.1200 608.8000 ;
      RECT 2497.4200 607.7200 3302.8200 608.8000 ;
      RECT 2446.4800 607.7200 2495.2200 608.8000 ;
      RECT 1007.4200 607.7200 2444.2800 608.8000 ;
      RECT 665.0200 607.7200 1005.2200 608.8000 ;
      RECT 507.4200 607.7200 662.8200 608.8000 ;
      RECT 5.3000 607.7200 505.2200 608.8000 ;
      RECT 0.0000 607.7200 1.7000 608.8000 ;
      RECT 0.0000 607.6700 3370.4200 607.7200 ;
      RECT 1.1000 606.7700 3370.4200 607.6700 ;
      RECT 0.0000 606.0800 3370.4200 606.7700 ;
      RECT 3364.7200 605.0000 3370.4200 606.0800 ;
      RECT 3307.6200 605.0000 3361.1200 606.0800 ;
      RECT 2494.8200 605.0000 3305.4200 606.0800 ;
      RECT 2449.0800 605.0000 2492.6200 606.0800 ;
      RECT 1004.8200 605.0000 2446.8800 606.0800 ;
      RECT 667.6200 605.0000 1002.6200 606.0800 ;
      RECT 504.8200 605.0000 665.4200 606.0800 ;
      RECT 9.3000 605.0000 502.6200 606.0800 ;
      RECT 0.0000 605.0000 5.7000 606.0800 ;
      RECT 0.0000 603.3600 3370.4200 605.0000 ;
      RECT 3368.7200 602.2800 3370.4200 603.3600 ;
      RECT 3305.0200 602.2800 3365.1200 603.3600 ;
      RECT 2497.4200 602.2800 3302.8200 603.3600 ;
      RECT 2446.4800 602.2800 2495.2200 603.3600 ;
      RECT 1007.4200 602.2800 2444.2800 603.3600 ;
      RECT 665.0200 602.2800 1005.2200 603.3600 ;
      RECT 507.4200 602.2800 662.8200 603.3600 ;
      RECT 5.3000 602.2800 505.2200 603.3600 ;
      RECT 0.0000 602.2800 1.7000 603.3600 ;
      RECT 0.0000 600.6400 3370.4200 602.2800 ;
      RECT 3364.7200 599.5600 3370.4200 600.6400 ;
      RECT 3307.6200 599.5600 3361.1200 600.6400 ;
      RECT 2494.8200 599.5600 3305.4200 600.6400 ;
      RECT 2449.0800 599.5600 2492.6200 600.6400 ;
      RECT 1004.8200 599.5600 2446.8800 600.6400 ;
      RECT 667.6200 599.5600 1002.6200 600.6400 ;
      RECT 504.8200 599.5600 665.4200 600.6400 ;
      RECT 9.3000 599.5600 502.6200 600.6400 ;
      RECT 0.0000 599.5600 5.7000 600.6400 ;
      RECT 0.0000 597.9200 3370.4200 599.5600 ;
      RECT 3368.7200 596.8400 3370.4200 597.9200 ;
      RECT 3305.0200 596.8400 3365.1200 597.9200 ;
      RECT 2497.4200 596.8400 3302.8200 597.9200 ;
      RECT 2446.4800 596.8400 2495.2200 597.9200 ;
      RECT 1007.4200 596.8400 2444.2800 597.9200 ;
      RECT 665.0200 596.8400 1005.2200 597.9200 ;
      RECT 507.4200 596.8400 662.8200 597.9200 ;
      RECT 5.3000 596.8400 505.2200 597.9200 ;
      RECT 0.0000 596.8400 1.7000 597.9200 ;
      RECT 0.0000 596.6900 3370.4200 596.8400 ;
      RECT 1.1000 595.7900 3370.4200 596.6900 ;
      RECT 0.0000 595.2000 3370.4200 595.7900 ;
      RECT 3364.7200 594.1200 3370.4200 595.2000 ;
      RECT 3307.6200 594.1200 3361.1200 595.2000 ;
      RECT 2494.8200 594.1200 3305.4200 595.2000 ;
      RECT 2449.0800 594.1200 2492.6200 595.2000 ;
      RECT 1004.8200 594.1200 2446.8800 595.2000 ;
      RECT 667.6200 594.1200 1002.6200 595.2000 ;
      RECT 504.8200 594.1200 665.4200 595.2000 ;
      RECT 9.3000 594.1200 502.6200 595.2000 ;
      RECT 0.0000 594.1200 5.7000 595.2000 ;
      RECT 0.0000 592.4800 3370.4200 594.1200 ;
      RECT 3368.7200 591.4000 3370.4200 592.4800 ;
      RECT 3305.0200 591.4000 3365.1200 592.4800 ;
      RECT 2497.4200 591.4000 3302.8200 592.4800 ;
      RECT 2446.4800 591.4000 2495.2200 592.4800 ;
      RECT 1007.4200 591.4000 2444.2800 592.4800 ;
      RECT 665.0200 591.4000 1005.2200 592.4800 ;
      RECT 507.4200 591.4000 662.8200 592.4800 ;
      RECT 5.3000 591.4000 505.2200 592.4800 ;
      RECT 0.0000 591.4000 1.7000 592.4800 ;
      RECT 0.0000 589.7600 3370.4200 591.4000 ;
      RECT 3364.7200 588.6800 3370.4200 589.7600 ;
      RECT 3307.6200 588.6800 3361.1200 589.7600 ;
      RECT 2494.8200 588.6800 3305.4200 589.7600 ;
      RECT 2449.0800 588.6800 2492.6200 589.7600 ;
      RECT 1004.8200 588.6800 2446.8800 589.7600 ;
      RECT 667.6200 588.6800 1002.6200 589.7600 ;
      RECT 504.8200 588.6800 665.4200 589.7600 ;
      RECT 9.3000 588.6800 502.6200 589.7600 ;
      RECT 0.0000 588.6800 5.7000 589.7600 ;
      RECT 0.0000 587.0400 3370.4200 588.6800 ;
      RECT 3368.7200 585.9600 3370.4200 587.0400 ;
      RECT 3305.0200 585.9600 3365.1200 587.0400 ;
      RECT 2497.4200 585.9600 3302.8200 587.0400 ;
      RECT 2446.4800 585.9600 2495.2200 587.0400 ;
      RECT 1007.4200 585.9600 2444.2800 587.0400 ;
      RECT 665.0200 585.9600 1005.2200 587.0400 ;
      RECT 507.4200 585.9600 662.8200 587.0400 ;
      RECT 5.3000 585.9600 505.2200 587.0400 ;
      RECT 0.0000 585.9600 1.7000 587.0400 ;
      RECT 0.0000 585.7100 3370.4200 585.9600 ;
      RECT 1.1000 584.8100 3370.4200 585.7100 ;
      RECT 0.0000 584.3200 3370.4200 584.8100 ;
      RECT 3364.7200 583.2400 3370.4200 584.3200 ;
      RECT 3307.6200 583.2400 3361.1200 584.3200 ;
      RECT 2494.8200 583.2400 3305.4200 584.3200 ;
      RECT 2449.0800 583.2400 2492.6200 584.3200 ;
      RECT 1004.8200 583.2400 2446.8800 584.3200 ;
      RECT 667.6200 583.2400 1002.6200 584.3200 ;
      RECT 504.8200 583.2400 665.4200 584.3200 ;
      RECT 9.3000 583.2400 502.6200 584.3200 ;
      RECT 0.0000 583.2400 5.7000 584.3200 ;
      RECT 0.0000 581.6000 3370.4200 583.2400 ;
      RECT 3368.7200 580.5200 3370.4200 581.6000 ;
      RECT 3305.0200 580.5200 3365.1200 581.6000 ;
      RECT 2497.4200 580.5200 3302.8200 581.6000 ;
      RECT 2446.4800 580.5200 2495.2200 581.6000 ;
      RECT 1007.4200 580.5200 2444.2800 581.6000 ;
      RECT 665.0200 580.5200 1005.2200 581.6000 ;
      RECT 507.4200 580.5200 662.8200 581.6000 ;
      RECT 5.3000 580.5200 505.2200 581.6000 ;
      RECT 0.0000 580.5200 1.7000 581.6000 ;
      RECT 0.0000 578.8800 3370.4200 580.5200 ;
      RECT 3364.7200 577.8000 3370.4200 578.8800 ;
      RECT 3307.6200 577.8000 3361.1200 578.8800 ;
      RECT 2494.8200 577.8000 3305.4200 578.8800 ;
      RECT 2449.0800 577.8000 2492.6200 578.8800 ;
      RECT 1004.8200 577.8000 2446.8800 578.8800 ;
      RECT 667.6200 577.8000 1002.6200 578.8800 ;
      RECT 504.8200 577.8000 665.4200 578.8800 ;
      RECT 9.3000 577.8000 502.6200 578.8800 ;
      RECT 0.0000 577.8000 5.7000 578.8800 ;
      RECT 0.0000 576.1600 3370.4200 577.8000 ;
      RECT 3368.7200 575.0800 3370.4200 576.1600 ;
      RECT 3305.0200 575.0800 3365.1200 576.1600 ;
      RECT 2497.4200 575.0800 3302.8200 576.1600 ;
      RECT 2446.4800 575.0800 2495.2200 576.1600 ;
      RECT 1007.4200 575.0800 2444.2800 576.1600 ;
      RECT 665.0200 575.0800 1005.2200 576.1600 ;
      RECT 507.4200 575.0800 662.8200 576.1600 ;
      RECT 5.3000 575.0800 505.2200 576.1600 ;
      RECT 0.0000 575.0800 1.7000 576.1600 ;
      RECT 0.0000 574.7300 3370.4200 575.0800 ;
      RECT 1.1000 573.8300 3370.4200 574.7300 ;
      RECT 0.0000 573.4400 3370.4200 573.8300 ;
      RECT 3364.7200 572.3600 3370.4200 573.4400 ;
      RECT 3307.6200 572.3600 3361.1200 573.4400 ;
      RECT 2494.8200 572.3600 3305.4200 573.4400 ;
      RECT 2449.0800 572.3600 2492.6200 573.4400 ;
      RECT 1004.8200 572.3600 2446.8800 573.4400 ;
      RECT 667.6200 572.3600 1002.6200 573.4400 ;
      RECT 504.8200 572.3600 665.4200 573.4400 ;
      RECT 9.3000 572.3600 502.6200 573.4400 ;
      RECT 0.0000 572.3600 5.7000 573.4400 ;
      RECT 0.0000 570.7200 3370.4200 572.3600 ;
      RECT 3368.7200 569.6400 3370.4200 570.7200 ;
      RECT 3305.0200 569.6400 3365.1200 570.7200 ;
      RECT 2497.4200 569.6400 3302.8200 570.7200 ;
      RECT 2446.4800 569.6400 2495.2200 570.7200 ;
      RECT 1007.4200 569.6400 2444.2800 570.7200 ;
      RECT 665.0200 569.6400 1005.2200 570.7200 ;
      RECT 507.4200 569.6400 662.8200 570.7200 ;
      RECT 5.3000 569.6400 505.2200 570.7200 ;
      RECT 0.0000 569.6400 1.7000 570.7200 ;
      RECT 0.0000 568.0000 3370.4200 569.6400 ;
      RECT 3364.7200 566.9200 3370.4200 568.0000 ;
      RECT 3307.6200 566.9200 3361.1200 568.0000 ;
      RECT 2494.8200 566.9200 3305.4200 568.0000 ;
      RECT 2449.0800 566.9200 2492.6200 568.0000 ;
      RECT 1004.8200 566.9200 2446.8800 568.0000 ;
      RECT 667.6200 566.9200 1002.6200 568.0000 ;
      RECT 504.8200 566.9200 665.4200 568.0000 ;
      RECT 9.3000 566.9200 502.6200 568.0000 ;
      RECT 0.0000 566.9200 5.7000 568.0000 ;
      RECT 0.0000 565.2800 3370.4200 566.9200 ;
      RECT 0.0000 564.3600 1.7000 565.2800 ;
      RECT 3368.7200 564.2000 3370.4200 565.2800 ;
      RECT 3305.0200 564.2000 3365.1200 565.2800 ;
      RECT 2497.4200 564.2000 3302.8200 565.2800 ;
      RECT 2446.4800 564.2000 2495.2200 565.2800 ;
      RECT 1007.4200 564.2000 2444.2800 565.2800 ;
      RECT 665.0200 564.2000 1005.2200 565.2800 ;
      RECT 507.4200 564.2000 662.8200 565.2800 ;
      RECT 5.3000 564.2000 505.2200 565.2800 ;
      RECT 1.1000 564.2000 1.7000 564.3600 ;
      RECT 1.1000 563.4600 3370.4200 564.2000 ;
      RECT 0.0000 562.5600 3370.4200 563.4600 ;
      RECT 3364.7200 561.4800 3370.4200 562.5600 ;
      RECT 3307.6200 561.4800 3361.1200 562.5600 ;
      RECT 2494.8200 561.4800 3305.4200 562.5600 ;
      RECT 2449.0800 561.4800 2492.6200 562.5600 ;
      RECT 1004.8200 561.4800 2446.8800 562.5600 ;
      RECT 667.6200 561.4800 1002.6200 562.5600 ;
      RECT 504.8200 561.4800 665.4200 562.5600 ;
      RECT 9.3000 561.4800 502.6200 562.5600 ;
      RECT 0.0000 561.4800 5.7000 562.5600 ;
      RECT 0.0000 559.8400 3370.4200 561.4800 ;
      RECT 3368.7200 558.7600 3370.4200 559.8400 ;
      RECT 3305.0200 558.7600 3365.1200 559.8400 ;
      RECT 2497.4200 558.7600 3302.8200 559.8400 ;
      RECT 2446.4800 558.7600 2495.2200 559.8400 ;
      RECT 1007.4200 558.7600 2444.2800 559.8400 ;
      RECT 665.0200 558.7600 1005.2200 559.8400 ;
      RECT 507.4200 558.7600 662.8200 559.8400 ;
      RECT 5.3000 558.7600 505.2200 559.8400 ;
      RECT 0.0000 558.7600 1.7000 559.8400 ;
      RECT 0.0000 557.1200 3370.4200 558.7600 ;
      RECT 3364.7200 556.0400 3370.4200 557.1200 ;
      RECT 3307.6200 556.0400 3361.1200 557.1200 ;
      RECT 2494.8200 556.0400 3305.4200 557.1200 ;
      RECT 2449.0800 556.0400 2492.6200 557.1200 ;
      RECT 1004.8200 556.0400 2446.8800 557.1200 ;
      RECT 667.6200 556.0400 1002.6200 557.1200 ;
      RECT 504.8200 556.0400 665.4200 557.1200 ;
      RECT 9.3000 556.0400 502.6200 557.1200 ;
      RECT 0.0000 556.0400 5.7000 557.1200 ;
      RECT 0.0000 554.4000 3370.4200 556.0400 ;
      RECT 0.0000 553.3800 1.7000 554.4000 ;
      RECT 3368.7200 553.3200 3370.4200 554.4000 ;
      RECT 3305.0200 553.3200 3365.1200 554.4000 ;
      RECT 2497.4200 553.3200 3302.8200 554.4000 ;
      RECT 2446.4800 553.3200 2495.2200 554.4000 ;
      RECT 1007.4200 553.3200 2444.2800 554.4000 ;
      RECT 665.0200 553.3200 1005.2200 554.4000 ;
      RECT 507.4200 553.3200 662.8200 554.4000 ;
      RECT 5.3000 553.3200 505.2200 554.4000 ;
      RECT 1.1000 553.3200 1.7000 553.3800 ;
      RECT 1.1000 552.4800 3370.4200 553.3200 ;
      RECT 0.0000 551.6800 3370.4200 552.4800 ;
      RECT 3364.7200 550.6000 3370.4200 551.6800 ;
      RECT 3307.6200 550.6000 3361.1200 551.6800 ;
      RECT 2494.8200 550.6000 3305.4200 551.6800 ;
      RECT 2449.0800 550.6000 2492.6200 551.6800 ;
      RECT 1004.8200 550.6000 2446.8800 551.6800 ;
      RECT 667.6200 550.6000 1002.6200 551.6800 ;
      RECT 504.8200 550.6000 665.4200 551.6800 ;
      RECT 9.3000 550.6000 502.6200 551.6800 ;
      RECT 0.0000 550.6000 5.7000 551.6800 ;
      RECT 0.0000 548.9600 3370.4200 550.6000 ;
      RECT 3368.7200 547.8800 3370.4200 548.9600 ;
      RECT 3305.0200 547.8800 3365.1200 548.9600 ;
      RECT 2497.4200 547.8800 3302.8200 548.9600 ;
      RECT 2446.4800 547.8800 2495.2200 548.9600 ;
      RECT 1007.4200 547.8800 2444.2800 548.9600 ;
      RECT 665.0200 547.8800 1005.2200 548.9600 ;
      RECT 507.4200 547.8800 662.8200 548.9600 ;
      RECT 5.3000 547.8800 505.2200 548.9600 ;
      RECT 0.0000 547.8800 1.7000 548.9600 ;
      RECT 0.0000 546.2400 3370.4200 547.8800 ;
      RECT 3364.7200 545.1600 3370.4200 546.2400 ;
      RECT 3307.6200 545.1600 3361.1200 546.2400 ;
      RECT 2494.8200 545.1600 3305.4200 546.2400 ;
      RECT 2449.0800 545.1600 2492.6200 546.2400 ;
      RECT 1004.8200 545.1600 2446.8800 546.2400 ;
      RECT 667.6200 545.1600 1002.6200 546.2400 ;
      RECT 504.8200 545.1600 665.4200 546.2400 ;
      RECT 9.3000 545.1600 502.6200 546.2400 ;
      RECT 0.0000 545.1600 5.7000 546.2400 ;
      RECT 0.0000 543.5200 3370.4200 545.1600 ;
      RECT 3368.7200 542.4400 3370.4200 543.5200 ;
      RECT 3305.0200 542.4400 3365.1200 543.5200 ;
      RECT 2497.4200 542.4400 3302.8200 543.5200 ;
      RECT 2446.4800 542.4400 2495.2200 543.5200 ;
      RECT 1007.4200 542.4400 2444.2800 543.5200 ;
      RECT 665.0200 542.4400 1005.2200 543.5200 ;
      RECT 507.4200 542.4400 662.8200 543.5200 ;
      RECT 5.3000 542.4400 505.2200 543.5200 ;
      RECT 0.0000 542.4400 1.7000 543.5200 ;
      RECT 0.0000 542.4000 3370.4200 542.4400 ;
      RECT 1.1000 541.5000 3370.4200 542.4000 ;
      RECT 0.0000 540.8000 3370.4200 541.5000 ;
      RECT 3364.7200 539.7200 3370.4200 540.8000 ;
      RECT 3307.6200 539.7200 3361.1200 540.8000 ;
      RECT 2494.8200 539.7200 3305.4200 540.8000 ;
      RECT 2449.0800 539.7200 2492.6200 540.8000 ;
      RECT 1004.8200 539.7200 2446.8800 540.8000 ;
      RECT 667.6200 539.7200 1002.6200 540.8000 ;
      RECT 504.8200 539.7200 665.4200 540.8000 ;
      RECT 9.3000 539.7200 502.6200 540.8000 ;
      RECT 0.0000 539.7200 5.7000 540.8000 ;
      RECT 0.0000 538.0800 3370.4200 539.7200 ;
      RECT 3368.7200 537.0000 3370.4200 538.0800 ;
      RECT 3305.0200 537.0000 3365.1200 538.0800 ;
      RECT 2497.4200 537.0000 3302.8200 538.0800 ;
      RECT 2446.4800 537.0000 2495.2200 538.0800 ;
      RECT 1007.4200 537.0000 2444.2800 538.0800 ;
      RECT 665.0200 537.0000 1005.2200 538.0800 ;
      RECT 507.4200 537.0000 662.8200 538.0800 ;
      RECT 5.3000 537.0000 505.2200 538.0800 ;
      RECT 0.0000 537.0000 1.7000 538.0800 ;
      RECT 0.0000 535.3600 3370.4200 537.0000 ;
      RECT 3364.7200 534.2800 3370.4200 535.3600 ;
      RECT 3307.6200 534.2800 3361.1200 535.3600 ;
      RECT 2494.8200 534.2800 3305.4200 535.3600 ;
      RECT 2449.0800 534.2800 2492.6200 535.3600 ;
      RECT 1004.8200 534.2800 2446.8800 535.3600 ;
      RECT 667.6200 534.2800 1002.6200 535.3600 ;
      RECT 504.8200 534.2800 665.4200 535.3600 ;
      RECT 9.3000 534.2800 502.6200 535.3600 ;
      RECT 0.0000 534.2800 5.7000 535.3600 ;
      RECT 0.0000 532.6400 3370.4200 534.2800 ;
      RECT 3368.7200 531.5600 3370.4200 532.6400 ;
      RECT 3305.0200 531.5600 3365.1200 532.6400 ;
      RECT 2497.4200 531.5600 3302.8200 532.6400 ;
      RECT 2446.4800 531.5600 2495.2200 532.6400 ;
      RECT 1007.4200 531.5600 2444.2800 532.6400 ;
      RECT 665.0200 531.5600 1005.2200 532.6400 ;
      RECT 507.4200 531.5600 662.8200 532.6400 ;
      RECT 5.3000 531.5600 505.2200 532.6400 ;
      RECT 0.0000 531.5600 1.7000 532.6400 ;
      RECT 0.0000 531.4200 3370.4200 531.5600 ;
      RECT 1.1000 530.5200 3370.4200 531.4200 ;
      RECT 0.0000 529.9200 3370.4200 530.5200 ;
      RECT 3364.7200 528.8400 3370.4200 529.9200 ;
      RECT 3307.6200 528.8400 3361.1200 529.9200 ;
      RECT 2494.8200 528.8400 3305.4200 529.9200 ;
      RECT 2449.0800 528.8400 2492.6200 529.9200 ;
      RECT 1004.8200 528.8400 2446.8800 529.9200 ;
      RECT 667.6200 528.8400 1002.6200 529.9200 ;
      RECT 504.8200 528.8400 665.4200 529.9200 ;
      RECT 9.3000 528.8400 502.6200 529.9200 ;
      RECT 0.0000 528.8400 5.7000 529.9200 ;
      RECT 0.0000 527.2000 3370.4200 528.8400 ;
      RECT 3368.7200 526.1200 3370.4200 527.2000 ;
      RECT 3305.0200 526.1200 3365.1200 527.2000 ;
      RECT 2497.4200 526.1200 3302.8200 527.2000 ;
      RECT 2446.4800 526.1200 2495.2200 527.2000 ;
      RECT 1007.4200 526.1200 2444.2800 527.2000 ;
      RECT 665.0200 526.1200 1005.2200 527.2000 ;
      RECT 507.4200 526.1200 662.8200 527.2000 ;
      RECT 5.3000 526.1200 505.2200 527.2000 ;
      RECT 0.0000 526.1200 1.7000 527.2000 ;
      RECT 0.0000 524.4800 3370.4200 526.1200 ;
      RECT 3364.7200 523.4000 3370.4200 524.4800 ;
      RECT 3307.6200 523.4000 3361.1200 524.4800 ;
      RECT 2494.8200 523.4000 3305.4200 524.4800 ;
      RECT 2449.0800 523.4000 2492.6200 524.4800 ;
      RECT 1004.8200 523.4000 2446.8800 524.4800 ;
      RECT 667.6200 523.4000 1002.6200 524.4800 ;
      RECT 504.8200 523.4000 665.4200 524.4800 ;
      RECT 9.3000 523.4000 502.6200 524.4800 ;
      RECT 0.0000 523.4000 5.7000 524.4800 ;
      RECT 0.0000 521.7600 3370.4200 523.4000 ;
      RECT 3368.7200 520.6800 3370.4200 521.7600 ;
      RECT 3305.0200 520.6800 3365.1200 521.7600 ;
      RECT 2497.4200 520.6800 3302.8200 521.7600 ;
      RECT 2446.4800 520.6800 2495.2200 521.7600 ;
      RECT 1007.4200 520.6800 2444.2800 521.7600 ;
      RECT 665.0200 520.6800 1005.2200 521.7600 ;
      RECT 507.4200 520.6800 662.8200 521.7600 ;
      RECT 5.3000 520.6800 505.2200 521.7600 ;
      RECT 0.0000 520.6800 1.7000 521.7600 ;
      RECT 0.0000 520.4400 3370.4200 520.6800 ;
      RECT 1.1000 519.5400 3370.4200 520.4400 ;
      RECT 0.0000 519.0400 3370.4200 519.5400 ;
      RECT 3364.7200 517.9600 3370.4200 519.0400 ;
      RECT 3307.6200 517.9600 3361.1200 519.0400 ;
      RECT 2494.8200 517.9600 3305.4200 519.0400 ;
      RECT 2449.0800 517.9600 2492.6200 519.0400 ;
      RECT 1004.8200 517.9600 2446.8800 519.0400 ;
      RECT 667.6200 517.9600 1002.6200 519.0400 ;
      RECT 504.8200 517.9600 665.4200 519.0400 ;
      RECT 9.3000 517.9600 502.6200 519.0400 ;
      RECT 0.0000 517.9600 5.7000 519.0400 ;
      RECT 0.0000 516.3200 3370.4200 517.9600 ;
      RECT 3368.7200 515.2400 3370.4200 516.3200 ;
      RECT 3305.0200 515.2400 3365.1200 516.3200 ;
      RECT 2497.4200 515.2400 3302.8200 516.3200 ;
      RECT 2446.4800 515.2400 2495.2200 516.3200 ;
      RECT 1007.4200 515.2400 2444.2800 516.3200 ;
      RECT 665.0200 515.2400 1005.2200 516.3200 ;
      RECT 507.4200 515.2400 662.8200 516.3200 ;
      RECT 5.3000 515.2400 505.2200 516.3200 ;
      RECT 0.0000 515.2400 1.7000 516.3200 ;
      RECT 0.0000 513.6000 3370.4200 515.2400 ;
      RECT 3364.7200 512.5200 3370.4200 513.6000 ;
      RECT 3307.6200 512.5200 3361.1200 513.6000 ;
      RECT 2494.8200 512.5200 3305.4200 513.6000 ;
      RECT 2449.0800 512.5200 2492.6200 513.6000 ;
      RECT 1004.8200 512.5200 2446.8800 513.6000 ;
      RECT 667.6200 512.5200 1002.6200 513.6000 ;
      RECT 504.8200 512.5200 665.4200 513.6000 ;
      RECT 9.3000 512.5200 502.6200 513.6000 ;
      RECT 0.0000 512.5200 5.7000 513.6000 ;
      RECT 0.0000 510.8800 3370.4200 512.5200 ;
      RECT 0.0000 510.0700 1.7000 510.8800 ;
      RECT 3368.7200 509.8000 3370.4200 510.8800 ;
      RECT 3305.0200 509.8000 3365.1200 510.8800 ;
      RECT 2497.4200 509.8000 3302.8200 510.8800 ;
      RECT 2446.4800 509.8000 2495.2200 510.8800 ;
      RECT 1007.4200 509.8000 2444.2800 510.8800 ;
      RECT 665.0200 509.8000 1005.2200 510.8800 ;
      RECT 507.4200 509.8000 662.8200 510.8800 ;
      RECT 5.3000 509.8000 505.2200 510.8800 ;
      RECT 1.1000 509.8000 1.7000 510.0700 ;
      RECT 1.1000 509.1700 3370.4200 509.8000 ;
      RECT 0.0000 508.1600 3370.4200 509.1700 ;
      RECT 3364.7200 507.0800 3370.4200 508.1600 ;
      RECT 3307.6200 507.0800 3361.1200 508.1600 ;
      RECT 2494.8200 507.0800 3305.4200 508.1600 ;
      RECT 2449.0800 507.0800 2492.6200 508.1600 ;
      RECT 1004.8200 507.0800 2446.8800 508.1600 ;
      RECT 667.6200 507.0800 1002.6200 508.1600 ;
      RECT 504.8200 507.0800 665.4200 508.1600 ;
      RECT 9.3000 507.0800 502.6200 508.1600 ;
      RECT 0.0000 507.0800 5.7000 508.1600 ;
      RECT 0.0000 505.4400 3370.4200 507.0800 ;
      RECT 3368.7200 504.3600 3370.4200 505.4400 ;
      RECT 3305.0200 504.3600 3365.1200 505.4400 ;
      RECT 2497.4200 504.3600 3302.8200 505.4400 ;
      RECT 2446.4800 504.3600 2495.2200 505.4400 ;
      RECT 1007.4200 504.3600 2444.2800 505.4400 ;
      RECT 665.0200 504.3600 1005.2200 505.4400 ;
      RECT 507.4200 504.3600 662.8200 505.4400 ;
      RECT 5.3000 504.3600 505.2200 505.4400 ;
      RECT 0.0000 504.3600 1.7000 505.4400 ;
      RECT 0.0000 502.7200 3370.4200 504.3600 ;
      RECT 3364.7200 501.6400 3370.4200 502.7200 ;
      RECT 3307.6200 501.6400 3361.1200 502.7200 ;
      RECT 2494.8200 501.6400 3305.4200 502.7200 ;
      RECT 2449.0800 501.6400 2492.6200 502.7200 ;
      RECT 1004.8200 501.6400 2446.8800 502.7200 ;
      RECT 667.6200 501.6400 1002.6200 502.7200 ;
      RECT 504.8200 501.6400 665.4200 502.7200 ;
      RECT 9.3000 501.6400 502.6200 502.7200 ;
      RECT 0.0000 501.6400 5.7000 502.7200 ;
      RECT 0.0000 500.0000 3370.4200 501.6400 ;
      RECT 0.0000 499.0900 1.7000 500.0000 ;
      RECT 3368.7200 498.9200 3370.4200 500.0000 ;
      RECT 3305.0200 498.9200 3365.1200 500.0000 ;
      RECT 2497.4200 498.9200 3302.8200 500.0000 ;
      RECT 2446.4800 498.9200 2495.2200 500.0000 ;
      RECT 1007.4200 498.9200 2444.2800 500.0000 ;
      RECT 665.0200 498.9200 1005.2200 500.0000 ;
      RECT 507.4200 498.9200 662.8200 500.0000 ;
      RECT 5.3000 498.9200 505.2200 500.0000 ;
      RECT 1.1000 498.9200 1.7000 499.0900 ;
      RECT 1.1000 498.1900 3370.4200 498.9200 ;
      RECT 0.0000 497.2800 3370.4200 498.1900 ;
      RECT 3364.7200 496.2000 3370.4200 497.2800 ;
      RECT 3307.6200 496.2000 3361.1200 497.2800 ;
      RECT 2494.8200 496.2000 3305.4200 497.2800 ;
      RECT 2449.0800 496.2000 2492.6200 497.2800 ;
      RECT 1004.8200 496.2000 2446.8800 497.2800 ;
      RECT 667.6200 496.2000 1002.6200 497.2800 ;
      RECT 504.8200 496.2000 665.4200 497.2800 ;
      RECT 9.3000 496.2000 502.6200 497.2800 ;
      RECT 0.0000 496.2000 5.7000 497.2800 ;
      RECT 0.0000 494.5600 3370.4200 496.2000 ;
      RECT 3368.7200 493.4800 3370.4200 494.5600 ;
      RECT 3305.0200 493.4800 3365.1200 494.5600 ;
      RECT 2497.4200 493.4800 3302.8200 494.5600 ;
      RECT 2446.4800 493.4800 2495.2200 494.5600 ;
      RECT 1007.4200 493.4800 2444.2800 494.5600 ;
      RECT 665.0200 493.4800 1005.2200 494.5600 ;
      RECT 507.4200 493.4800 662.8200 494.5600 ;
      RECT 5.3000 493.4800 505.2200 494.5600 ;
      RECT 0.0000 493.4800 1.7000 494.5600 ;
      RECT 0.0000 491.8400 3370.4200 493.4800 ;
      RECT 3364.7200 490.7600 3370.4200 491.8400 ;
      RECT 3307.6200 490.7600 3361.1200 491.8400 ;
      RECT 2494.8200 490.7600 3305.4200 491.8400 ;
      RECT 2449.0800 490.7600 2492.6200 491.8400 ;
      RECT 1004.8200 490.7600 2446.8800 491.8400 ;
      RECT 667.6200 490.7600 1002.6200 491.8400 ;
      RECT 504.8200 490.7600 665.4200 491.8400 ;
      RECT 9.3000 490.7600 502.6200 491.8400 ;
      RECT 0.0000 490.7600 5.7000 491.8400 ;
      RECT 0.0000 489.1200 3370.4200 490.7600 ;
      RECT 0.0000 488.1100 1.7000 489.1200 ;
      RECT 3368.7200 488.0400 3370.4200 489.1200 ;
      RECT 3305.0200 488.0400 3365.1200 489.1200 ;
      RECT 2497.4200 488.0400 3302.8200 489.1200 ;
      RECT 2446.4800 488.0400 2495.2200 489.1200 ;
      RECT 1007.4200 488.0400 2444.2800 489.1200 ;
      RECT 665.0200 488.0400 1005.2200 489.1200 ;
      RECT 507.4200 488.0400 662.8200 489.1200 ;
      RECT 5.3000 488.0400 505.2200 489.1200 ;
      RECT 1.1000 488.0400 1.7000 488.1100 ;
      RECT 1.1000 487.2100 3370.4200 488.0400 ;
      RECT 0.0000 486.4000 3370.4200 487.2100 ;
      RECT 3364.7200 485.3200 3370.4200 486.4000 ;
      RECT 3307.6200 485.3200 3361.1200 486.4000 ;
      RECT 2494.8200 485.3200 3305.4200 486.4000 ;
      RECT 2449.0800 485.3200 2492.6200 486.4000 ;
      RECT 1004.8200 485.3200 2446.8800 486.4000 ;
      RECT 667.6200 485.3200 1002.6200 486.4000 ;
      RECT 504.8200 485.3200 665.4200 486.4000 ;
      RECT 9.3000 485.3200 502.6200 486.4000 ;
      RECT 0.0000 485.3200 5.7000 486.4000 ;
      RECT 0.0000 483.6800 3370.4200 485.3200 ;
      RECT 3368.7200 482.6000 3370.4200 483.6800 ;
      RECT 3305.0200 482.6000 3365.1200 483.6800 ;
      RECT 2497.4200 482.6000 3302.8200 483.6800 ;
      RECT 2446.4800 482.6000 2495.2200 483.6800 ;
      RECT 1007.4200 482.6000 2444.2800 483.6800 ;
      RECT 665.0200 482.6000 1005.2200 483.6800 ;
      RECT 507.4200 482.6000 662.8200 483.6800 ;
      RECT 5.3000 482.6000 505.2200 483.6800 ;
      RECT 0.0000 482.6000 1.7000 483.6800 ;
      RECT 0.0000 480.9600 3370.4200 482.6000 ;
      RECT 3364.7200 479.8800 3370.4200 480.9600 ;
      RECT 3307.6200 479.8800 3361.1200 480.9600 ;
      RECT 2494.8200 479.8800 3305.4200 480.9600 ;
      RECT 2449.0800 479.8800 2492.6200 480.9600 ;
      RECT 1004.8200 479.8800 2446.8800 480.9600 ;
      RECT 667.6200 479.8800 1002.6200 480.9600 ;
      RECT 504.8200 479.8800 665.4200 480.9600 ;
      RECT 9.3000 479.8800 502.6200 480.9600 ;
      RECT 0.0000 479.8800 5.7000 480.9600 ;
      RECT 0.0000 478.2400 3370.4200 479.8800 ;
      RECT 3368.7200 477.1600 3370.4200 478.2400 ;
      RECT 3305.0200 477.1600 3365.1200 478.2400 ;
      RECT 2497.4200 477.1600 3302.8200 478.2400 ;
      RECT 2446.4800 477.1600 2495.2200 478.2400 ;
      RECT 1007.4200 477.1600 2444.2800 478.2400 ;
      RECT 665.0200 477.1600 1005.2200 478.2400 ;
      RECT 507.4200 477.1600 662.8200 478.2400 ;
      RECT 5.3000 477.1600 505.2200 478.2400 ;
      RECT 0.0000 477.1600 1.7000 478.2400 ;
      RECT 0.0000 477.1300 3370.4200 477.1600 ;
      RECT 1.1000 476.2300 3370.4200 477.1300 ;
      RECT 0.0000 475.5200 3370.4200 476.2300 ;
      RECT 3364.7200 474.4400 3370.4200 475.5200 ;
      RECT 3307.6200 474.4400 3361.1200 475.5200 ;
      RECT 2494.8200 474.4400 3305.4200 475.5200 ;
      RECT 2449.0800 474.4400 2492.6200 475.5200 ;
      RECT 1004.8200 474.4400 2446.8800 475.5200 ;
      RECT 667.6200 474.4400 1002.6200 475.5200 ;
      RECT 504.8200 474.4400 665.4200 475.5200 ;
      RECT 9.3000 474.4400 502.6200 475.5200 ;
      RECT 0.0000 474.4400 5.7000 475.5200 ;
      RECT 0.0000 472.8000 3370.4200 474.4400 ;
      RECT 3368.7200 471.7200 3370.4200 472.8000 ;
      RECT 3305.0200 471.7200 3365.1200 472.8000 ;
      RECT 2497.4200 471.7200 3302.8200 472.8000 ;
      RECT 2446.4800 471.7200 2495.2200 472.8000 ;
      RECT 1007.4200 471.7200 2444.2800 472.8000 ;
      RECT 665.0200 471.7200 1005.2200 472.8000 ;
      RECT 507.4200 471.7200 662.8200 472.8000 ;
      RECT 5.3000 471.7200 505.2200 472.8000 ;
      RECT 0.0000 471.7200 1.7000 472.8000 ;
      RECT 0.0000 470.0800 3370.4200 471.7200 ;
      RECT 3364.7200 469.0000 3370.4200 470.0800 ;
      RECT 3307.6200 469.0000 3361.1200 470.0800 ;
      RECT 2494.8200 469.0000 3305.4200 470.0800 ;
      RECT 2449.0800 469.0000 2492.6200 470.0800 ;
      RECT 1004.8200 469.0000 2446.8800 470.0800 ;
      RECT 667.6200 469.0000 1002.6200 470.0800 ;
      RECT 504.8200 469.0000 665.4200 470.0800 ;
      RECT 9.3000 469.0000 502.6200 470.0800 ;
      RECT 0.0000 469.0000 5.7000 470.0800 ;
      RECT 0.0000 467.3600 3370.4200 469.0000 ;
      RECT 3368.7200 466.2800 3370.4200 467.3600 ;
      RECT 3305.0200 466.2800 3365.1200 467.3600 ;
      RECT 2497.4200 466.2800 3302.8200 467.3600 ;
      RECT 2446.4800 466.2800 2495.2200 467.3600 ;
      RECT 1007.4200 466.2800 2444.2800 467.3600 ;
      RECT 665.0200 466.2800 1005.2200 467.3600 ;
      RECT 507.4200 466.2800 662.8200 467.3600 ;
      RECT 5.3000 466.2800 505.2200 467.3600 ;
      RECT 0.0000 466.2800 1.7000 467.3600 ;
      RECT 0.0000 466.1500 3370.4200 466.2800 ;
      RECT 1.1000 465.2500 3370.4200 466.1500 ;
      RECT 0.0000 464.6400 3370.4200 465.2500 ;
      RECT 3364.7200 463.5600 3370.4200 464.6400 ;
      RECT 3307.6200 463.5600 3361.1200 464.6400 ;
      RECT 2494.8200 463.5600 3305.4200 464.6400 ;
      RECT 2449.0800 463.5600 2492.6200 464.6400 ;
      RECT 1004.8200 463.5600 2446.8800 464.6400 ;
      RECT 667.6200 463.5600 1002.6200 464.6400 ;
      RECT 504.8200 463.5600 665.4200 464.6400 ;
      RECT 9.3000 463.5600 502.6200 464.6400 ;
      RECT 0.0000 463.5600 5.7000 464.6400 ;
      RECT 0.0000 461.9200 3370.4200 463.5600 ;
      RECT 3368.7200 460.8400 3370.4200 461.9200 ;
      RECT 3305.0200 460.8400 3365.1200 461.9200 ;
      RECT 2497.4200 460.8400 3302.8200 461.9200 ;
      RECT 2446.4800 460.8400 2495.2200 461.9200 ;
      RECT 1007.4200 460.8400 2444.2800 461.9200 ;
      RECT 665.0200 460.8400 1005.2200 461.9200 ;
      RECT 507.4200 460.8400 662.8200 461.9200 ;
      RECT 5.3000 460.8400 505.2200 461.9200 ;
      RECT 0.0000 460.8400 1.7000 461.9200 ;
      RECT 0.0000 459.2000 3370.4200 460.8400 ;
      RECT 3364.7200 458.1200 3370.4200 459.2000 ;
      RECT 3307.6200 458.1200 3361.1200 459.2000 ;
      RECT 2494.8200 458.1200 3305.4200 459.2000 ;
      RECT 2449.0800 458.1200 2492.6200 459.2000 ;
      RECT 1004.8200 458.1200 2446.8800 459.2000 ;
      RECT 667.6200 458.1200 1002.6200 459.2000 ;
      RECT 504.8200 458.1200 665.4200 459.2000 ;
      RECT 9.3000 458.1200 502.6200 459.2000 ;
      RECT 0.0000 458.1200 5.7000 459.2000 ;
      RECT 0.0000 456.4800 3370.4200 458.1200 ;
      RECT 0.0000 455.7800 1.7000 456.4800 ;
      RECT 3368.7200 455.4000 3370.4200 456.4800 ;
      RECT 3305.0200 455.4000 3365.1200 456.4800 ;
      RECT 2497.4200 455.4000 3302.8200 456.4800 ;
      RECT 2446.4800 455.4000 2495.2200 456.4800 ;
      RECT 1007.4200 455.4000 2444.2800 456.4800 ;
      RECT 665.0200 455.4000 1005.2200 456.4800 ;
      RECT 507.4200 455.4000 662.8200 456.4800 ;
      RECT 5.3000 455.4000 505.2200 456.4800 ;
      RECT 1.1000 455.4000 1.7000 455.7800 ;
      RECT 1.1000 454.8800 3370.4200 455.4000 ;
      RECT 0.0000 453.7600 3370.4200 454.8800 ;
      RECT 3364.7200 452.6800 3370.4200 453.7600 ;
      RECT 3307.6200 452.6800 3361.1200 453.7600 ;
      RECT 2494.8200 452.6800 3305.4200 453.7600 ;
      RECT 2449.0800 452.6800 2492.6200 453.7600 ;
      RECT 1004.8200 452.6800 2446.8800 453.7600 ;
      RECT 667.6200 452.6800 1002.6200 453.7600 ;
      RECT 504.8200 452.6800 665.4200 453.7600 ;
      RECT 9.3000 452.6800 502.6200 453.7600 ;
      RECT 0.0000 452.6800 5.7000 453.7600 ;
      RECT 0.0000 451.0400 3370.4200 452.6800 ;
      RECT 3368.7200 449.9600 3370.4200 451.0400 ;
      RECT 3305.0200 449.9600 3365.1200 451.0400 ;
      RECT 2497.4200 449.9600 3302.8200 451.0400 ;
      RECT 2446.4800 449.9600 2495.2200 451.0400 ;
      RECT 1007.4200 449.9600 2444.2800 451.0400 ;
      RECT 665.0200 449.9600 1005.2200 451.0400 ;
      RECT 507.4200 449.9600 662.8200 451.0400 ;
      RECT 5.3000 449.9600 505.2200 451.0400 ;
      RECT 0.0000 449.9600 1.7000 451.0400 ;
      RECT 0.0000 448.3200 3370.4200 449.9600 ;
      RECT 3364.7200 447.2400 3370.4200 448.3200 ;
      RECT 3307.6200 447.2400 3361.1200 448.3200 ;
      RECT 2494.8200 447.2400 3305.4200 448.3200 ;
      RECT 2449.0800 447.2400 2492.6200 448.3200 ;
      RECT 1004.8200 447.2400 2446.8800 448.3200 ;
      RECT 667.6200 447.2400 1002.6200 448.3200 ;
      RECT 504.8200 447.2400 665.4200 448.3200 ;
      RECT 9.3000 447.2400 502.6200 448.3200 ;
      RECT 0.0000 447.2400 5.7000 448.3200 ;
      RECT 0.0000 445.6000 3370.4200 447.2400 ;
      RECT 0.0000 444.8000 1.7000 445.6000 ;
      RECT 3368.7200 444.5200 3370.4200 445.6000 ;
      RECT 3305.0200 444.5200 3365.1200 445.6000 ;
      RECT 2497.4200 444.5200 3302.8200 445.6000 ;
      RECT 2446.4800 444.5200 2495.2200 445.6000 ;
      RECT 1007.4200 444.5200 2444.2800 445.6000 ;
      RECT 665.0200 444.5200 1005.2200 445.6000 ;
      RECT 507.4200 444.5200 662.8200 445.6000 ;
      RECT 5.3000 444.5200 505.2200 445.6000 ;
      RECT 1.1000 444.5200 1.7000 444.8000 ;
      RECT 1.1000 443.9000 3370.4200 444.5200 ;
      RECT 0.0000 442.8800 3370.4200 443.9000 ;
      RECT 3364.7200 441.8000 3370.4200 442.8800 ;
      RECT 3307.6200 441.8000 3361.1200 442.8800 ;
      RECT 2494.8200 441.8000 3305.4200 442.8800 ;
      RECT 2449.0800 441.8000 2492.6200 442.8800 ;
      RECT 1004.8200 441.8000 2446.8800 442.8800 ;
      RECT 667.6200 441.8000 1002.6200 442.8800 ;
      RECT 504.8200 441.8000 665.4200 442.8800 ;
      RECT 9.3000 441.8000 502.6200 442.8800 ;
      RECT 0.0000 441.8000 5.7000 442.8800 ;
      RECT 0.0000 440.1600 3370.4200 441.8000 ;
      RECT 3368.7200 439.0800 3370.4200 440.1600 ;
      RECT 3305.0200 439.0800 3365.1200 440.1600 ;
      RECT 2497.4200 439.0800 3302.8200 440.1600 ;
      RECT 2446.4800 439.0800 2495.2200 440.1600 ;
      RECT 1007.4200 439.0800 2444.2800 440.1600 ;
      RECT 665.0200 439.0800 1005.2200 440.1600 ;
      RECT 507.4200 439.0800 662.8200 440.1600 ;
      RECT 5.3000 439.0800 505.2200 440.1600 ;
      RECT 0.0000 439.0800 1.7000 440.1600 ;
      RECT 0.0000 437.4400 3370.4200 439.0800 ;
      RECT 3364.7200 436.3600 3370.4200 437.4400 ;
      RECT 3307.6200 436.3600 3361.1200 437.4400 ;
      RECT 2494.8200 436.3600 3305.4200 437.4400 ;
      RECT 2449.0800 436.3600 2492.6200 437.4400 ;
      RECT 1004.8200 436.3600 2446.8800 437.4400 ;
      RECT 667.6200 436.3600 1002.6200 437.4400 ;
      RECT 504.8200 436.3600 665.4200 437.4400 ;
      RECT 9.3000 436.3600 502.6200 437.4400 ;
      RECT 0.0000 436.3600 5.7000 437.4400 ;
      RECT 0.0000 434.7200 3370.4200 436.3600 ;
      RECT 0.0000 433.8200 1.7000 434.7200 ;
      RECT 3368.7200 433.6400 3370.4200 434.7200 ;
      RECT 3305.0200 433.6400 3365.1200 434.7200 ;
      RECT 2497.4200 433.6400 3302.8200 434.7200 ;
      RECT 2446.4800 433.6400 2495.2200 434.7200 ;
      RECT 1007.4200 433.6400 2444.2800 434.7200 ;
      RECT 665.0200 433.6400 1005.2200 434.7200 ;
      RECT 507.4200 433.6400 662.8200 434.7200 ;
      RECT 5.3000 433.6400 505.2200 434.7200 ;
      RECT 1.1000 433.6400 1.7000 433.8200 ;
      RECT 1.1000 432.9200 3370.4200 433.6400 ;
      RECT 0.0000 432.0000 3370.4200 432.9200 ;
      RECT 3364.7200 430.9200 3370.4200 432.0000 ;
      RECT 3307.6200 430.9200 3361.1200 432.0000 ;
      RECT 2494.8200 430.9200 3305.4200 432.0000 ;
      RECT 2449.0800 430.9200 2492.6200 432.0000 ;
      RECT 1004.8200 430.9200 2446.8800 432.0000 ;
      RECT 667.6200 430.9200 1002.6200 432.0000 ;
      RECT 504.8200 430.9200 665.4200 432.0000 ;
      RECT 9.3000 430.9200 502.6200 432.0000 ;
      RECT 0.0000 430.9200 5.7000 432.0000 ;
      RECT 0.0000 429.2800 3370.4200 430.9200 ;
      RECT 3368.7200 428.2000 3370.4200 429.2800 ;
      RECT 3305.0200 428.2000 3365.1200 429.2800 ;
      RECT 2497.4200 428.2000 3302.8200 429.2800 ;
      RECT 2446.4800 428.2000 2495.2200 429.2800 ;
      RECT 1007.4200 428.2000 2444.2800 429.2800 ;
      RECT 665.0200 428.2000 1005.2200 429.2800 ;
      RECT 507.4200 428.2000 662.8200 429.2800 ;
      RECT 5.3000 428.2000 505.2200 429.2800 ;
      RECT 0.0000 428.2000 1.7000 429.2800 ;
      RECT 0.0000 426.5600 3370.4200 428.2000 ;
      RECT 3364.7200 425.4800 3370.4200 426.5600 ;
      RECT 3307.6200 425.4800 3361.1200 426.5600 ;
      RECT 2494.8200 425.4800 3305.4200 426.5600 ;
      RECT 2449.0800 425.4800 2492.6200 426.5600 ;
      RECT 1004.8200 425.4800 2446.8800 426.5600 ;
      RECT 667.6200 425.4800 1002.6200 426.5600 ;
      RECT 504.8200 425.4800 665.4200 426.5600 ;
      RECT 9.3000 425.4800 502.6200 426.5600 ;
      RECT 0.0000 425.4800 5.7000 426.5600 ;
      RECT 0.0000 423.8400 3370.4200 425.4800 ;
      RECT 1007.4200 423.5000 2444.2800 423.8400 ;
      RECT 1017.4800 423.2400 2444.2800 423.5000 ;
      RECT 0.0000 422.8400 1.7000 423.8400 ;
      RECT 3368.7200 422.7600 3370.4200 423.8400 ;
      RECT 3305.0200 422.7600 3365.1200 423.8400 ;
      RECT 2497.4200 422.7600 3302.8200 423.8400 ;
      RECT 2446.4800 422.7600 2495.2200 423.8400 ;
      RECT 2436.3200 422.7600 2444.2800 423.2400 ;
      RECT 1007.4200 422.7600 1015.2800 423.5000 ;
      RECT 665.0200 422.7600 1005.2200 423.8400 ;
      RECT 507.4200 422.7600 662.8200 423.8400 ;
      RECT 5.3000 422.7600 505.2200 423.8400 ;
      RECT 1.1000 422.7600 1.7000 422.8400 ;
      RECT 1017.4800 422.4200 1295.6000 423.2400 ;
      RECT 1.1000 422.4200 1015.2800 422.7600 ;
      RECT 2436.3200 422.1600 3370.4200 422.7600 ;
      RECT 2178.6800 422.1600 2434.1200 423.2400 ;
      RECT 1738.2400 422.1600 2176.4800 423.2400 ;
      RECT 1518.0200 422.1600 1736.0400 423.2400 ;
      RECT 1297.8000 422.1600 1515.8200 423.2400 ;
      RECT 1.1000 422.1600 1295.6000 422.4200 ;
      RECT 1.1000 421.9400 3370.4200 422.1600 ;
      RECT 0.0000 421.1200 3370.4200 421.9400 ;
      RECT 1004.8200 420.3300 2446.8800 421.1200 ;
      RECT 1065.1600 420.1700 2446.8800 420.3300 ;
      RECT 3364.7200 420.0400 3370.4200 421.1200 ;
      RECT 3307.6200 420.0400 3361.1200 421.1200 ;
      RECT 2494.8200 420.0400 3305.4200 421.1200 ;
      RECT 2449.0800 420.0400 2492.6200 421.1200 ;
      RECT 2446.4800 420.0400 2446.8800 420.1700 ;
      RECT 1004.8200 420.0400 1005.2200 420.3300 ;
      RECT 667.6200 420.0400 1002.6200 421.1200 ;
      RECT 504.8200 420.0400 665.4200 421.1200 ;
      RECT 9.3000 420.0400 502.6200 421.1200 ;
      RECT 0.0000 420.0400 5.7000 421.1200 ;
      RECT 2446.4800 418.4000 3370.4200 420.0400 ;
      RECT 0.0000 418.4000 1005.2200 420.0400 ;
      RECT 1065.1600 418.1300 1283.0400 420.1700 ;
      RECT 1011.2200 418.1300 1059.1600 420.3300 ;
      RECT 2392.5400 417.9700 2440.4800 420.1700 ;
      RECT 2172.3200 417.9700 2380.3400 420.1700 ;
      RECT 1945.9000 417.9700 2163.9200 420.1700 ;
      RECT 1731.8800 417.9700 1939.9000 420.1700 ;
      RECT 1511.6600 417.9700 1719.6800 420.1700 ;
      RECT 1291.4400 417.9700 1499.4600 420.1700 ;
      RECT 1007.4200 417.9700 1283.0400 418.1300 ;
      RECT 1007.4200 417.9300 2444.2800 417.9700 ;
      RECT 665.0200 417.9300 1005.2200 418.4000 ;
      RECT 2446.4800 417.5700 2495.2200 418.4000 ;
      RECT 1067.7600 417.5700 2444.2800 417.9300 ;
      RECT 3368.7200 417.3200 3370.4200 418.4000 ;
      RECT 3305.0200 417.3200 3365.1200 418.4000 ;
      RECT 2497.4200 417.3200 3302.8200 418.4000 ;
      RECT 2449.0800 417.3200 2495.2200 417.5700 ;
      RECT 665.0200 417.3200 1002.6200 417.9300 ;
      RECT 507.4200 417.3200 662.8200 418.4000 ;
      RECT 5.3000 417.3200 505.2200 418.4000 ;
      RECT 0.0000 417.3200 1.7000 418.4000 ;
      RECT 1067.7600 415.7300 1285.6400 417.5700 ;
      RECT 1011.2200 415.7300 1059.1600 417.9300 ;
      RECT 0.0000 415.7300 1002.6200 417.3200 ;
      RECT 2449.0800 415.6800 3370.4200 417.3200 ;
      RECT 0.0000 415.6800 1285.6400 415.7300 ;
      RECT 2449.0800 415.3700 2449.3400 415.6800 ;
      RECT 2392.5400 415.3700 2440.4800 417.5700 ;
      RECT 2172.3200 415.3700 2380.3400 417.5700 ;
      RECT 1948.5000 415.3700 2166.5200 417.5700 ;
      RECT 1731.8800 415.3700 1939.9000 417.5700 ;
      RECT 1511.6600 415.3700 1719.6800 417.5700 ;
      RECT 1291.4400 415.3700 1505.8600 417.5700 ;
      RECT 1004.8200 415.3700 1285.6400 415.6800 ;
      RECT 3364.7200 414.6000 3370.4200 415.6800 ;
      RECT 3307.6200 414.6000 3361.1200 415.6800 ;
      RECT 2494.8200 414.6000 3305.4200 415.6800 ;
      RECT 2450.4400 414.6000 2492.6200 415.6800 ;
      RECT 1004.8200 414.6000 2449.3400 415.3700 ;
      RECT 667.6200 414.6000 1002.6200 415.6800 ;
      RECT 504.8200 414.6000 665.4200 415.6800 ;
      RECT 9.3000 414.6000 502.6200 415.6800 ;
      RECT 0.0000 414.6000 5.7000 415.6800 ;
      RECT 0.0000 412.9600 3370.4200 414.6000 ;
      RECT 3368.7200 411.8800 3370.4200 412.9600 ;
      RECT 3305.0200 411.8800 3365.1200 412.9600 ;
      RECT 2497.4200 411.8800 3302.8200 412.9600 ;
      RECT 2446.4800 411.8800 2495.2200 412.9600 ;
      RECT 1007.4200 411.8800 2444.2800 412.9600 ;
      RECT 665.0200 411.8800 1005.2200 412.9600 ;
      RECT 507.4200 411.8800 662.8200 412.9600 ;
      RECT 5.3000 411.8800 505.2200 412.9600 ;
      RECT 0.0000 411.8800 1.7000 412.9600 ;
      RECT 0.0000 411.8600 3370.4200 411.8800 ;
      RECT 1.1000 411.3400 3370.4200 411.8600 ;
      RECT 1.1000 410.9600 5.7000 411.3400 ;
      RECT 1004.8200 410.4000 3370.4200 411.3400 ;
      RECT 667.6200 410.4000 1002.6200 411.3400 ;
      RECT 504.8200 410.4000 665.4200 411.3400 ;
      RECT 9.3000 410.4000 502.6200 411.3400 ;
      RECT 0.0000 410.4000 5.7000 410.9600 ;
      RECT 1065.1600 410.2400 3370.4200 410.4000 ;
      RECT 1065.1600 410.1400 2446.8800 410.2400 ;
      RECT 3364.7200 409.1600 3370.4200 410.2400 ;
      RECT 3307.6200 409.1600 3361.1200 410.2400 ;
      RECT 2494.8200 409.1600 3305.4200 410.2400 ;
      RECT 2449.0800 409.1600 2492.6200 410.2400 ;
      RECT 2446.4800 409.1600 2446.8800 410.1400 ;
      RECT 1065.1600 408.2000 1283.0400 410.1400 ;
      RECT 516.8150 408.2000 656.5450 410.4000 ;
      RECT 0.0000 408.2000 1.7000 410.4000 ;
      RECT 1945.9000 407.9400 2163.9200 410.1400 ;
      RECT 1007.4200 407.9400 1283.0400 408.2000 ;
      RECT 1007.4200 407.8200 2444.2800 407.9400 ;
      RECT 665.0200 407.8200 1005.2200 408.2000 ;
      RECT 507.4200 407.8200 662.8200 408.2000 ;
      RECT 0.0000 407.8200 505.2200 408.2000 ;
      RECT 0.0000 407.8000 2444.2800 407.8200 ;
      RECT 2446.4800 407.6300 3370.4200 409.1600 ;
      RECT 1067.7600 407.6300 2444.2800 407.8000 ;
      RECT 1067.7600 407.5400 3370.4200 407.6300 ;
      RECT 2449.0800 407.5200 3370.4200 407.5400 ;
      RECT 0.0000 407.5200 5.7000 407.8000 ;
      RECT 3368.7200 406.4400 3370.4200 407.5200 ;
      RECT 3305.0200 406.4400 3365.1200 407.5200 ;
      RECT 2497.4200 406.4400 3302.8200 407.5200 ;
      RECT 2449.0800 406.4400 2495.2200 407.5200 ;
      RECT 5.3000 406.4400 5.7000 407.5200 ;
      RECT 0.0000 406.4400 1.7000 407.5200 ;
      RECT 1067.7600 405.6000 1285.6400 407.5400 ;
      RECT 516.8150 405.6000 656.5450 407.8000 ;
      RECT 0.0000 405.6000 5.7000 406.4400 ;
      RECT 2449.0800 405.3400 3370.4200 406.4400 ;
      RECT 1948.5000 405.3400 2166.5200 407.5400 ;
      RECT 0.0000 405.3400 1285.6400 405.6000 ;
      RECT 0.0000 404.8000 3370.4200 405.3400 ;
      RECT 3364.7200 403.7200 3370.4200 404.8000 ;
      RECT 3307.6200 403.7200 3361.1200 404.8000 ;
      RECT 2494.8200 403.7200 3305.4200 404.8000 ;
      RECT 2449.0800 403.7200 2492.6200 404.8000 ;
      RECT 1004.8200 403.7200 2446.8800 404.8000 ;
      RECT 667.6200 403.7200 1002.6200 404.8000 ;
      RECT 504.8200 403.7200 665.4200 404.8000 ;
      RECT 9.3000 403.7200 502.6200 404.8000 ;
      RECT 0.0000 403.7200 5.7000 404.8000 ;
      RECT 0.0000 402.0800 3370.4200 403.7200 ;
      RECT 0.0000 401.4900 1.7000 402.0800 ;
      RECT 3368.7200 401.0000 3370.4200 402.0800 ;
      RECT 3305.0200 401.0000 3365.1200 402.0800 ;
      RECT 2497.4200 401.0000 3302.8200 402.0800 ;
      RECT 2446.4800 401.0000 2495.2200 402.0800 ;
      RECT 1007.4200 401.0000 2444.2800 402.0800 ;
      RECT 665.0200 401.0000 1005.2200 402.0800 ;
      RECT 507.4200 401.0000 662.8200 402.0800 ;
      RECT 5.3000 401.0000 505.2200 402.0800 ;
      RECT 1.1000 401.0000 1.7000 401.4900 ;
      RECT 1.1000 400.5900 3370.4200 401.0000 ;
      RECT 0.0000 399.7900 3370.4200 400.5900 ;
      RECT 1067.7600 399.6300 3370.4200 399.7900 ;
      RECT 2449.0800 399.3600 3370.4200 399.6300 ;
      RECT 0.0000 399.3600 1002.6200 399.7900 ;
      RECT 3364.7200 398.2800 3370.4200 399.3600 ;
      RECT 3307.6200 398.2800 3361.1200 399.3600 ;
      RECT 2494.8200 398.2800 3305.4200 399.3600 ;
      RECT 2449.0800 398.2800 2492.6200 399.3600 ;
      RECT 667.6200 398.2800 1002.6200 399.3600 ;
      RECT 504.8200 398.2800 665.4200 399.3600 ;
      RECT 9.3000 398.2800 502.6200 399.3600 ;
      RECT 0.0000 398.2800 5.7000 399.3600 ;
      RECT 1067.7600 397.5900 1285.6400 399.6300 ;
      RECT 1011.2200 397.5900 1059.1600 399.7900 ;
      RECT 0.0000 397.5900 1002.6200 398.2800 ;
      RECT 2449.0800 397.4300 3370.4200 398.2800 ;
      RECT 2392.5400 397.4300 2440.4800 399.6300 ;
      RECT 2172.3200 397.4300 2380.3400 399.6300 ;
      RECT 1948.5000 397.4300 2166.5200 399.6300 ;
      RECT 1731.8800 397.4300 1939.9000 399.6300 ;
      RECT 1511.6600 397.4300 1719.6800 399.6300 ;
      RECT 1291.4400 397.4300 1499.4600 399.6300 ;
      RECT 0.0000 397.4300 1285.6400 397.5900 ;
      RECT 0.0000 397.3900 3370.4200 397.4300 ;
      RECT 1065.1600 397.0300 3370.4200 397.3900 ;
      RECT 2446.4800 396.6400 3370.4200 397.0300 ;
      RECT 0.0000 396.6400 1005.2200 397.3900 ;
      RECT 3368.7200 395.5600 3370.4200 396.6400 ;
      RECT 3305.0200 395.5600 3365.1200 396.6400 ;
      RECT 2497.4200 395.5600 3302.8200 396.6400 ;
      RECT 2446.4800 395.5600 2495.2200 396.6400 ;
      RECT 665.0200 395.5600 1005.2200 396.6400 ;
      RECT 507.4200 395.5600 662.8200 396.6400 ;
      RECT 5.3000 395.5600 505.2200 396.6400 ;
      RECT 0.0000 395.5600 1.7000 396.6400 ;
      RECT 1065.1600 395.1900 1283.0400 397.0300 ;
      RECT 1011.2200 395.1900 1059.1600 397.3900 ;
      RECT 0.0000 395.1900 1005.2200 395.5600 ;
      RECT 2446.4800 394.8300 3370.4200 395.5600 ;
      RECT 2392.5400 394.8300 2440.4800 397.0300 ;
      RECT 2172.3200 394.8300 2380.3400 397.0300 ;
      RECT 1945.9000 394.8300 2163.9200 397.0300 ;
      RECT 1731.8800 394.8300 1939.9000 397.0300 ;
      RECT 1511.6600 394.8300 1719.6800 397.0300 ;
      RECT 1291.4400 394.8300 1499.4600 397.0300 ;
      RECT 0.0000 394.8300 1283.0400 395.1900 ;
      RECT 0.0000 393.9200 3370.4200 394.8300 ;
      RECT 3364.7200 392.8400 3370.4200 393.9200 ;
      RECT 3307.6200 392.8400 3361.1200 393.9200 ;
      RECT 2494.8200 392.8400 3305.4200 393.9200 ;
      RECT 2449.0800 392.8400 2492.6200 393.9200 ;
      RECT 1004.8200 392.8400 2446.8800 393.9200 ;
      RECT 667.6200 392.8400 1002.6200 393.9200 ;
      RECT 504.8200 392.8400 665.4200 393.9200 ;
      RECT 9.3000 392.8400 502.6200 393.9200 ;
      RECT 0.0000 392.8400 5.7000 393.9200 ;
      RECT 0.0000 392.4200 3370.4200 392.8400 ;
      RECT 1015.0800 392.1600 3370.4200 392.4200 ;
      RECT 1015.0800 391.3400 1293.0000 392.1600 ;
      RECT 0.0000 391.3400 1012.8800 392.4200 ;
      RECT 2396.3000 391.2000 3370.4200 392.1600 ;
      RECT 0.0000 391.2000 1293.0000 391.3400 ;
      RECT 2396.3000 391.0800 2444.2800 391.2000 ;
      RECT 2176.0800 391.0800 2394.1000 392.1600 ;
      RECT 1735.6400 391.0800 2173.8800 392.1600 ;
      RECT 1515.4200 391.0800 1733.4400 392.1600 ;
      RECT 1295.2000 391.0800 1513.2200 392.1600 ;
      RECT 1007.4200 391.0800 1293.0000 391.2000 ;
      RECT 0.0000 390.5100 1.7000 391.2000 ;
      RECT 3368.7200 390.1200 3370.4200 391.2000 ;
      RECT 3305.0200 390.1200 3365.1200 391.2000 ;
      RECT 2497.4200 390.1200 3302.8200 391.2000 ;
      RECT 2446.4800 390.1200 2495.2200 391.2000 ;
      RECT 1007.4200 390.1200 2444.2800 391.0800 ;
      RECT 665.0200 390.1200 1005.2200 391.2000 ;
      RECT 507.4200 390.1200 662.8200 391.2000 ;
      RECT 5.3000 390.1200 505.2200 391.2000 ;
      RECT 1.1000 390.1200 1.7000 390.5100 ;
      RECT 1.1000 389.6100 3370.4200 390.1200 ;
      RECT 0.0000 388.4800 3370.4200 389.6100 ;
      RECT 3364.7200 387.4000 3370.4200 388.4800 ;
      RECT 3307.6200 387.4000 3361.1200 388.4800 ;
      RECT 2494.8200 387.4000 3305.4200 388.4800 ;
      RECT 2449.0800 387.4000 2492.6200 388.4800 ;
      RECT 1004.8200 387.4000 2446.8800 388.4800 ;
      RECT 667.6200 387.4000 1002.6200 388.4800 ;
      RECT 504.8200 387.4000 665.4200 388.4800 ;
      RECT 9.3000 387.4000 502.6200 388.4800 ;
      RECT 0.0000 387.4000 5.7000 388.4800 ;
      RECT 0.0000 385.7600 3370.4200 387.4000 ;
      RECT 3368.7200 384.6800 3370.4200 385.7600 ;
      RECT 3305.0200 384.6800 3365.1200 385.7600 ;
      RECT 2497.4200 384.6800 3302.8200 385.7600 ;
      RECT 2446.4800 384.6800 2495.2200 385.7600 ;
      RECT 1007.4200 384.6800 2444.2800 385.7600 ;
      RECT 665.0200 384.6800 1005.2200 385.7600 ;
      RECT 507.4200 384.6800 662.8200 385.7600 ;
      RECT 5.3000 384.6800 505.2200 385.7600 ;
      RECT 0.0000 384.6800 1.7000 385.7600 ;
      RECT 0.0000 383.0400 3370.4200 384.6800 ;
      RECT 3364.7200 381.9600 3370.4200 383.0400 ;
      RECT 3307.6200 381.9600 3361.1200 383.0400 ;
      RECT 2494.8200 381.9600 3305.4200 383.0400 ;
      RECT 2449.0800 381.9600 2492.6200 383.0400 ;
      RECT 1004.8200 381.9600 2446.8800 383.0400 ;
      RECT 667.6200 381.9600 1002.6200 383.0400 ;
      RECT 504.8200 381.9600 665.4200 383.0400 ;
      RECT 9.3000 381.9600 502.6200 383.0400 ;
      RECT 0.0000 381.9600 5.7000 383.0400 ;
      RECT 0.0000 380.3200 3370.4200 381.9600 ;
      RECT 0.0000 379.5300 1.7000 380.3200 ;
      RECT 3368.7200 379.2400 3370.4200 380.3200 ;
      RECT 3305.0200 379.2400 3365.1200 380.3200 ;
      RECT 2497.4200 379.2400 3302.8200 380.3200 ;
      RECT 2446.4800 379.2400 2495.2200 380.3200 ;
      RECT 1007.4200 379.2400 2444.2800 380.3200 ;
      RECT 665.0200 379.2400 1005.2200 380.3200 ;
      RECT 507.4200 379.2400 662.8200 380.3200 ;
      RECT 5.3000 379.2400 505.2200 380.3200 ;
      RECT 1.1000 379.2400 1.7000 379.5300 ;
      RECT 1.1000 378.6300 3370.4200 379.2400 ;
      RECT 0.0000 377.6000 3370.4200 378.6300 ;
      RECT 3364.7200 376.5200 3370.4200 377.6000 ;
      RECT 3307.6200 376.5200 3361.1200 377.6000 ;
      RECT 2494.8200 376.5200 3305.4200 377.6000 ;
      RECT 2449.0800 376.5200 2492.6200 377.6000 ;
      RECT 1004.8200 376.5200 2446.8800 377.6000 ;
      RECT 667.6200 376.5200 1002.6200 377.6000 ;
      RECT 504.8200 376.5200 665.4200 377.6000 ;
      RECT 9.3000 376.5200 502.6200 377.6000 ;
      RECT 0.0000 376.5200 5.7000 377.6000 ;
      RECT 0.0000 374.8800 3370.4200 376.5200 ;
      RECT 3368.7200 373.8000 3370.4200 374.8800 ;
      RECT 3305.0200 373.8000 3365.1200 374.8800 ;
      RECT 2497.4200 373.8000 3302.8200 374.8800 ;
      RECT 2446.4800 373.8000 2495.2200 374.8800 ;
      RECT 1007.4200 373.8000 2444.2800 374.8800 ;
      RECT 665.0200 373.8000 1005.2200 374.8800 ;
      RECT 507.4200 373.8000 662.8200 374.8800 ;
      RECT 5.3000 373.8000 505.2200 374.8800 ;
      RECT 0.0000 373.8000 1.7000 374.8800 ;
      RECT 0.0000 372.1600 3370.4200 373.8000 ;
      RECT 3364.7200 371.0800 3370.4200 372.1600 ;
      RECT 3307.6200 371.0800 3361.1200 372.1600 ;
      RECT 2494.8200 371.0800 3305.4200 372.1600 ;
      RECT 2449.0800 371.0800 2492.6200 372.1600 ;
      RECT 1004.8200 371.0800 2446.8800 372.1600 ;
      RECT 667.6200 371.0800 1002.6200 372.1600 ;
      RECT 504.8200 371.0800 665.4200 372.1600 ;
      RECT 9.3000 371.0800 502.6200 372.1600 ;
      RECT 0.0000 371.0800 5.7000 372.1600 ;
      RECT 0.0000 369.4400 3370.4200 371.0800 ;
      RECT 0.0000 368.5500 1.7000 369.4400 ;
      RECT 3368.7200 368.3600 3370.4200 369.4400 ;
      RECT 3305.0200 368.3600 3365.1200 369.4400 ;
      RECT 2497.4200 368.3600 3302.8200 369.4400 ;
      RECT 2446.4800 368.3600 2495.2200 369.4400 ;
      RECT 1007.4200 368.3600 2444.2800 369.4400 ;
      RECT 665.0200 368.3600 1005.2200 369.4400 ;
      RECT 507.4200 368.3600 662.8200 369.4400 ;
      RECT 5.3000 368.3600 505.2200 369.4400 ;
      RECT 1.1000 368.3600 1.7000 368.5500 ;
      RECT 1.1000 367.6500 3370.4200 368.3600 ;
      RECT 0.0000 366.7200 3370.4200 367.6500 ;
      RECT 3364.7200 365.6400 3370.4200 366.7200 ;
      RECT 3307.6200 365.6400 3361.1200 366.7200 ;
      RECT 2494.8200 365.6400 3305.4200 366.7200 ;
      RECT 2449.0800 365.6400 2492.6200 366.7200 ;
      RECT 1004.8200 365.6400 2446.8800 366.7200 ;
      RECT 667.6200 365.6400 1002.6200 366.7200 ;
      RECT 504.8200 365.6400 665.4200 366.7200 ;
      RECT 9.3000 365.6400 502.6200 366.7200 ;
      RECT 0.0000 365.6400 5.7000 366.7200 ;
      RECT 0.0000 364.0000 3370.4200 365.6400 ;
      RECT 3368.7200 362.9200 3370.4200 364.0000 ;
      RECT 3305.0200 362.9200 3365.1200 364.0000 ;
      RECT 2497.4200 362.9200 3302.8200 364.0000 ;
      RECT 2446.4800 362.9200 2495.2200 364.0000 ;
      RECT 1007.4200 362.9200 2444.2800 364.0000 ;
      RECT 665.0200 362.9200 1005.2200 364.0000 ;
      RECT 507.4200 362.9200 662.8200 364.0000 ;
      RECT 5.3000 362.9200 505.2200 364.0000 ;
      RECT 0.0000 362.9200 1.7000 364.0000 ;
      RECT 0.0000 361.2800 3370.4200 362.9200 ;
      RECT 3364.7200 360.2000 3370.4200 361.2800 ;
      RECT 3307.6200 360.2000 3361.1200 361.2800 ;
      RECT 2494.8200 360.2000 3305.4200 361.2800 ;
      RECT 2449.0800 360.2000 2492.6200 361.2800 ;
      RECT 1004.8200 360.2000 2446.8800 361.2800 ;
      RECT 667.6200 360.2000 1002.6200 361.2800 ;
      RECT 504.8200 360.2000 665.4200 361.2800 ;
      RECT 9.3000 360.2000 502.6200 361.2800 ;
      RECT 0.0000 360.2000 5.7000 361.2800 ;
      RECT 0.0000 358.5600 3370.4200 360.2000 ;
      RECT 0.0000 357.5700 1.7000 358.5600 ;
      RECT 3368.7200 357.4800 3370.4200 358.5600 ;
      RECT 3305.0200 357.4800 3365.1200 358.5600 ;
      RECT 2497.4200 357.4800 3302.8200 358.5600 ;
      RECT 2446.4800 357.4800 2495.2200 358.5600 ;
      RECT 1007.4200 357.4800 2444.2800 358.5600 ;
      RECT 665.0200 357.4800 1005.2200 358.5600 ;
      RECT 507.4200 357.4800 662.8200 358.5600 ;
      RECT 5.3000 357.4800 505.2200 358.5600 ;
      RECT 1.1000 357.4800 1.7000 357.5700 ;
      RECT 1.1000 356.6700 3370.4200 357.4800 ;
      RECT 0.0000 355.8400 3370.4200 356.6700 ;
      RECT 3364.7200 354.7600 3370.4200 355.8400 ;
      RECT 3307.6200 354.7600 3361.1200 355.8400 ;
      RECT 2494.8200 354.7600 3305.4200 355.8400 ;
      RECT 2449.0800 354.7600 2492.6200 355.8400 ;
      RECT 1004.8200 354.7600 2446.8800 355.8400 ;
      RECT 667.6200 354.7600 1002.6200 355.8400 ;
      RECT 504.8200 354.7600 665.4200 355.8400 ;
      RECT 9.3000 354.7600 502.6200 355.8400 ;
      RECT 0.0000 354.7600 5.7000 355.8400 ;
      RECT 0.0000 353.1200 3370.4200 354.7600 ;
      RECT 3368.7200 352.0400 3370.4200 353.1200 ;
      RECT 3305.0200 352.0400 3365.1200 353.1200 ;
      RECT 2497.4200 352.0400 3302.8200 353.1200 ;
      RECT 2446.4800 352.0400 2495.2200 353.1200 ;
      RECT 1007.4200 352.0400 2444.2800 353.1200 ;
      RECT 665.0200 352.0400 1005.2200 353.1200 ;
      RECT 507.4200 352.0400 662.8200 353.1200 ;
      RECT 5.3000 352.0400 505.2200 353.1200 ;
      RECT 0.0000 352.0400 1.7000 353.1200 ;
      RECT 0.0000 350.4000 3370.4200 352.0400 ;
      RECT 3364.7200 349.3200 3370.4200 350.4000 ;
      RECT 3307.6200 349.3200 3361.1200 350.4000 ;
      RECT 2494.8200 349.3200 3305.4200 350.4000 ;
      RECT 2449.0800 349.3200 2492.6200 350.4000 ;
      RECT 1004.8200 349.3200 2446.8800 350.4000 ;
      RECT 667.6200 349.3200 1002.6200 350.4000 ;
      RECT 504.8200 349.3200 665.4200 350.4000 ;
      RECT 9.3000 349.3200 502.6200 350.4000 ;
      RECT 0.0000 349.3200 5.7000 350.4000 ;
      RECT 0.0000 347.6800 3370.4200 349.3200 ;
      RECT 0.0000 347.2000 1.7000 347.6800 ;
      RECT 3368.7200 346.6000 3370.4200 347.6800 ;
      RECT 3305.0200 346.6000 3365.1200 347.6800 ;
      RECT 2497.4200 346.6000 3302.8200 347.6800 ;
      RECT 2446.4800 346.6000 2495.2200 347.6800 ;
      RECT 1007.4200 346.6000 2444.2800 347.6800 ;
      RECT 665.0200 346.6000 1005.2200 347.6800 ;
      RECT 507.4200 346.6000 662.8200 347.6800 ;
      RECT 5.3000 346.6000 505.2200 347.6800 ;
      RECT 1.1000 346.6000 1.7000 347.2000 ;
      RECT 1.1000 346.3000 3370.4200 346.6000 ;
      RECT 0.0000 344.9600 3370.4200 346.3000 ;
      RECT 3364.7200 343.8800 3370.4200 344.9600 ;
      RECT 3307.6200 343.8800 3361.1200 344.9600 ;
      RECT 2494.8200 343.8800 3305.4200 344.9600 ;
      RECT 2449.0800 343.8800 2492.6200 344.9600 ;
      RECT 1004.8200 343.8800 2446.8800 344.9600 ;
      RECT 667.6200 343.8800 1002.6200 344.9600 ;
      RECT 504.8200 343.8800 665.4200 344.9600 ;
      RECT 9.3000 343.8800 502.6200 344.9600 ;
      RECT 0.0000 343.8800 5.7000 344.9600 ;
      RECT 0.0000 342.2400 3370.4200 343.8800 ;
      RECT 3368.7200 341.1600 3370.4200 342.2400 ;
      RECT 3305.0200 341.1600 3365.1200 342.2400 ;
      RECT 2497.4200 341.1600 3302.8200 342.2400 ;
      RECT 2446.4800 341.1600 2495.2200 342.2400 ;
      RECT 1007.4200 341.1600 2444.2800 342.2400 ;
      RECT 665.0200 341.1600 1005.2200 342.2400 ;
      RECT 507.4200 341.1600 662.8200 342.2400 ;
      RECT 5.3000 341.1600 505.2200 342.2400 ;
      RECT 0.0000 341.1600 1.7000 342.2400 ;
      RECT 0.0000 339.5200 3370.4200 341.1600 ;
      RECT 3364.7200 338.4400 3370.4200 339.5200 ;
      RECT 3307.6200 338.4400 3361.1200 339.5200 ;
      RECT 2494.8200 338.4400 3305.4200 339.5200 ;
      RECT 2449.0800 338.4400 2492.6200 339.5200 ;
      RECT 1004.8200 338.4400 2446.8800 339.5200 ;
      RECT 667.6200 338.4400 1002.6200 339.5200 ;
      RECT 504.8200 338.4400 665.4200 339.5200 ;
      RECT 9.3000 338.4400 502.6200 339.5200 ;
      RECT 0.0000 338.4400 5.7000 339.5200 ;
      RECT 0.0000 336.8000 3370.4200 338.4400 ;
      RECT 0.0000 336.2200 1.7000 336.8000 ;
      RECT 3368.7200 335.7200 3370.4200 336.8000 ;
      RECT 3305.0200 335.7200 3365.1200 336.8000 ;
      RECT 2497.4200 335.7200 3302.8200 336.8000 ;
      RECT 2446.4800 335.7200 2495.2200 336.8000 ;
      RECT 1007.4200 335.7200 2444.2800 336.8000 ;
      RECT 665.0200 335.7200 1005.2200 336.8000 ;
      RECT 507.4200 335.7200 662.8200 336.8000 ;
      RECT 5.3000 335.7200 505.2200 336.8000 ;
      RECT 1.1000 335.7200 1.7000 336.2200 ;
      RECT 1.1000 335.3200 3370.4200 335.7200 ;
      RECT 0.0000 334.0800 3370.4200 335.3200 ;
      RECT 3364.7200 333.0000 3370.4200 334.0800 ;
      RECT 3307.6200 333.0000 3361.1200 334.0800 ;
      RECT 2494.8200 333.0000 3305.4200 334.0800 ;
      RECT 2449.0800 333.0000 2492.6200 334.0800 ;
      RECT 1004.8200 333.0000 2446.8800 334.0800 ;
      RECT 667.6200 333.0000 1002.6200 334.0800 ;
      RECT 504.8200 333.0000 665.4200 334.0800 ;
      RECT 9.3000 333.0000 502.6200 334.0800 ;
      RECT 0.0000 333.0000 5.7000 334.0800 ;
      RECT 0.0000 331.3600 3370.4200 333.0000 ;
      RECT 3368.7200 330.2800 3370.4200 331.3600 ;
      RECT 3305.0200 330.2800 3365.1200 331.3600 ;
      RECT 2497.4200 330.2800 3302.8200 331.3600 ;
      RECT 2446.4800 330.2800 2495.2200 331.3600 ;
      RECT 1007.4200 330.2800 2444.2800 331.3600 ;
      RECT 665.0200 330.2800 1005.2200 331.3600 ;
      RECT 507.4200 330.2800 662.8200 331.3600 ;
      RECT 5.3000 330.2800 505.2200 331.3600 ;
      RECT 0.0000 330.2800 1.7000 331.3600 ;
      RECT 0.0000 328.6400 3370.4200 330.2800 ;
      RECT 3364.7200 327.5600 3370.4200 328.6400 ;
      RECT 3307.6200 327.5600 3361.1200 328.6400 ;
      RECT 2494.8200 327.5600 3305.4200 328.6400 ;
      RECT 2449.0800 327.5600 2492.6200 328.6400 ;
      RECT 1004.8200 327.5600 2446.8800 328.6400 ;
      RECT 667.6200 327.5600 1002.6200 328.6400 ;
      RECT 504.8200 327.5600 665.4200 328.6400 ;
      RECT 9.3000 327.5600 502.6200 328.6400 ;
      RECT 0.0000 327.5600 5.7000 328.6400 ;
      RECT 0.0000 325.9200 3370.4200 327.5600 ;
      RECT 0.0000 325.2400 1.7000 325.9200 ;
      RECT 3368.7200 324.8400 3370.4200 325.9200 ;
      RECT 3305.0200 324.8400 3365.1200 325.9200 ;
      RECT 2497.4200 324.8400 3302.8200 325.9200 ;
      RECT 2446.4800 324.8400 2495.2200 325.9200 ;
      RECT 1007.4200 324.8400 2444.2800 325.9200 ;
      RECT 665.0200 324.8400 1005.2200 325.9200 ;
      RECT 507.4200 324.8400 662.8200 325.9200 ;
      RECT 5.3000 324.8400 505.2200 325.9200 ;
      RECT 1.1000 324.8400 1.7000 325.2400 ;
      RECT 1.1000 324.3400 3370.4200 324.8400 ;
      RECT 0.0000 323.2000 3370.4200 324.3400 ;
      RECT 3364.7200 322.1200 3370.4200 323.2000 ;
      RECT 3307.6200 322.1200 3361.1200 323.2000 ;
      RECT 2494.8200 322.1200 3305.4200 323.2000 ;
      RECT 2449.0800 322.1200 2492.6200 323.2000 ;
      RECT 1004.8200 322.1200 2446.8800 323.2000 ;
      RECT 667.6200 322.1200 1002.6200 323.2000 ;
      RECT 504.8200 322.1200 665.4200 323.2000 ;
      RECT 9.3000 322.1200 502.6200 323.2000 ;
      RECT 0.0000 322.1200 5.7000 323.2000 ;
      RECT 0.0000 320.4800 3370.4200 322.1200 ;
      RECT 3368.7200 319.4000 3370.4200 320.4800 ;
      RECT 3305.0200 319.4000 3365.1200 320.4800 ;
      RECT 2497.4200 319.4000 3302.8200 320.4800 ;
      RECT 2446.4800 319.4000 2495.2200 320.4800 ;
      RECT 1007.4200 319.4000 2444.2800 320.4800 ;
      RECT 665.0200 319.4000 1005.2200 320.4800 ;
      RECT 507.4200 319.4000 662.8200 320.4800 ;
      RECT 5.3000 319.4000 505.2200 320.4800 ;
      RECT 0.0000 319.4000 1.7000 320.4800 ;
      RECT 0.0000 317.7600 3370.4200 319.4000 ;
      RECT 3364.7200 316.6800 3370.4200 317.7600 ;
      RECT 3307.6200 316.6800 3361.1200 317.7600 ;
      RECT 2494.8200 316.6800 3305.4200 317.7600 ;
      RECT 2449.0800 316.6800 2492.6200 317.7600 ;
      RECT 1004.8200 316.6800 2446.8800 317.7600 ;
      RECT 667.6200 316.6800 1002.6200 317.7600 ;
      RECT 504.8200 316.6800 665.4200 317.7600 ;
      RECT 9.3000 316.6800 502.6200 317.7600 ;
      RECT 0.0000 316.6800 5.7000 317.7600 ;
      RECT 0.0000 315.0400 3370.4200 316.6800 ;
      RECT 0.0000 314.2600 1.7000 315.0400 ;
      RECT 3368.7200 313.9600 3370.4200 315.0400 ;
      RECT 3305.0200 313.9600 3365.1200 315.0400 ;
      RECT 2497.4200 313.9600 3302.8200 315.0400 ;
      RECT 2446.4800 313.9600 2495.2200 315.0400 ;
      RECT 1007.4200 313.9600 2444.2800 315.0400 ;
      RECT 665.0200 313.9600 1005.2200 315.0400 ;
      RECT 507.4200 313.9600 662.8200 315.0400 ;
      RECT 5.3000 313.9600 505.2200 315.0400 ;
      RECT 1.1000 313.9600 1.7000 314.2600 ;
      RECT 1.1000 313.3600 3370.4200 313.9600 ;
      RECT 0.0000 312.3200 3370.4200 313.3600 ;
      RECT 3364.7200 311.2400 3370.4200 312.3200 ;
      RECT 3307.6200 311.2400 3361.1200 312.3200 ;
      RECT 2494.8200 311.2400 3305.4200 312.3200 ;
      RECT 2449.0800 311.2400 2492.6200 312.3200 ;
      RECT 1004.8200 311.2400 2446.8800 312.3200 ;
      RECT 667.6200 311.2400 1002.6200 312.3200 ;
      RECT 504.8200 311.2400 665.4200 312.3200 ;
      RECT 9.3000 311.2400 502.6200 312.3200 ;
      RECT 0.0000 311.2400 5.7000 312.3200 ;
      RECT 0.0000 309.6000 3370.4200 311.2400 ;
      RECT 3368.7200 308.5200 3370.4200 309.6000 ;
      RECT 3305.0200 308.5200 3365.1200 309.6000 ;
      RECT 2497.4200 308.5200 3302.8200 309.6000 ;
      RECT 2446.4800 308.5200 2495.2200 309.6000 ;
      RECT 1007.4200 308.5200 2444.2800 309.6000 ;
      RECT 665.0200 308.5200 1005.2200 309.6000 ;
      RECT 507.4200 308.5200 662.8200 309.6000 ;
      RECT 5.3000 308.5200 505.2200 309.6000 ;
      RECT 0.0000 308.5200 1.7000 309.6000 ;
      RECT 0.0000 306.8800 3370.4200 308.5200 ;
      RECT 3364.7200 305.8000 3370.4200 306.8800 ;
      RECT 3307.6200 305.8000 3361.1200 306.8800 ;
      RECT 2494.8200 305.8000 3305.4200 306.8800 ;
      RECT 2449.0800 305.8000 2492.6200 306.8800 ;
      RECT 1004.8200 305.8000 2446.8800 306.8800 ;
      RECT 667.6200 305.8000 1002.6200 306.8800 ;
      RECT 504.8200 305.8000 665.4200 306.8800 ;
      RECT 9.3000 305.8000 502.6200 306.8800 ;
      RECT 0.0000 305.8000 5.7000 306.8800 ;
      RECT 0.0000 304.1600 3370.4200 305.8000 ;
      RECT 0.0000 303.2800 1.7000 304.1600 ;
      RECT 3368.7200 303.0800 3370.4200 304.1600 ;
      RECT 3305.0200 303.0800 3365.1200 304.1600 ;
      RECT 2497.4200 303.0800 3302.8200 304.1600 ;
      RECT 2446.4800 303.0800 2495.2200 304.1600 ;
      RECT 1007.4200 303.0800 2444.2800 304.1600 ;
      RECT 665.0200 303.0800 1005.2200 304.1600 ;
      RECT 507.4200 303.0800 662.8200 304.1600 ;
      RECT 5.3000 303.0800 505.2200 304.1600 ;
      RECT 1.1000 303.0800 1.7000 303.2800 ;
      RECT 1.1000 302.3800 3370.4200 303.0800 ;
      RECT 0.0000 301.4400 3370.4200 302.3800 ;
      RECT 3364.7200 300.3600 3370.4200 301.4400 ;
      RECT 3307.6200 300.3600 3361.1200 301.4400 ;
      RECT 2494.8200 300.3600 3305.4200 301.4400 ;
      RECT 2449.0800 300.3600 2492.6200 301.4400 ;
      RECT 1004.8200 300.3600 2446.8800 301.4400 ;
      RECT 667.6200 300.3600 1002.6200 301.4400 ;
      RECT 504.8200 300.3600 665.4200 301.4400 ;
      RECT 9.3000 300.3600 502.6200 301.4400 ;
      RECT 0.0000 300.3600 5.7000 301.4400 ;
      RECT 0.0000 298.7200 3370.4200 300.3600 ;
      RECT 3368.7200 297.6400 3370.4200 298.7200 ;
      RECT 3305.0200 297.6400 3365.1200 298.7200 ;
      RECT 2497.4200 297.6400 3302.8200 298.7200 ;
      RECT 2446.4800 297.6400 2495.2200 298.7200 ;
      RECT 1007.4200 297.6400 2444.2800 298.7200 ;
      RECT 665.0200 297.6400 1005.2200 298.7200 ;
      RECT 507.4200 297.6400 662.8200 298.7200 ;
      RECT 5.3000 297.6400 505.2200 298.7200 ;
      RECT 0.0000 297.6400 1.7000 298.7200 ;
      RECT 0.0000 296.0000 3370.4200 297.6400 ;
      RECT 3364.7200 294.9200 3370.4200 296.0000 ;
      RECT 3307.6200 294.9200 3361.1200 296.0000 ;
      RECT 2494.8200 294.9200 3305.4200 296.0000 ;
      RECT 2449.0800 294.9200 2492.6200 296.0000 ;
      RECT 1004.8200 294.9200 2446.8800 296.0000 ;
      RECT 667.6200 294.9200 1002.6200 296.0000 ;
      RECT 504.8200 294.9200 665.4200 296.0000 ;
      RECT 9.3000 294.9200 502.6200 296.0000 ;
      RECT 0.0000 294.9200 5.7000 296.0000 ;
      RECT 0.0000 293.2800 3370.4200 294.9200 ;
      RECT 0.0000 292.9100 1.7000 293.2800 ;
      RECT 3368.7200 292.2000 3370.4200 293.2800 ;
      RECT 3305.0200 292.2000 3365.1200 293.2800 ;
      RECT 2497.4200 292.2000 3302.8200 293.2800 ;
      RECT 2446.4800 292.2000 2495.2200 293.2800 ;
      RECT 1007.4200 292.2000 2444.2800 293.2800 ;
      RECT 665.0200 292.2000 1005.2200 293.2800 ;
      RECT 507.4200 292.2000 662.8200 293.2800 ;
      RECT 5.3000 292.2000 505.2200 293.2800 ;
      RECT 1.1000 292.2000 1.7000 292.9100 ;
      RECT 1.1000 292.0100 3370.4200 292.2000 ;
      RECT 0.0000 290.5600 3370.4200 292.0100 ;
      RECT 3364.7200 289.4800 3370.4200 290.5600 ;
      RECT 3307.6200 289.4800 3361.1200 290.5600 ;
      RECT 2494.8200 289.4800 3305.4200 290.5600 ;
      RECT 2449.0800 289.4800 2492.6200 290.5600 ;
      RECT 1004.8200 289.4800 2446.8800 290.5600 ;
      RECT 667.6200 289.4800 1002.6200 290.5600 ;
      RECT 504.8200 289.4800 665.4200 290.5600 ;
      RECT 9.3000 289.4800 502.6200 290.5600 ;
      RECT 0.0000 289.4800 5.7000 290.5600 ;
      RECT 0.0000 287.8400 3370.4200 289.4800 ;
      RECT 3368.7200 286.7600 3370.4200 287.8400 ;
      RECT 3305.0200 286.7600 3365.1200 287.8400 ;
      RECT 2497.4200 286.7600 3302.8200 287.8400 ;
      RECT 2446.4800 286.7600 2495.2200 287.8400 ;
      RECT 1007.4200 286.7600 2444.2800 287.8400 ;
      RECT 665.0200 286.7600 1005.2200 287.8400 ;
      RECT 507.4200 286.7600 662.8200 287.8400 ;
      RECT 5.3000 286.7600 505.2200 287.8400 ;
      RECT 0.0000 286.7600 1.7000 287.8400 ;
      RECT 0.0000 285.1200 3370.4200 286.7600 ;
      RECT 3364.7200 284.0400 3370.4200 285.1200 ;
      RECT 3307.6200 284.0400 3361.1200 285.1200 ;
      RECT 2494.8200 284.0400 3305.4200 285.1200 ;
      RECT 2449.0800 284.0400 2492.6200 285.1200 ;
      RECT 1004.8200 284.0400 2446.8800 285.1200 ;
      RECT 667.6200 284.0400 1002.6200 285.1200 ;
      RECT 504.8200 284.0400 665.4200 285.1200 ;
      RECT 9.3000 284.0400 502.6200 285.1200 ;
      RECT 0.0000 284.0400 5.7000 285.1200 ;
      RECT 0.0000 282.4000 3370.4200 284.0400 ;
      RECT 0.0000 281.9300 1.7000 282.4000 ;
      RECT 3368.7200 281.3200 3370.4200 282.4000 ;
      RECT 3305.0200 281.3200 3365.1200 282.4000 ;
      RECT 2497.4200 281.3200 3302.8200 282.4000 ;
      RECT 2446.4800 281.3200 2495.2200 282.4000 ;
      RECT 1007.4200 281.3200 2444.2800 282.4000 ;
      RECT 665.0200 281.3200 1005.2200 282.4000 ;
      RECT 507.4200 281.3200 662.8200 282.4000 ;
      RECT 5.3000 281.3200 505.2200 282.4000 ;
      RECT 1.1000 281.3200 1.7000 281.9300 ;
      RECT 1.1000 281.0300 3370.4200 281.3200 ;
      RECT 0.0000 279.6800 3370.4200 281.0300 ;
      RECT 3364.7200 278.6000 3370.4200 279.6800 ;
      RECT 3307.6200 278.6000 3361.1200 279.6800 ;
      RECT 2494.8200 278.6000 3305.4200 279.6800 ;
      RECT 2449.0800 278.6000 2492.6200 279.6800 ;
      RECT 1004.8200 278.6000 2446.8800 279.6800 ;
      RECT 667.6200 278.6000 1002.6200 279.6800 ;
      RECT 504.8200 278.6000 665.4200 279.6800 ;
      RECT 9.3000 278.6000 502.6200 279.6800 ;
      RECT 0.0000 278.6000 5.7000 279.6800 ;
      RECT 0.0000 276.9600 3370.4200 278.6000 ;
      RECT 3368.7200 275.8800 3370.4200 276.9600 ;
      RECT 3305.0200 275.8800 3365.1200 276.9600 ;
      RECT 2497.4200 275.8800 3302.8200 276.9600 ;
      RECT 2446.4800 275.8800 2495.2200 276.9600 ;
      RECT 1007.4200 275.8800 2444.2800 276.9600 ;
      RECT 665.0200 275.8800 1005.2200 276.9600 ;
      RECT 507.4200 275.8800 662.8200 276.9600 ;
      RECT 5.3000 275.8800 505.2200 276.9600 ;
      RECT 0.0000 275.8800 1.7000 276.9600 ;
      RECT 0.0000 274.2400 3370.4200 275.8800 ;
      RECT 3364.7200 273.1600 3370.4200 274.2400 ;
      RECT 3307.6200 273.1600 3361.1200 274.2400 ;
      RECT 2494.8200 273.1600 3305.4200 274.2400 ;
      RECT 2449.0800 273.1600 2492.6200 274.2400 ;
      RECT 1004.8200 273.1600 2446.8800 274.2400 ;
      RECT 667.6200 273.1600 1002.6200 274.2400 ;
      RECT 504.8200 273.1600 665.4200 274.2400 ;
      RECT 9.3000 273.1600 502.6200 274.2400 ;
      RECT 0.0000 273.1600 5.7000 274.2400 ;
      RECT 0.0000 271.5200 3370.4200 273.1600 ;
      RECT 0.0000 270.9500 1.7000 271.5200 ;
      RECT 3368.7200 270.4400 3370.4200 271.5200 ;
      RECT 3305.0200 270.4400 3365.1200 271.5200 ;
      RECT 2497.4200 270.4400 3302.8200 271.5200 ;
      RECT 2446.4800 270.4400 2495.2200 271.5200 ;
      RECT 1007.4200 270.4400 2444.2800 271.5200 ;
      RECT 665.0200 270.4400 1005.2200 271.5200 ;
      RECT 507.4200 270.4400 662.8200 271.5200 ;
      RECT 5.3000 270.4400 505.2200 271.5200 ;
      RECT 1.1000 270.4400 1.7000 270.9500 ;
      RECT 1.1000 270.0500 3370.4200 270.4400 ;
      RECT 0.0000 268.8000 3370.4200 270.0500 ;
      RECT 3364.7200 267.7200 3370.4200 268.8000 ;
      RECT 3307.6200 267.7200 3361.1200 268.8000 ;
      RECT 2494.8200 267.7200 3305.4200 268.8000 ;
      RECT 2449.0800 267.7200 2492.6200 268.8000 ;
      RECT 1004.8200 267.7200 2446.8800 268.8000 ;
      RECT 667.6200 267.7200 1002.6200 268.8000 ;
      RECT 504.8200 267.7200 665.4200 268.8000 ;
      RECT 9.3000 267.7200 502.6200 268.8000 ;
      RECT 0.0000 267.7200 5.7000 268.8000 ;
      RECT 0.0000 266.0800 3370.4200 267.7200 ;
      RECT 3368.7200 265.0000 3370.4200 266.0800 ;
      RECT 3305.0200 265.0000 3365.1200 266.0800 ;
      RECT 2497.4200 265.0000 3302.8200 266.0800 ;
      RECT 2446.4800 265.0000 2495.2200 266.0800 ;
      RECT 1007.4200 265.0000 2444.2800 266.0800 ;
      RECT 665.0200 265.0000 1005.2200 266.0800 ;
      RECT 507.4200 265.0000 662.8200 266.0800 ;
      RECT 5.3000 265.0000 505.2200 266.0800 ;
      RECT 0.0000 265.0000 1.7000 266.0800 ;
      RECT 0.0000 263.3600 3370.4200 265.0000 ;
      RECT 3364.7200 262.2800 3370.4200 263.3600 ;
      RECT 3307.6200 262.2800 3361.1200 263.3600 ;
      RECT 2494.8200 262.2800 3305.4200 263.3600 ;
      RECT 2449.0800 262.2800 2492.6200 263.3600 ;
      RECT 1004.8200 262.2800 2446.8800 263.3600 ;
      RECT 667.6200 262.2800 1002.6200 263.3600 ;
      RECT 504.8200 262.2800 665.4200 263.3600 ;
      RECT 9.3000 262.2800 502.6200 263.3600 ;
      RECT 0.0000 262.2800 5.7000 263.3600 ;
      RECT 0.0000 260.6400 3370.4200 262.2800 ;
      RECT 0.0000 259.9700 1.7000 260.6400 ;
      RECT 3368.7200 259.5600 3370.4200 260.6400 ;
      RECT 3305.0200 259.5600 3365.1200 260.6400 ;
      RECT 2497.4200 259.5600 3302.8200 260.6400 ;
      RECT 2446.4800 259.5600 2495.2200 260.6400 ;
      RECT 1007.4200 259.5600 2444.2800 260.6400 ;
      RECT 665.0200 259.5600 1005.2200 260.6400 ;
      RECT 507.4200 259.5600 662.8200 260.6400 ;
      RECT 5.3000 259.5600 505.2200 260.6400 ;
      RECT 1.1000 259.5600 1.7000 259.9700 ;
      RECT 1.1000 259.0700 3370.4200 259.5600 ;
      RECT 0.0000 257.9200 3370.4200 259.0700 ;
      RECT 3364.7200 256.8400 3370.4200 257.9200 ;
      RECT 3307.6200 256.8400 3361.1200 257.9200 ;
      RECT 2494.8200 256.8400 3305.4200 257.9200 ;
      RECT 2449.0800 256.8400 2492.6200 257.9200 ;
      RECT 1004.8200 256.8400 2446.8800 257.9200 ;
      RECT 667.6200 256.8400 1002.6200 257.9200 ;
      RECT 504.8200 256.8400 665.4200 257.9200 ;
      RECT 9.3000 256.8400 502.6200 257.9200 ;
      RECT 0.0000 256.8400 5.7000 257.9200 ;
      RECT 0.0000 255.2000 3370.4200 256.8400 ;
      RECT 3368.7200 254.1200 3370.4200 255.2000 ;
      RECT 3305.0200 254.1200 3365.1200 255.2000 ;
      RECT 2497.4200 254.1200 3302.8200 255.2000 ;
      RECT 2446.4800 254.1200 2495.2200 255.2000 ;
      RECT 1007.4200 254.1200 2444.2800 255.2000 ;
      RECT 665.0200 254.1200 1005.2200 255.2000 ;
      RECT 507.4200 254.1200 662.8200 255.2000 ;
      RECT 5.3000 254.1200 505.2200 255.2000 ;
      RECT 0.0000 254.1200 1.7000 255.2000 ;
      RECT 0.0000 252.4800 3370.4200 254.1200 ;
      RECT 3364.7200 251.4000 3370.4200 252.4800 ;
      RECT 3307.6200 251.4000 3361.1200 252.4800 ;
      RECT 2494.8200 251.4000 3305.4200 252.4800 ;
      RECT 2449.0800 251.4000 2492.6200 252.4800 ;
      RECT 1004.8200 251.4000 2446.8800 252.4800 ;
      RECT 667.6200 251.4000 1002.6200 252.4800 ;
      RECT 504.8200 251.4000 665.4200 252.4800 ;
      RECT 9.3000 251.4000 502.6200 252.4800 ;
      RECT 0.0000 251.4000 5.7000 252.4800 ;
      RECT 0.0000 249.7600 3370.4200 251.4000 ;
      RECT 0.0000 248.9900 1.7000 249.7600 ;
      RECT 3368.7200 248.6800 3370.4200 249.7600 ;
      RECT 3305.0200 248.6800 3365.1200 249.7600 ;
      RECT 2497.4200 248.6800 3302.8200 249.7600 ;
      RECT 2446.4800 248.6800 2495.2200 249.7600 ;
      RECT 1007.4200 248.6800 2444.2800 249.7600 ;
      RECT 665.0200 248.6800 1005.2200 249.7600 ;
      RECT 507.4200 248.6800 662.8200 249.7600 ;
      RECT 5.3000 248.6800 505.2200 249.7600 ;
      RECT 1.1000 248.6800 1.7000 248.9900 ;
      RECT 1.1000 248.0900 3370.4200 248.6800 ;
      RECT 0.0000 247.0400 3370.4200 248.0900 ;
      RECT 3364.7200 245.9600 3370.4200 247.0400 ;
      RECT 3307.6200 245.9600 3361.1200 247.0400 ;
      RECT 2494.8200 245.9600 3305.4200 247.0400 ;
      RECT 2449.0800 245.9600 2492.6200 247.0400 ;
      RECT 1004.8200 245.9600 2446.8800 247.0400 ;
      RECT 667.6200 245.9600 1002.6200 247.0400 ;
      RECT 504.8200 245.9600 665.4200 247.0400 ;
      RECT 9.3000 245.9600 502.6200 247.0400 ;
      RECT 0.0000 245.9600 5.7000 247.0400 ;
      RECT 0.0000 244.3200 3370.4200 245.9600 ;
      RECT 3368.7200 243.2400 3370.4200 244.3200 ;
      RECT 3305.0200 243.2400 3365.1200 244.3200 ;
      RECT 2497.4200 243.2400 3302.8200 244.3200 ;
      RECT 2446.4800 243.2400 2495.2200 244.3200 ;
      RECT 1007.4200 243.2400 2444.2800 244.3200 ;
      RECT 665.0200 243.2400 1005.2200 244.3200 ;
      RECT 507.4200 243.2400 662.8200 244.3200 ;
      RECT 5.3000 243.2400 505.2200 244.3200 ;
      RECT 0.0000 243.2400 1.7000 244.3200 ;
      RECT 0.0000 241.6000 3370.4200 243.2400 ;
      RECT 3364.7200 240.5200 3370.4200 241.6000 ;
      RECT 3307.6200 240.5200 3361.1200 241.6000 ;
      RECT 2494.8200 240.5200 3305.4200 241.6000 ;
      RECT 2449.0800 240.5200 2492.6200 241.6000 ;
      RECT 1004.8200 240.5200 2446.8800 241.6000 ;
      RECT 667.6200 240.5200 1002.6200 241.6000 ;
      RECT 504.8200 240.5200 665.4200 241.6000 ;
      RECT 9.3000 240.5200 502.6200 241.6000 ;
      RECT 0.0000 240.5200 5.7000 241.6000 ;
      RECT 0.0000 238.8800 3370.4200 240.5200 ;
      RECT 0.0000 238.6200 1.7000 238.8800 ;
      RECT 3368.7200 237.8000 3370.4200 238.8800 ;
      RECT 3305.0200 237.8000 3365.1200 238.8800 ;
      RECT 2497.4200 237.8000 3302.8200 238.8800 ;
      RECT 2446.4800 237.8000 2495.2200 238.8800 ;
      RECT 1007.4200 237.8000 2444.2800 238.8800 ;
      RECT 665.0200 237.8000 1005.2200 238.8800 ;
      RECT 507.4200 237.8000 662.8200 238.8800 ;
      RECT 5.3000 237.8000 505.2200 238.8800 ;
      RECT 1.1000 237.8000 1.7000 238.6200 ;
      RECT 1.1000 237.7200 3370.4200 237.8000 ;
      RECT 0.0000 236.1600 3370.4200 237.7200 ;
      RECT 3364.7200 235.0800 3370.4200 236.1600 ;
      RECT 3307.6200 235.0800 3361.1200 236.1600 ;
      RECT 2494.8200 235.0800 3305.4200 236.1600 ;
      RECT 2449.0800 235.0800 2492.6200 236.1600 ;
      RECT 1004.8200 235.0800 2446.8800 236.1600 ;
      RECT 667.6200 235.0800 1002.6200 236.1600 ;
      RECT 504.8200 235.0800 665.4200 236.1600 ;
      RECT 9.3000 235.0800 502.6200 236.1600 ;
      RECT 0.0000 235.0800 5.7000 236.1600 ;
      RECT 0.0000 233.4400 3370.4200 235.0800 ;
      RECT 3368.7200 232.3600 3370.4200 233.4400 ;
      RECT 3305.0200 232.3600 3365.1200 233.4400 ;
      RECT 2497.4200 232.3600 3302.8200 233.4400 ;
      RECT 2446.4800 232.3600 2495.2200 233.4400 ;
      RECT 1007.4200 232.3600 2444.2800 233.4400 ;
      RECT 665.0200 232.3600 1005.2200 233.4400 ;
      RECT 507.4200 232.3600 662.8200 233.4400 ;
      RECT 5.3000 232.3600 505.2200 233.4400 ;
      RECT 0.0000 232.3600 1.7000 233.4400 ;
      RECT 0.0000 230.7200 3370.4200 232.3600 ;
      RECT 3364.7200 229.6400 3370.4200 230.7200 ;
      RECT 3307.6200 229.6400 3361.1200 230.7200 ;
      RECT 2494.8200 229.6400 3305.4200 230.7200 ;
      RECT 2449.0800 229.6400 2492.6200 230.7200 ;
      RECT 1004.8200 229.6400 2446.8800 230.7200 ;
      RECT 667.6200 229.6400 1002.6200 230.7200 ;
      RECT 504.8200 229.6400 665.4200 230.7200 ;
      RECT 9.3000 229.6400 502.6200 230.7200 ;
      RECT 0.0000 229.6400 5.7000 230.7200 ;
      RECT 0.0000 228.0000 3370.4200 229.6400 ;
      RECT 0.0000 227.6400 1.7000 228.0000 ;
      RECT 3368.7200 226.9200 3370.4200 228.0000 ;
      RECT 3305.0200 226.9200 3365.1200 228.0000 ;
      RECT 2497.4200 226.9200 3302.8200 228.0000 ;
      RECT 2446.4800 226.9200 2495.2200 228.0000 ;
      RECT 1007.4200 226.9200 2444.2800 228.0000 ;
      RECT 665.0200 226.9200 1005.2200 228.0000 ;
      RECT 507.4200 226.9200 662.8200 228.0000 ;
      RECT 5.3000 226.9200 505.2200 228.0000 ;
      RECT 1.1000 226.9200 1.7000 227.6400 ;
      RECT 1.1000 226.7400 3370.4200 226.9200 ;
      RECT 0.0000 225.2800 3370.4200 226.7400 ;
      RECT 3364.7200 224.2000 3370.4200 225.2800 ;
      RECT 3307.6200 224.2000 3361.1200 225.2800 ;
      RECT 2494.8200 224.2000 3305.4200 225.2800 ;
      RECT 2449.0800 224.2000 2492.6200 225.2800 ;
      RECT 1004.8200 224.2000 2446.8800 225.2800 ;
      RECT 667.6200 224.2000 1002.6200 225.2800 ;
      RECT 504.8200 224.2000 665.4200 225.2800 ;
      RECT 9.3000 224.2000 502.6200 225.2800 ;
      RECT 0.0000 224.2000 5.7000 225.2800 ;
      RECT 0.0000 222.5600 3370.4200 224.2000 ;
      RECT 3368.7200 221.4800 3370.4200 222.5600 ;
      RECT 3305.0200 221.4800 3365.1200 222.5600 ;
      RECT 2497.4200 221.4800 3302.8200 222.5600 ;
      RECT 2446.4800 221.4800 2495.2200 222.5600 ;
      RECT 1007.4200 221.4800 2444.2800 222.5600 ;
      RECT 665.0200 221.4800 1005.2200 222.5600 ;
      RECT 507.4200 221.4800 662.8200 222.5600 ;
      RECT 5.3000 221.4800 505.2200 222.5600 ;
      RECT 0.0000 221.4800 1.7000 222.5600 ;
      RECT 0.0000 219.8400 3370.4200 221.4800 ;
      RECT 3364.7200 218.7600 3370.4200 219.8400 ;
      RECT 3307.6200 218.7600 3361.1200 219.8400 ;
      RECT 2494.8200 218.7600 3305.4200 219.8400 ;
      RECT 2449.0800 218.7600 2492.6200 219.8400 ;
      RECT 1004.8200 218.7600 2446.8800 219.8400 ;
      RECT 667.6200 218.7600 1002.6200 219.8400 ;
      RECT 504.8200 218.7600 665.4200 219.8400 ;
      RECT 9.3000 218.7600 502.6200 219.8400 ;
      RECT 0.0000 218.7600 5.7000 219.8400 ;
      RECT 0.0000 217.1200 3370.4200 218.7600 ;
      RECT 0.0000 216.6600 1.7000 217.1200 ;
      RECT 3368.7200 216.0400 3370.4200 217.1200 ;
      RECT 3305.0200 216.0400 3365.1200 217.1200 ;
      RECT 2497.4200 216.0400 3302.8200 217.1200 ;
      RECT 2446.4800 216.0400 2495.2200 217.1200 ;
      RECT 1007.4200 216.0400 2444.2800 217.1200 ;
      RECT 665.0200 216.0400 1005.2200 217.1200 ;
      RECT 507.4200 216.0400 662.8200 217.1200 ;
      RECT 5.3000 216.0400 505.2200 217.1200 ;
      RECT 1.1000 216.0400 1.7000 216.6600 ;
      RECT 1.1000 215.7600 3370.4200 216.0400 ;
      RECT 0.0000 214.4000 3370.4200 215.7600 ;
      RECT 3364.7200 213.3200 3370.4200 214.4000 ;
      RECT 3307.6200 213.3200 3361.1200 214.4000 ;
      RECT 2494.8200 213.3200 3305.4200 214.4000 ;
      RECT 2449.0800 213.3200 2492.6200 214.4000 ;
      RECT 1004.8200 213.3200 2446.8800 214.4000 ;
      RECT 667.6200 213.3200 1002.6200 214.4000 ;
      RECT 504.8200 213.3200 665.4200 214.4000 ;
      RECT 9.3000 213.3200 502.6200 214.4000 ;
      RECT 0.0000 213.3200 5.7000 214.4000 ;
      RECT 0.0000 211.6800 3370.4200 213.3200 ;
      RECT 3368.7200 210.6000 3370.4200 211.6800 ;
      RECT 3305.0200 210.6000 3365.1200 211.6800 ;
      RECT 2497.4200 210.6000 3302.8200 211.6800 ;
      RECT 2446.4800 210.6000 2495.2200 211.6800 ;
      RECT 1007.4200 210.6000 2444.2800 211.6800 ;
      RECT 665.0200 210.6000 1005.2200 211.6800 ;
      RECT 507.4200 210.6000 662.8200 211.6800 ;
      RECT 5.3000 210.6000 505.2200 211.6800 ;
      RECT 0.0000 210.6000 1.7000 211.6800 ;
      RECT 0.0000 208.9600 3370.4200 210.6000 ;
      RECT 3364.7200 207.8800 3370.4200 208.9600 ;
      RECT 3307.6200 207.8800 3361.1200 208.9600 ;
      RECT 2494.8200 207.8800 3305.4200 208.9600 ;
      RECT 2449.0800 207.8800 2492.6200 208.9600 ;
      RECT 1004.8200 207.8800 2446.8800 208.9600 ;
      RECT 667.6200 207.8800 1002.6200 208.9600 ;
      RECT 504.8200 207.8800 665.4200 208.9600 ;
      RECT 9.3000 207.8800 502.6200 208.9600 ;
      RECT 0.0000 207.8800 5.7000 208.9600 ;
      RECT 0.0000 206.2400 3370.4200 207.8800 ;
      RECT 0.0000 205.6800 1.7000 206.2400 ;
      RECT 3368.7200 205.1600 3370.4200 206.2400 ;
      RECT 3305.0200 205.1600 3365.1200 206.2400 ;
      RECT 2497.4200 205.1600 3302.8200 206.2400 ;
      RECT 2446.4800 205.1600 2495.2200 206.2400 ;
      RECT 1007.4200 205.1600 2444.2800 206.2400 ;
      RECT 665.0200 205.1600 1005.2200 206.2400 ;
      RECT 507.4200 205.1600 662.8200 206.2400 ;
      RECT 5.3000 205.1600 505.2200 206.2400 ;
      RECT 1.1000 205.1600 1.7000 205.6800 ;
      RECT 1.1000 204.7800 3370.4200 205.1600 ;
      RECT 0.0000 203.5200 3370.4200 204.7800 ;
      RECT 3364.7200 202.4400 3370.4200 203.5200 ;
      RECT 3307.6200 202.4400 3361.1200 203.5200 ;
      RECT 2494.8200 202.4400 3305.4200 203.5200 ;
      RECT 2449.0800 202.4400 2492.6200 203.5200 ;
      RECT 1004.8200 202.4400 2446.8800 203.5200 ;
      RECT 667.6200 202.4400 1002.6200 203.5200 ;
      RECT 504.8200 202.4400 665.4200 203.5200 ;
      RECT 9.3000 202.4400 502.6200 203.5200 ;
      RECT 0.0000 202.4400 5.7000 203.5200 ;
      RECT 0.0000 200.8000 3370.4200 202.4400 ;
      RECT 3368.7200 199.7200 3370.4200 200.8000 ;
      RECT 3305.0200 199.7200 3365.1200 200.8000 ;
      RECT 2497.4200 199.7200 3302.8200 200.8000 ;
      RECT 2446.4800 199.7200 2495.2200 200.8000 ;
      RECT 1007.4200 199.7200 2444.2800 200.8000 ;
      RECT 665.0200 199.7200 1005.2200 200.8000 ;
      RECT 507.4200 199.7200 662.8200 200.8000 ;
      RECT 5.3000 199.7200 505.2200 200.8000 ;
      RECT 0.0000 199.7200 1.7000 200.8000 ;
      RECT 0.0000 198.0800 3370.4200 199.7200 ;
      RECT 3364.7200 197.0000 3370.4200 198.0800 ;
      RECT 3307.6200 197.0000 3361.1200 198.0800 ;
      RECT 2494.8200 197.0000 3305.4200 198.0800 ;
      RECT 2449.0800 197.0000 2492.6200 198.0800 ;
      RECT 1004.8200 197.0000 2446.8800 198.0800 ;
      RECT 667.6200 197.0000 1002.6200 198.0800 ;
      RECT 504.8200 197.0000 665.4200 198.0800 ;
      RECT 9.3000 197.0000 502.6200 198.0800 ;
      RECT 0.0000 197.0000 5.7000 198.0800 ;
      RECT 0.0000 195.3600 3370.4200 197.0000 ;
      RECT 0.0000 194.7000 1.7000 195.3600 ;
      RECT 3368.7200 194.2800 3370.4200 195.3600 ;
      RECT 3305.0200 194.2800 3365.1200 195.3600 ;
      RECT 2497.4200 194.2800 3302.8200 195.3600 ;
      RECT 2446.4800 194.2800 2495.2200 195.3600 ;
      RECT 1007.4200 194.2800 2444.2800 195.3600 ;
      RECT 665.0200 194.2800 1005.2200 195.3600 ;
      RECT 507.4200 194.2800 662.8200 195.3600 ;
      RECT 5.3000 194.2800 505.2200 195.3600 ;
      RECT 1.1000 194.2800 1.7000 194.7000 ;
      RECT 1.1000 193.8600 3370.4200 194.2800 ;
      RECT 1.1000 193.8000 1015.2800 193.8600 ;
      RECT 1077.7200 193.6000 3370.4200 193.8600 ;
      RECT 1077.7200 192.7800 1295.6000 193.6000 ;
      RECT 1017.4800 192.7800 1075.5200 193.8600 ;
      RECT 0.0000 192.7800 1015.2800 193.8000 ;
      RECT 2436.3200 192.6400 3370.4200 193.6000 ;
      RECT 0.0000 192.6400 1295.6000 192.7800 ;
      RECT 2436.3200 192.5200 2446.8800 192.6400 ;
      RECT 2178.6800 192.5200 2434.1200 193.6000 ;
      RECT 1958.4600 192.5200 2176.4800 193.6000 ;
      RECT 1738.2400 192.5200 1956.2600 193.6000 ;
      RECT 1518.0200 192.5200 1736.0400 193.6000 ;
      RECT 1297.8000 192.5200 1515.8200 193.6000 ;
      RECT 1004.8200 192.5200 1295.6000 192.6400 ;
      RECT 3364.7200 191.5600 3370.4200 192.6400 ;
      RECT 3307.6200 191.5600 3361.1200 192.6400 ;
      RECT 2494.8200 191.5600 3305.4200 192.6400 ;
      RECT 2449.0800 191.5600 2492.6200 192.6400 ;
      RECT 1004.8200 191.5600 2446.8800 192.5200 ;
      RECT 667.6200 191.5600 1002.6200 192.6400 ;
      RECT 504.8200 191.5600 665.4200 192.6400 ;
      RECT 9.3000 191.5600 502.6200 192.6400 ;
      RECT 0.0000 191.5600 5.7000 192.6400 ;
      RECT 0.0000 190.7900 3370.4200 191.5600 ;
      RECT 0.0000 190.6900 1062.9600 190.7900 ;
      RECT 1285.3800 190.5300 3370.4200 190.7900 ;
      RECT 2446.4800 189.9200 3370.4200 190.5300 ;
      RECT 0.0000 189.9200 1005.2200 190.6900 ;
      RECT 3368.7200 188.8400 3370.4200 189.9200 ;
      RECT 3305.0200 188.8400 3365.1200 189.9200 ;
      RECT 2497.4200 188.8400 3302.8200 189.9200 ;
      RECT 2446.4800 188.8400 2495.2200 189.9200 ;
      RECT 665.0200 188.8400 1005.2200 189.9200 ;
      RECT 507.4200 188.8400 662.8200 189.9200 ;
      RECT 5.3000 188.8400 505.2200 189.9200 ;
      RECT 0.0000 188.8400 1.7000 189.9200 ;
      RECT 1071.3600 188.5900 1279.3800 190.7900 ;
      RECT 1065.1600 188.4900 1283.0400 188.5900 ;
      RECT 1011.2200 188.4900 1059.1600 190.6900 ;
      RECT 0.0000 188.4900 1005.2200 188.8400 ;
      RECT 2446.4800 188.3300 3370.4200 188.8400 ;
      RECT 2392.5400 188.3300 2440.4800 190.5300 ;
      RECT 2172.3200 188.3300 2384.1400 190.5300 ;
      RECT 1952.1000 188.3300 2160.1200 190.5300 ;
      RECT 1731.8800 188.3300 1943.7000 190.5300 ;
      RECT 1511.6600 188.3300 1723.4800 190.5300 ;
      RECT 1291.4400 188.3300 1503.2600 190.5300 ;
      RECT 0.0000 188.3300 1283.0400 188.4900 ;
      RECT 0.0000 188.2900 3370.4200 188.3300 ;
      RECT 1067.7600 188.1900 3370.4200 188.2900 ;
      RECT 1287.9800 187.9300 3370.4200 188.1900 ;
      RECT 2392.5400 187.2000 3370.4200 187.9300 ;
      RECT 0.0000 187.2000 1002.6200 188.2900 ;
      RECT 3364.7200 186.1200 3370.4200 187.2000 ;
      RECT 3307.6200 186.1200 3361.1200 187.2000 ;
      RECT 2494.8200 186.1200 3305.4200 187.2000 ;
      RECT 2449.0800 186.1200 2492.6200 187.2000 ;
      RECT 2392.5400 186.1200 2446.8800 187.2000 ;
      RECT 667.6200 186.1200 1002.6200 187.2000 ;
      RECT 504.8200 186.1200 665.4200 187.2000 ;
      RECT 9.3000 186.1200 502.6200 187.2000 ;
      RECT 0.0000 186.1200 5.7000 187.2000 ;
      RECT 1011.2200 186.0900 1059.1600 188.2900 ;
      RECT 0.0000 186.0900 1002.6200 186.1200 ;
      RECT 1071.3600 185.9900 1279.3800 188.1900 ;
      RECT 0.0000 185.9900 1065.5600 186.0900 ;
      RECT 2392.5400 185.7300 3370.4200 186.1200 ;
      RECT 2172.3200 185.7300 2386.7400 187.9300 ;
      RECT 1952.1000 185.7300 2166.5200 187.9300 ;
      RECT 1731.8800 185.7300 1946.3000 187.9300 ;
      RECT 1511.6600 185.7300 1726.0800 187.9300 ;
      RECT 1291.4400 185.7300 1505.8600 187.9300 ;
      RECT 0.0000 185.7300 1285.6400 185.9900 ;
      RECT 0.0000 184.4800 3370.4200 185.7300 ;
      RECT 0.0000 184.3300 1.7000 184.4800 ;
      RECT 1.1000 183.4300 1.7000 184.3300 ;
      RECT 3368.7200 183.4000 3370.4200 184.4800 ;
      RECT 3305.0200 183.4000 3365.1200 184.4800 ;
      RECT 2497.4200 183.4000 3302.8200 184.4800 ;
      RECT 2446.4800 183.4000 2495.2200 184.4800 ;
      RECT 1007.4200 183.4000 2444.2800 184.4800 ;
      RECT 665.0200 183.4000 1005.2200 184.4800 ;
      RECT 507.4200 183.4000 662.8200 184.4800 ;
      RECT 5.3000 183.4000 505.2200 184.4800 ;
      RECT 0.0000 183.4000 1.7000 183.4300 ;
      RECT 0.0000 181.7600 3370.4200 183.4000 ;
      RECT 1004.8200 180.7600 2446.8800 181.7600 ;
      RECT 667.6200 180.7600 1002.6200 181.7600 ;
      RECT 504.8200 180.7600 665.4200 181.7600 ;
      RECT 9.3000 180.7600 502.6200 181.7600 ;
      RECT 0.0000 180.7600 5.7000 181.7600 ;
      RECT 3364.7200 180.6800 3370.4200 181.7600 ;
      RECT 3307.6200 180.6800 3361.1200 181.7600 ;
      RECT 2494.8200 180.6800 3305.4200 181.7600 ;
      RECT 2449.0800 180.6800 2492.6200 181.7600 ;
      RECT 1285.3800 180.6800 2446.8800 180.7600 ;
      RECT 1285.3800 180.5000 3370.4200 180.6800 ;
      RECT 2446.4800 179.0400 3370.4200 180.5000 ;
      RECT 5.3000 178.3000 1283.0400 178.5600 ;
      RECT 5.3000 178.2600 2444.2800 178.3000 ;
      RECT 1065.0600 178.1600 2444.2800 178.2600 ;
      RECT 5.3000 178.1600 1062.6600 178.2600 ;
      RECT 5.3000 178.1300 5.7000 178.1600 ;
      RECT 0.0000 178.1300 1.7000 180.7600 ;
      RECT 3368.7200 177.9600 3370.4200 179.0400 ;
      RECT 3305.0200 177.9600 3365.1200 179.0400 ;
      RECT 2497.4200 177.9600 3302.8200 179.0400 ;
      RECT 2446.4800 177.9600 2495.2200 179.0400 ;
      RECT 1287.9800 177.9600 2444.2800 178.1600 ;
      RECT 1287.9800 177.9000 3370.4200 177.9600 ;
      RECT 2449.0800 176.3200 3370.4200 177.9000 ;
      RECT 1065.0600 175.7000 1285.6400 175.9600 ;
      RECT 3364.7200 175.2400 3370.4200 176.3200 ;
      RECT 3307.6200 175.2400 3361.1200 176.3200 ;
      RECT 2494.8200 175.2400 3305.4200 176.3200 ;
      RECT 2449.0800 175.2400 2492.6200 176.3200 ;
      RECT 1065.0600 175.2400 2446.8800 175.7000 ;
      RECT 9.3000 175.0700 1062.6600 175.9600 ;
      RECT 0.0000 175.0700 5.7000 178.1300 ;
      RECT 1065.0600 174.2600 3370.4200 175.2400 ;
      RECT 0.0000 174.2600 1062.6600 175.0700 ;
      RECT 0.0000 173.6000 3370.4200 174.2600 ;
      RECT 0.0000 173.3500 1.7000 173.6000 ;
      RECT 3368.7200 172.5200 3370.4200 173.6000 ;
      RECT 3305.0200 172.5200 3365.1200 173.6000 ;
      RECT 2497.4200 172.5200 3302.8200 173.6000 ;
      RECT 2446.4800 172.5200 2495.2200 173.6000 ;
      RECT 2386.3400 172.5200 2444.2800 173.6000 ;
      RECT 1065.1600 172.5200 2384.1400 173.6000 ;
      RECT 5.3000 172.5200 1062.9600 173.6000 ;
      RECT 1.1000 172.5200 1.7000 173.3500 ;
      RECT 1.1000 172.4500 3370.4200 172.5200 ;
      RECT 0.0000 171.0000 3370.4200 172.4500 ;
      RECT 1287.9800 170.8800 3370.4200 171.0000 ;
      RECT 0.0000 170.8800 1065.5600 171.0000 ;
      RECT 1287.9800 170.7400 2386.7400 170.8800 ;
      RECT 3364.7200 169.8000 3370.4200 170.8800 ;
      RECT 3307.6200 169.8000 3361.1200 170.8800 ;
      RECT 2494.8200 169.8000 3305.4200 170.8800 ;
      RECT 2449.0800 169.8000 2492.6200 170.8800 ;
      RECT 2388.9400 169.8000 2446.8800 170.8800 ;
      RECT 9.3000 169.8000 1065.5600 170.8800 ;
      RECT 0.0000 169.8000 5.7000 170.8800 ;
      RECT 1071.3600 168.8000 1279.3800 171.0000 ;
      RECT 0.0000 168.8000 1065.5600 169.8000 ;
      RECT 0.0000 168.6000 1285.6400 168.8000 ;
      RECT 2388.9400 168.5400 3370.4200 169.8000 ;
      RECT 2172.3200 168.5400 2380.3400 170.7400 ;
      RECT 1952.1000 168.5400 2160.1200 170.7400 ;
      RECT 1731.8800 168.5400 1939.9000 170.7400 ;
      RECT 1511.6600 168.5400 1719.6800 170.7400 ;
      RECT 1291.4400 168.5400 1499.4600 170.7400 ;
      RECT 1285.3800 168.5400 1285.6400 168.6000 ;
      RECT 1285.3800 168.3400 3370.4200 168.5400 ;
      RECT 2386.3400 168.1600 3370.4200 168.3400 ;
      RECT 0.0000 168.1600 1062.9600 168.6000 ;
      RECT 3368.7200 167.0800 3370.4200 168.1600 ;
      RECT 3305.0200 167.0800 3365.1200 168.1600 ;
      RECT 2497.4200 167.0800 3302.8200 168.1600 ;
      RECT 2446.4800 167.0800 2495.2200 168.1600 ;
      RECT 2386.3400 167.0800 2444.2800 168.1600 ;
      RECT 5.3000 167.0800 1062.9600 168.1600 ;
      RECT 0.0000 167.0800 1.7000 168.1600 ;
      RECT 1071.3600 166.4000 1279.3800 168.6000 ;
      RECT 0.0000 166.4000 1062.9600 167.0800 ;
      RECT 2386.3400 166.1400 3370.4200 167.0800 ;
      RECT 2172.3200 166.1400 2380.3400 168.3400 ;
      RECT 1952.1000 166.1400 2160.1200 168.3400 ;
      RECT 1731.8800 166.1400 1939.9000 168.3400 ;
      RECT 1511.6600 166.1400 1719.6800 168.3400 ;
      RECT 1291.4400 166.1400 1499.4600 168.3400 ;
      RECT 0.0000 166.1400 1283.0400 166.4000 ;
      RECT 0.0000 165.4400 3370.4200 166.1400 ;
      RECT 1067.7600 164.4800 2386.7400 165.4400 ;
      RECT 3364.7200 164.3600 3370.4200 165.4400 ;
      RECT 3307.6200 164.3600 3361.1200 165.4400 ;
      RECT 2494.8200 164.3600 3305.4200 165.4400 ;
      RECT 2449.0800 164.3600 2492.6200 165.4400 ;
      RECT 2388.9400 164.3600 2446.8800 165.4400 ;
      RECT 1075.2200 164.3600 2386.7400 164.4800 ;
      RECT 1067.7600 164.3600 1073.0200 164.4800 ;
      RECT 9.3000 164.3600 1065.5600 165.4400 ;
      RECT 0.0000 164.3600 5.7000 165.4400 ;
      RECT 1075.2200 164.2200 3370.4200 164.3600 ;
      RECT 1075.2200 163.4000 1293.1000 164.2200 ;
      RECT 0.0000 163.4000 1073.0200 164.3600 ;
      RECT 2176.1800 163.1400 3370.4200 164.2200 ;
      RECT 1955.9600 163.1400 2173.9800 164.2200 ;
      RECT 1735.7400 163.1400 1953.7600 164.2200 ;
      RECT 1515.5200 163.1400 1733.5400 164.2200 ;
      RECT 1295.3000 163.1400 1513.3200 164.2200 ;
      RECT 0.0000 163.1400 1293.1000 163.4000 ;
      RECT 0.0000 162.7200 3370.4200 163.1400 ;
      RECT 0.0000 162.3700 1.7000 162.7200 ;
      RECT 3368.7200 161.6400 3370.4200 162.7200 ;
      RECT 3305.0200 161.6400 3365.1200 162.7200 ;
      RECT 2497.4200 161.6400 3302.8200 162.7200 ;
      RECT 2446.4800 161.6400 2495.2200 162.7200 ;
      RECT 2386.3400 161.6400 2444.2800 162.7200 ;
      RECT 1065.1600 161.6400 2384.1400 162.7200 ;
      RECT 5.3000 161.6400 1062.9600 162.7200 ;
      RECT 1.1000 161.6400 1.7000 162.3700 ;
      RECT 1.1000 161.4700 3370.4200 161.6400 ;
      RECT 0.0000 160.0000 3370.4200 161.4700 ;
      RECT 3364.7200 158.9200 3370.4200 160.0000 ;
      RECT 3307.6200 158.9200 3361.1200 160.0000 ;
      RECT 2494.8200 158.9200 3305.4200 160.0000 ;
      RECT 2449.0800 158.9200 2492.6200 160.0000 ;
      RECT 2388.9400 158.9200 2446.8800 160.0000 ;
      RECT 1067.7600 158.9200 2386.7400 160.0000 ;
      RECT 9.3000 158.9200 1065.5600 160.0000 ;
      RECT 0.0000 158.9200 5.7000 160.0000 ;
      RECT 0.0000 157.2800 3370.4200 158.9200 ;
      RECT 3368.7200 156.2000 3370.4200 157.2800 ;
      RECT 3305.0200 156.2000 3365.1200 157.2800 ;
      RECT 2497.4200 156.2000 3302.8200 157.2800 ;
      RECT 2446.4800 156.2000 2495.2200 157.2800 ;
      RECT 2386.3400 156.2000 2444.2800 157.2800 ;
      RECT 1065.1600 156.2000 2384.1400 157.2800 ;
      RECT 5.3000 156.2000 1062.9600 157.2800 ;
      RECT 0.0000 156.2000 1.7000 157.2800 ;
      RECT 0.0000 154.5600 3370.4200 156.2000 ;
      RECT 3364.7200 153.4800 3370.4200 154.5600 ;
      RECT 3307.6200 153.4800 3361.1200 154.5600 ;
      RECT 2494.8200 153.4800 3305.4200 154.5600 ;
      RECT 2449.0800 153.4800 2492.6200 154.5600 ;
      RECT 2388.9400 153.4800 2446.8800 154.5600 ;
      RECT 1067.7600 153.4800 2386.7400 154.5600 ;
      RECT 9.3000 153.4800 1065.5600 154.5600 ;
      RECT 0.0000 153.4800 5.7000 154.5600 ;
      RECT 0.0000 151.8400 3370.4200 153.4800 ;
      RECT 0.0000 151.3900 1.7000 151.8400 ;
      RECT 1065.1600 150.8800 2384.1400 151.8400 ;
      RECT 3368.7200 150.7600 3370.4200 151.8400 ;
      RECT 3305.0200 150.7600 3365.1200 151.8400 ;
      RECT 2497.4200 150.7600 3302.8200 151.8400 ;
      RECT 2446.4800 150.7600 2495.2200 151.8400 ;
      RECT 2386.3400 150.7600 2444.2800 151.8400 ;
      RECT 1275.3200 150.7600 2384.1400 150.8800 ;
      RECT 1065.1600 150.7600 1273.1200 150.8800 ;
      RECT 5.3000 150.7600 1062.9600 151.8400 ;
      RECT 1.1000 150.7600 1.7000 151.3900 ;
      RECT 1275.3200 150.6200 3370.4200 150.7600 ;
      RECT 1.1000 150.4900 1273.1200 150.7600 ;
      RECT 0.0000 149.9700 1273.1200 150.4900 ;
      RECT 1275.3200 149.8000 1493.2000 150.6200 ;
      RECT 1067.7600 149.8000 1273.1200 149.9700 ;
      RECT 2376.2800 149.5400 3370.4200 150.6200 ;
      RECT 2156.0600 149.5400 2374.0800 150.6200 ;
      RECT 1935.8400 149.5400 2153.8600 150.6200 ;
      RECT 1715.6200 149.5400 1933.6400 150.6200 ;
      RECT 1495.4000 149.5400 1713.4200 150.6200 ;
      RECT 1067.7600 149.5400 1493.2000 149.8000 ;
      RECT 1067.7600 149.1200 3370.4200 149.5400 ;
      RECT 0.0000 149.1200 1065.5600 149.9700 ;
      RECT 1067.7600 149.0700 2386.7400 149.1200 ;
      RECT 9.3000 149.0700 1065.5600 149.1200 ;
      RECT 1285.3800 148.8100 2386.7400 149.0700 ;
      RECT 3364.7200 148.0400 3370.4200 149.1200 ;
      RECT 3307.6200 148.0400 3361.1200 149.1200 ;
      RECT 2494.8200 148.0400 3305.4200 149.1200 ;
      RECT 2449.0800 148.0400 2492.6200 149.1200 ;
      RECT 2388.9400 148.0400 2446.8800 149.1200 ;
      RECT 2386.3400 148.0400 2386.7400 148.8100 ;
      RECT 9.3000 148.0400 1062.9600 149.0700 ;
      RECT 0.0000 148.0400 5.7000 149.1200 ;
      RECT 1071.3600 146.8700 1279.3800 149.0700 ;
      RECT 0.0000 146.8700 1062.9600 148.0400 ;
      RECT 0.0000 146.6700 1283.0400 146.8700 ;
      RECT 2386.3400 146.6100 3370.4200 148.0400 ;
      RECT 2172.3200 146.6100 2380.3400 148.8100 ;
      RECT 1952.1000 146.6100 2160.1200 148.8100 ;
      RECT 1731.8800 146.6100 1939.9000 148.8100 ;
      RECT 1511.6600 146.6100 1719.6800 148.8100 ;
      RECT 1291.4400 146.6100 1499.4600 148.8100 ;
      RECT 1071.3600 146.6100 1283.0400 146.6700 ;
      RECT 1071.3600 146.4100 3370.4200 146.6100 ;
      RECT 2172.3200 146.4000 3370.4200 146.4100 ;
      RECT 0.0000 146.4000 1065.5600 146.6700 ;
      RECT 3368.7200 145.3200 3370.4200 146.4000 ;
      RECT 3305.0200 145.3200 3365.1200 146.4000 ;
      RECT 2497.4200 145.3200 3302.8200 146.4000 ;
      RECT 2446.4800 145.3200 2495.2200 146.4000 ;
      RECT 2386.3400 145.3200 2444.2800 146.4000 ;
      RECT 2172.3200 145.3200 2384.1400 146.4000 ;
      RECT 1065.1600 145.3200 1065.5600 146.4000 ;
      RECT 5.3000 145.3200 1062.9600 146.4000 ;
      RECT 0.0000 145.3200 1.7000 146.4000 ;
      RECT 1071.3600 144.4700 1285.6400 146.4100 ;
      RECT 0.0000 144.4700 1065.5600 145.3200 ;
      RECT 2172.3200 144.2100 3370.4200 145.3200 ;
      RECT 1952.1000 144.2100 2160.1200 146.4100 ;
      RECT 1731.8800 144.2100 1946.3000 146.4100 ;
      RECT 1511.6600 144.2100 1726.0800 146.4100 ;
      RECT 1291.4400 144.2100 1499.4600 146.4100 ;
      RECT 0.0000 144.2100 1285.6400 144.4700 ;
      RECT 0.0000 143.6800 3370.4200 144.2100 ;
      RECT 3364.7200 142.6000 3370.4200 143.6800 ;
      RECT 3307.6200 142.6000 3361.1200 143.6800 ;
      RECT 2494.8200 142.6000 3305.4200 143.6800 ;
      RECT 2449.0800 142.6000 2492.6200 143.6800 ;
      RECT 2388.9400 142.6000 2446.8800 143.6800 ;
      RECT 1067.7600 142.6000 2386.7400 143.6800 ;
      RECT 9.3000 142.6000 1065.5600 143.6800 ;
      RECT 0.0000 142.6000 5.7000 143.6800 ;
      RECT 0.0000 141.1100 3370.4200 142.6000 ;
      RECT 2386.3400 140.9600 3370.4200 141.1100 ;
      RECT 0.0000 140.9600 2384.1400 141.1100 ;
      RECT 1065.1600 140.5000 2384.1400 140.9600 ;
      RECT 0.0000 140.4100 1.7000 140.9600 ;
      RECT 1285.3800 140.2400 2384.1400 140.5000 ;
      RECT 3368.7200 139.8800 3370.4200 140.9600 ;
      RECT 3305.0200 139.8800 3365.1200 140.9600 ;
      RECT 2497.4200 139.8800 3302.8200 140.9600 ;
      RECT 2446.4800 139.8800 2495.2200 140.9600 ;
      RECT 2386.3400 139.8800 2444.2800 140.9600 ;
      RECT 5.3000 139.8800 1062.9600 140.9600 ;
      RECT 1.1000 139.8800 1.7000 140.4100 ;
      RECT 1.1000 139.5100 1062.9600 139.8800 ;
      RECT 0.0000 138.3000 1062.9600 139.5100 ;
      RECT 2386.3400 138.2400 3370.4200 139.8800 ;
      RECT 0.0000 138.2400 1283.0400 138.3000 ;
      RECT 2386.3400 138.0400 2389.2000 138.2400 ;
      RECT 1067.7600 138.0400 1283.0400 138.2400 ;
      RECT 1067.7600 137.9000 2389.2000 138.0400 ;
      RECT 1287.9800 137.6400 2389.2000 137.9000 ;
      RECT 3364.7200 137.1600 3370.4200 138.2400 ;
      RECT 3307.6200 137.1600 3361.1200 138.2400 ;
      RECT 2494.8200 137.1600 3305.4200 138.2400 ;
      RECT 2449.0800 137.1600 2492.6200 138.2400 ;
      RECT 2390.3000 137.1600 2446.8800 138.2400 ;
      RECT 2388.9400 137.1600 2389.2000 137.6400 ;
      RECT 9.3000 137.1600 1065.5600 138.2400 ;
      RECT 0.0000 137.1600 5.7000 138.2400 ;
      RECT 0.0000 135.7000 1065.5600 137.1600 ;
      RECT 2388.9400 135.5200 3370.4200 137.1600 ;
      RECT 0.0000 135.5200 1285.6400 135.7000 ;
      RECT 2388.9400 135.4400 2444.2800 135.5200 ;
      RECT 1065.1600 135.4400 1285.6400 135.5200 ;
      RECT 3368.7200 134.4400 3370.4200 135.5200 ;
      RECT 3305.0200 134.4400 3365.1200 135.5200 ;
      RECT 2497.4200 134.4400 3302.8200 135.5200 ;
      RECT 2446.4800 134.4400 2495.2200 135.5200 ;
      RECT 2386.3400 134.4400 2444.2800 135.4400 ;
      RECT 1065.1600 134.4400 2384.1400 135.4400 ;
      RECT 5.3000 134.4400 1062.9600 135.5200 ;
      RECT 0.0000 134.4400 1.7000 135.5200 ;
      RECT 0.0000 132.8000 3370.4200 134.4400 ;
      RECT 3364.7200 131.7200 3370.4200 132.8000 ;
      RECT 3307.6200 131.7200 3361.1200 132.8000 ;
      RECT 2494.8200 131.7200 3305.4200 132.8000 ;
      RECT 2449.0800 131.7200 2492.6200 132.8000 ;
      RECT 2388.9400 131.7200 2446.8800 132.8000 ;
      RECT 2168.7200 131.7200 2386.7400 132.8000 ;
      RECT 1948.5000 131.7200 2166.5200 132.8000 ;
      RECT 1728.2800 131.7200 1946.3000 132.8000 ;
      RECT 1508.0600 131.7200 1726.0800 132.8000 ;
      RECT 1287.9800 131.7200 1505.8600 132.8000 ;
      RECT 1067.7600 131.7200 1285.6400 132.8000 ;
      RECT 9.3000 131.7200 1065.5600 132.8000 ;
      RECT 0.0000 131.7200 5.7000 132.8000 ;
      RECT 0.0000 130.0800 3370.4200 131.7200 ;
      RECT 0.0000 130.0400 1.7000 130.0800 ;
      RECT 1.1000 129.1400 1.7000 130.0400 ;
      RECT 3368.7200 129.0000 3370.4200 130.0800 ;
      RECT 3305.0200 129.0000 3365.1200 130.0800 ;
      RECT 2497.4200 129.0000 3302.8200 130.0800 ;
      RECT 2446.4800 129.0000 2495.2200 130.0800 ;
      RECT 2386.3400 129.0000 2444.2800 130.0800 ;
      RECT 2166.1200 129.0000 2384.1400 130.0800 ;
      RECT 1945.9000 129.0000 2163.9200 130.0800 ;
      RECT 1725.6800 129.0000 1943.7000 130.0800 ;
      RECT 1505.4600 129.0000 1723.4800 130.0800 ;
      RECT 1285.3800 129.0000 1503.2600 130.0800 ;
      RECT 1065.1600 129.0000 1283.0400 130.0800 ;
      RECT 5.3000 129.0000 1062.9600 130.0800 ;
      RECT 0.0000 129.0000 1.7000 129.1400 ;
      RECT 0.0000 127.3600 3370.4200 129.0000 ;
      RECT 3364.7200 126.2800 3370.4200 127.3600 ;
      RECT 3307.6200 126.2800 3361.1200 127.3600 ;
      RECT 2494.8200 126.2800 3305.4200 127.3600 ;
      RECT 2449.0800 126.2800 2492.6200 127.3600 ;
      RECT 2388.9400 126.2800 2446.8800 127.3600 ;
      RECT 2168.7200 126.2800 2386.7400 127.3600 ;
      RECT 1948.5000 126.2800 2166.5200 127.3600 ;
      RECT 1728.2800 126.2800 1946.3000 127.3600 ;
      RECT 1508.0600 126.2800 1726.0800 127.3600 ;
      RECT 1287.9800 126.2800 1505.8600 127.3600 ;
      RECT 1067.7600 126.2800 1285.6400 127.3600 ;
      RECT 9.3000 126.2800 1065.5600 127.3600 ;
      RECT 0.0000 126.2800 5.7000 127.3600 ;
      RECT 0.0000 124.6400 3370.4200 126.2800 ;
      RECT 3368.7200 123.5600 3370.4200 124.6400 ;
      RECT 3305.0200 123.5600 3365.1200 124.6400 ;
      RECT 2497.4200 123.5600 3302.8200 124.6400 ;
      RECT 2446.4800 123.5600 2495.2200 124.6400 ;
      RECT 2386.3400 123.5600 2444.2800 124.6400 ;
      RECT 2166.1200 123.5600 2384.1400 124.6400 ;
      RECT 1945.9000 123.5600 2163.9200 124.6400 ;
      RECT 1725.6800 123.5600 1943.7000 124.6400 ;
      RECT 1505.4600 123.5600 1723.4800 124.6400 ;
      RECT 1285.3800 123.5600 1503.2600 124.6400 ;
      RECT 1065.1600 123.5600 1283.0400 124.6400 ;
      RECT 5.3000 123.5600 1062.9600 124.6400 ;
      RECT 0.0000 123.5600 1.7000 124.6400 ;
      RECT 0.0000 121.9200 3370.4200 123.5600 ;
      RECT 3364.7200 120.8400 3370.4200 121.9200 ;
      RECT 3307.6200 120.8400 3361.1200 121.9200 ;
      RECT 2494.8200 120.8400 3305.4200 121.9200 ;
      RECT 2449.0800 120.8400 2492.6200 121.9200 ;
      RECT 2388.9400 120.8400 2446.8800 121.9200 ;
      RECT 2168.7200 120.8400 2386.7400 121.9200 ;
      RECT 1948.5000 120.8400 2166.5200 121.9200 ;
      RECT 1728.2800 120.8400 1946.3000 121.9200 ;
      RECT 1508.0600 120.8400 1726.0800 121.9200 ;
      RECT 1287.9800 120.8400 1505.8600 121.9200 ;
      RECT 1067.7600 120.8400 1285.6400 121.9200 ;
      RECT 9.3000 120.8400 1065.5600 121.9200 ;
      RECT 0.0000 120.8400 5.7000 121.9200 ;
      RECT 0.0000 119.2000 3370.4200 120.8400 ;
      RECT 0.0000 119.0600 1.7000 119.2000 ;
      RECT 1.1000 118.1600 1.7000 119.0600 ;
      RECT 3368.7200 118.1200 3370.4200 119.2000 ;
      RECT 3305.0200 118.1200 3365.1200 119.2000 ;
      RECT 2497.4200 118.1200 3302.8200 119.2000 ;
      RECT 2446.4800 118.1200 2495.2200 119.2000 ;
      RECT 2386.3400 118.1200 2444.2800 119.2000 ;
      RECT 2166.1200 118.1200 2384.1400 119.2000 ;
      RECT 1945.9000 118.1200 2163.9200 119.2000 ;
      RECT 1725.6800 118.1200 1943.7000 119.2000 ;
      RECT 1505.4600 118.1200 1723.4800 119.2000 ;
      RECT 1285.3800 118.1200 1503.2600 119.2000 ;
      RECT 1065.1600 118.1200 1283.0400 119.2000 ;
      RECT 5.3000 118.1200 1062.9600 119.2000 ;
      RECT 0.0000 118.1200 1.7000 118.1600 ;
      RECT 0.0000 116.4800 3370.4200 118.1200 ;
      RECT 3364.7200 115.4000 3370.4200 116.4800 ;
      RECT 3307.6200 115.4000 3361.1200 116.4800 ;
      RECT 2494.8200 115.4000 3305.4200 116.4800 ;
      RECT 2449.0800 115.4000 2492.6200 116.4800 ;
      RECT 2388.9400 115.4000 2446.8800 116.4800 ;
      RECT 2168.7200 115.4000 2386.7400 116.4800 ;
      RECT 1948.5000 115.4000 2166.5200 116.4800 ;
      RECT 1728.2800 115.4000 1946.3000 116.4800 ;
      RECT 1508.0600 115.4000 1726.0800 116.4800 ;
      RECT 1287.9800 115.4000 1505.8600 116.4800 ;
      RECT 1067.7600 115.4000 1285.6400 116.4800 ;
      RECT 9.3000 115.4000 1065.5600 116.4800 ;
      RECT 0.0000 115.4000 5.7000 116.4800 ;
      RECT 0.0000 113.7600 3370.4200 115.4000 ;
      RECT 3368.7200 112.6800 3370.4200 113.7600 ;
      RECT 3305.0200 112.6800 3365.1200 113.7600 ;
      RECT 2497.4200 112.6800 3302.8200 113.7600 ;
      RECT 2446.4800 112.6800 2495.2200 113.7600 ;
      RECT 2386.3400 112.6800 2444.2800 113.7600 ;
      RECT 2166.1200 112.6800 2384.1400 113.7600 ;
      RECT 1945.9000 112.6800 2163.9200 113.7600 ;
      RECT 1725.6800 112.6800 1943.7000 113.7600 ;
      RECT 1505.4600 112.6800 1723.4800 113.7600 ;
      RECT 1285.3800 112.6800 1503.2600 113.7600 ;
      RECT 1065.1600 112.6800 1283.0400 113.7600 ;
      RECT 5.3000 112.6800 1062.9600 113.7600 ;
      RECT 0.0000 112.6800 1.7000 113.7600 ;
      RECT 0.0000 111.0400 3370.4200 112.6800 ;
      RECT 3364.7200 109.9600 3370.4200 111.0400 ;
      RECT 3307.6200 109.9600 3361.1200 111.0400 ;
      RECT 2494.8200 109.9600 3305.4200 111.0400 ;
      RECT 2449.0800 109.9600 2492.6200 111.0400 ;
      RECT 2388.9400 109.9600 2446.8800 111.0400 ;
      RECT 2168.7200 109.9600 2386.7400 111.0400 ;
      RECT 1948.5000 109.9600 2166.5200 111.0400 ;
      RECT 1728.2800 109.9600 1946.3000 111.0400 ;
      RECT 1508.0600 109.9600 1726.0800 111.0400 ;
      RECT 1287.9800 109.9600 1505.8600 111.0400 ;
      RECT 1067.7600 109.9600 1285.6400 111.0400 ;
      RECT 9.3000 109.9600 1065.5600 111.0400 ;
      RECT 0.0000 109.9600 5.7000 111.0400 ;
      RECT 0.0000 108.3200 3370.4200 109.9600 ;
      RECT 0.0000 108.0800 1.7000 108.3200 ;
      RECT 3368.7200 107.2400 3370.4200 108.3200 ;
      RECT 3305.0200 107.2400 3365.1200 108.3200 ;
      RECT 2497.4200 107.2400 3302.8200 108.3200 ;
      RECT 2446.4800 107.2400 2495.2200 108.3200 ;
      RECT 2386.3400 107.2400 2444.2800 108.3200 ;
      RECT 2166.1200 107.2400 2384.1400 108.3200 ;
      RECT 1945.9000 107.2400 2163.9200 108.3200 ;
      RECT 1725.6800 107.2400 1943.7000 108.3200 ;
      RECT 1505.4600 107.2400 1723.4800 108.3200 ;
      RECT 1285.3800 107.2400 1503.2600 108.3200 ;
      RECT 1065.1600 107.2400 1283.0400 108.3200 ;
      RECT 5.3000 107.2400 1062.9600 108.3200 ;
      RECT 1.1000 107.2400 1.7000 108.0800 ;
      RECT 1.1000 107.1800 3370.4200 107.2400 ;
      RECT 0.0000 105.6000 3370.4200 107.1800 ;
      RECT 3364.7200 104.5200 3370.4200 105.6000 ;
      RECT 3307.6200 104.5200 3361.1200 105.6000 ;
      RECT 2494.8200 104.5200 3305.4200 105.6000 ;
      RECT 2449.0800 104.5200 2492.6200 105.6000 ;
      RECT 2388.9400 104.5200 2446.8800 105.6000 ;
      RECT 2168.7200 104.5200 2386.7400 105.6000 ;
      RECT 1948.5000 104.5200 2166.5200 105.6000 ;
      RECT 1728.2800 104.5200 1946.3000 105.6000 ;
      RECT 1508.0600 104.5200 1726.0800 105.6000 ;
      RECT 1287.9800 104.5200 1505.8600 105.6000 ;
      RECT 1067.7600 104.5200 1285.6400 105.6000 ;
      RECT 9.3000 104.5200 1065.5600 105.6000 ;
      RECT 0.0000 104.5200 5.7000 105.6000 ;
      RECT 0.0000 102.8800 3370.4200 104.5200 ;
      RECT 3368.7200 101.8000 3370.4200 102.8800 ;
      RECT 3305.0200 101.8000 3365.1200 102.8800 ;
      RECT 2497.4200 101.8000 3302.8200 102.8800 ;
      RECT 2446.4800 101.8000 2495.2200 102.8800 ;
      RECT 2386.3400 101.8000 2444.2800 102.8800 ;
      RECT 2166.1200 101.8000 2384.1400 102.8800 ;
      RECT 1945.9000 101.8000 2163.9200 102.8800 ;
      RECT 1725.6800 101.8000 1943.7000 102.8800 ;
      RECT 1505.4600 101.8000 1723.4800 102.8800 ;
      RECT 1285.3800 101.8000 1503.2600 102.8800 ;
      RECT 1065.1600 101.8000 1283.0400 102.8800 ;
      RECT 5.3000 101.8000 1062.9600 102.8800 ;
      RECT 0.0000 101.8000 1.7000 102.8800 ;
      RECT 0.0000 100.1600 3370.4200 101.8000 ;
      RECT 3364.7200 99.0800 3370.4200 100.1600 ;
      RECT 3307.6200 99.0800 3361.1200 100.1600 ;
      RECT 2494.8200 99.0800 3305.4200 100.1600 ;
      RECT 2449.0800 99.0800 2492.6200 100.1600 ;
      RECT 2388.9400 99.0800 2446.8800 100.1600 ;
      RECT 2168.7200 99.0800 2386.7400 100.1600 ;
      RECT 1948.5000 99.0800 2166.5200 100.1600 ;
      RECT 1728.2800 99.0800 1946.3000 100.1600 ;
      RECT 1508.0600 99.0800 1726.0800 100.1600 ;
      RECT 1287.9800 99.0800 1505.8600 100.1600 ;
      RECT 1067.7600 99.0800 1285.6400 100.1600 ;
      RECT 9.3000 99.0800 1065.5600 100.1600 ;
      RECT 0.0000 99.0800 5.7000 100.1600 ;
      RECT 0.0000 97.4400 3370.4200 99.0800 ;
      RECT 0.0000 97.1000 1.7000 97.4400 ;
      RECT 3368.7200 96.3600 3370.4200 97.4400 ;
      RECT 3305.0200 96.3600 3365.1200 97.4400 ;
      RECT 2497.4200 96.3600 3302.8200 97.4400 ;
      RECT 2446.4800 96.3600 2495.2200 97.4400 ;
      RECT 2386.3400 96.3600 2444.2800 97.4400 ;
      RECT 2166.1200 96.3600 2384.1400 97.4400 ;
      RECT 1945.9000 96.3600 2163.9200 97.4400 ;
      RECT 1725.6800 96.3600 1943.7000 97.4400 ;
      RECT 1505.4600 96.3600 1723.4800 97.4400 ;
      RECT 1285.3800 96.3600 1503.2600 97.4400 ;
      RECT 1065.1600 96.3600 1283.0400 97.4400 ;
      RECT 5.3000 96.3600 1062.9600 97.4400 ;
      RECT 1.1000 96.3600 1.7000 97.1000 ;
      RECT 1.1000 96.2000 3370.4200 96.3600 ;
      RECT 0.0000 94.7200 3370.4200 96.2000 ;
      RECT 3364.7200 93.6400 3370.4200 94.7200 ;
      RECT 3307.6200 93.6400 3361.1200 94.7200 ;
      RECT 2494.8200 93.6400 3305.4200 94.7200 ;
      RECT 2449.0800 93.6400 2492.6200 94.7200 ;
      RECT 2388.9400 93.6400 2446.8800 94.7200 ;
      RECT 2168.7200 93.6400 2386.7400 94.7200 ;
      RECT 1948.5000 93.6400 2166.5200 94.7200 ;
      RECT 1728.2800 93.6400 1946.3000 94.7200 ;
      RECT 1508.0600 93.6400 1726.0800 94.7200 ;
      RECT 1287.9800 93.6400 1505.8600 94.7200 ;
      RECT 1067.7600 93.6400 1285.6400 94.7200 ;
      RECT 9.3000 93.6400 1065.5600 94.7200 ;
      RECT 0.0000 93.6400 5.7000 94.7200 ;
      RECT 0.0000 92.0000 3370.4200 93.6400 ;
      RECT 3368.7200 90.9200 3370.4200 92.0000 ;
      RECT 3305.0200 90.9200 3365.1200 92.0000 ;
      RECT 2497.4200 90.9200 3302.8200 92.0000 ;
      RECT 2446.4800 90.9200 2495.2200 92.0000 ;
      RECT 2386.3400 90.9200 2444.2800 92.0000 ;
      RECT 2166.1200 90.9200 2384.1400 92.0000 ;
      RECT 1945.9000 90.9200 2163.9200 92.0000 ;
      RECT 1725.6800 90.9200 1943.7000 92.0000 ;
      RECT 1505.4600 90.9200 1723.4800 92.0000 ;
      RECT 1285.3800 90.9200 1503.2600 92.0000 ;
      RECT 1065.1600 90.9200 1283.0400 92.0000 ;
      RECT 5.3000 90.9200 1062.9600 92.0000 ;
      RECT 0.0000 90.9200 1.7000 92.0000 ;
      RECT 0.0000 89.2800 3370.4200 90.9200 ;
      RECT 3364.7200 88.2000 3370.4200 89.2800 ;
      RECT 3307.6200 88.2000 3361.1200 89.2800 ;
      RECT 2494.8200 88.2000 3305.4200 89.2800 ;
      RECT 2449.0800 88.2000 2492.6200 89.2800 ;
      RECT 2388.9400 88.2000 2446.8800 89.2800 ;
      RECT 2168.7200 88.2000 2386.7400 89.2800 ;
      RECT 1948.5000 88.2000 2166.5200 89.2800 ;
      RECT 1728.2800 88.2000 1946.3000 89.2800 ;
      RECT 1508.0600 88.2000 1726.0800 89.2800 ;
      RECT 1287.9800 88.2000 1505.8600 89.2800 ;
      RECT 1067.7600 88.2000 1285.6400 89.2800 ;
      RECT 9.3000 88.2000 1065.5600 89.2800 ;
      RECT 0.0000 88.2000 5.7000 89.2800 ;
      RECT 0.0000 86.5600 3370.4200 88.2000 ;
      RECT 0.0000 86.1200 1.7000 86.5600 ;
      RECT 3368.7200 85.4800 3370.4200 86.5600 ;
      RECT 3305.0200 85.4800 3365.1200 86.5600 ;
      RECT 2497.4200 85.4800 3302.8200 86.5600 ;
      RECT 2446.4800 85.4800 2495.2200 86.5600 ;
      RECT 2386.3400 85.4800 2444.2800 86.5600 ;
      RECT 2166.1200 85.4800 2384.1400 86.5600 ;
      RECT 1945.9000 85.4800 2163.9200 86.5600 ;
      RECT 1725.6800 85.4800 1943.7000 86.5600 ;
      RECT 1505.4600 85.4800 1723.4800 86.5600 ;
      RECT 1285.3800 85.4800 1503.2600 86.5600 ;
      RECT 1065.1600 85.4800 1283.0400 86.5600 ;
      RECT 5.3000 85.4800 1062.9600 86.5600 ;
      RECT 1.1000 85.4800 1.7000 86.1200 ;
      RECT 1.1000 85.2200 3370.4200 85.4800 ;
      RECT 0.0000 83.8400 3370.4200 85.2200 ;
      RECT 3364.7200 82.7600 3370.4200 83.8400 ;
      RECT 3307.6200 82.7600 3361.1200 83.8400 ;
      RECT 2494.8200 82.7600 3305.4200 83.8400 ;
      RECT 2449.0800 82.7600 2492.6200 83.8400 ;
      RECT 2388.9400 82.7600 2446.8800 83.8400 ;
      RECT 2168.7200 82.7600 2386.7400 83.8400 ;
      RECT 1948.5000 82.7600 2166.5200 83.8400 ;
      RECT 1728.2800 82.7600 1946.3000 83.8400 ;
      RECT 1508.0600 82.7600 1726.0800 83.8400 ;
      RECT 1287.9800 82.7600 1505.8600 83.8400 ;
      RECT 1067.7600 82.7600 1285.6400 83.8400 ;
      RECT 9.3000 82.7600 1065.5600 83.8400 ;
      RECT 0.0000 82.7600 5.7000 83.8400 ;
      RECT 0.0000 81.1200 3370.4200 82.7600 ;
      RECT 3368.7200 80.0400 3370.4200 81.1200 ;
      RECT 3305.0200 80.0400 3365.1200 81.1200 ;
      RECT 2497.4200 80.0400 3302.8200 81.1200 ;
      RECT 2446.4800 80.0400 2495.2200 81.1200 ;
      RECT 2386.3400 80.0400 2444.2800 81.1200 ;
      RECT 2166.1200 80.0400 2384.1400 81.1200 ;
      RECT 1945.9000 80.0400 2163.9200 81.1200 ;
      RECT 1725.6800 80.0400 1943.7000 81.1200 ;
      RECT 1505.4600 80.0400 1723.4800 81.1200 ;
      RECT 1285.3800 80.0400 1503.2600 81.1200 ;
      RECT 1065.1600 80.0400 1283.0400 81.1200 ;
      RECT 5.3000 80.0400 1062.9600 81.1200 ;
      RECT 0.0000 80.0400 1.7000 81.1200 ;
      RECT 0.0000 78.4000 3370.4200 80.0400 ;
      RECT 3364.7200 77.3200 3370.4200 78.4000 ;
      RECT 3307.6200 77.3200 3361.1200 78.4000 ;
      RECT 2494.8200 77.3200 3305.4200 78.4000 ;
      RECT 2449.0800 77.3200 2492.6200 78.4000 ;
      RECT 2388.9400 77.3200 2446.8800 78.4000 ;
      RECT 2168.7200 77.3200 2386.7400 78.4000 ;
      RECT 1948.5000 77.3200 2166.5200 78.4000 ;
      RECT 1728.2800 77.3200 1946.3000 78.4000 ;
      RECT 1508.0600 77.3200 1726.0800 78.4000 ;
      RECT 1287.9800 77.3200 1505.8600 78.4000 ;
      RECT 1067.7600 77.3200 1285.6400 78.4000 ;
      RECT 9.3000 77.3200 1065.5600 78.4000 ;
      RECT 0.0000 77.3200 5.7000 78.4000 ;
      RECT 0.0000 75.7500 3370.4200 77.3200 ;
      RECT 1.1000 75.6800 3370.4200 75.7500 ;
      RECT 1.1000 74.8500 1.7000 75.6800 ;
      RECT 3368.7200 74.6000 3370.4200 75.6800 ;
      RECT 3305.0200 74.6000 3365.1200 75.6800 ;
      RECT 2497.4200 74.6000 3302.8200 75.6800 ;
      RECT 2446.4800 74.6000 2495.2200 75.6800 ;
      RECT 2386.3400 74.6000 2444.2800 75.6800 ;
      RECT 2166.1200 74.6000 2384.1400 75.6800 ;
      RECT 1945.9000 74.6000 2163.9200 75.6800 ;
      RECT 1725.6800 74.6000 1943.7000 75.6800 ;
      RECT 1505.4600 74.6000 1723.4800 75.6800 ;
      RECT 1285.3800 74.6000 1503.2600 75.6800 ;
      RECT 1065.1600 74.6000 1283.0400 75.6800 ;
      RECT 5.3000 74.6000 1062.9600 75.6800 ;
      RECT 0.0000 74.6000 1.7000 74.8500 ;
      RECT 0.0000 72.9600 3370.4200 74.6000 ;
      RECT 3364.7200 71.8800 3370.4200 72.9600 ;
      RECT 3307.6200 71.8800 3361.1200 72.9600 ;
      RECT 2494.8200 71.8800 3305.4200 72.9600 ;
      RECT 2449.0800 71.8800 2492.6200 72.9600 ;
      RECT 2388.9400 71.8800 2446.8800 72.9600 ;
      RECT 2168.7200 71.8800 2386.7400 72.9600 ;
      RECT 1948.5000 71.8800 2166.5200 72.9600 ;
      RECT 1728.2800 71.8800 1946.3000 72.9600 ;
      RECT 1508.0600 71.8800 1726.0800 72.9600 ;
      RECT 1287.9800 71.8800 1505.8600 72.9600 ;
      RECT 1067.7600 71.8800 1285.6400 72.9600 ;
      RECT 9.3000 71.8800 1065.5600 72.9600 ;
      RECT 0.0000 71.8800 5.7000 72.9600 ;
      RECT 0.0000 70.2400 3370.4200 71.8800 ;
      RECT 3368.7200 69.1600 3370.4200 70.2400 ;
      RECT 3305.0200 69.1600 3365.1200 70.2400 ;
      RECT 2497.4200 69.1600 3302.8200 70.2400 ;
      RECT 2446.4800 69.1600 2495.2200 70.2400 ;
      RECT 2386.3400 69.1600 2444.2800 70.2400 ;
      RECT 2166.1200 69.1600 2384.1400 70.2400 ;
      RECT 1945.9000 69.1600 2163.9200 70.2400 ;
      RECT 1725.6800 69.1600 1943.7000 70.2400 ;
      RECT 1505.4600 69.1600 1723.4800 70.2400 ;
      RECT 1285.3800 69.1600 1503.2600 70.2400 ;
      RECT 1065.1600 69.1600 1283.0400 70.2400 ;
      RECT 5.3000 69.1600 1062.9600 70.2400 ;
      RECT 0.0000 69.1600 1.7000 70.2400 ;
      RECT 0.0000 67.5200 3370.4200 69.1600 ;
      RECT 3364.7200 66.4400 3370.4200 67.5200 ;
      RECT 3307.6200 66.4400 3361.1200 67.5200 ;
      RECT 2494.8200 66.4400 3305.4200 67.5200 ;
      RECT 2449.0800 66.4400 2492.6200 67.5200 ;
      RECT 2388.9400 66.4400 2446.8800 67.5200 ;
      RECT 2168.7200 66.4400 2386.7400 67.5200 ;
      RECT 1948.5000 66.4400 2166.5200 67.5200 ;
      RECT 1728.2800 66.4400 1946.3000 67.5200 ;
      RECT 1508.0600 66.4400 1726.0800 67.5200 ;
      RECT 1287.9800 66.4400 1505.8600 67.5200 ;
      RECT 1067.7600 66.4400 1285.6400 67.5200 ;
      RECT 9.3000 66.4400 1065.5600 67.5200 ;
      RECT 0.0000 66.4400 5.7000 67.5200 ;
      RECT 0.0000 64.8000 3370.4200 66.4400 ;
      RECT 0.0000 64.7700 1.7000 64.8000 ;
      RECT 1.1000 63.8700 1.7000 64.7700 ;
      RECT 3368.7200 63.7200 3370.4200 64.8000 ;
      RECT 3305.0200 63.7200 3365.1200 64.8000 ;
      RECT 2497.4200 63.7200 3302.8200 64.8000 ;
      RECT 2446.4800 63.7200 2495.2200 64.8000 ;
      RECT 2386.3400 63.7200 2444.2800 64.8000 ;
      RECT 2166.1200 63.7200 2384.1400 64.8000 ;
      RECT 1945.9000 63.7200 2163.9200 64.8000 ;
      RECT 1725.6800 63.7200 1943.7000 64.8000 ;
      RECT 1505.4600 63.7200 1723.4800 64.8000 ;
      RECT 1285.3800 63.7200 1503.2600 64.8000 ;
      RECT 1065.1600 63.7200 1283.0400 64.8000 ;
      RECT 5.3000 63.7200 1062.9600 64.8000 ;
      RECT 0.0000 63.7200 1.7000 63.8700 ;
      RECT 0.0000 62.0800 3370.4200 63.7200 ;
      RECT 3364.7200 61.0000 3370.4200 62.0800 ;
      RECT 3307.6200 61.0000 3361.1200 62.0800 ;
      RECT 2494.8200 61.0000 3305.4200 62.0800 ;
      RECT 2449.0800 61.0000 2492.6200 62.0800 ;
      RECT 2388.9400 61.0000 2446.8800 62.0800 ;
      RECT 2168.7200 61.0000 2386.7400 62.0800 ;
      RECT 1948.5000 61.0000 2166.5200 62.0800 ;
      RECT 1728.2800 61.0000 1946.3000 62.0800 ;
      RECT 1508.0600 61.0000 1726.0800 62.0800 ;
      RECT 1287.9800 61.0000 1505.8600 62.0800 ;
      RECT 1067.7600 61.0000 1285.6400 62.0800 ;
      RECT 9.3000 61.0000 1065.5600 62.0800 ;
      RECT 0.0000 61.0000 5.7000 62.0800 ;
      RECT 0.0000 59.3600 3370.4200 61.0000 ;
      RECT 3368.7200 58.2800 3370.4200 59.3600 ;
      RECT 3305.0200 58.2800 3365.1200 59.3600 ;
      RECT 2497.4200 58.2800 3302.8200 59.3600 ;
      RECT 2446.4800 58.2800 2495.2200 59.3600 ;
      RECT 2386.3400 58.2800 2444.2800 59.3600 ;
      RECT 2166.1200 58.2800 2384.1400 59.3600 ;
      RECT 1945.9000 58.2800 2163.9200 59.3600 ;
      RECT 1725.6800 58.2800 1943.7000 59.3600 ;
      RECT 1505.4600 58.2800 1723.4800 59.3600 ;
      RECT 1285.3800 58.2800 1503.2600 59.3600 ;
      RECT 1065.1600 58.2800 1283.0400 59.3600 ;
      RECT 5.3000 58.2800 1062.9600 59.3600 ;
      RECT 0.0000 58.2800 1.7000 59.3600 ;
      RECT 0.0000 56.6400 3370.4200 58.2800 ;
      RECT 3364.7200 55.5600 3370.4200 56.6400 ;
      RECT 3307.6200 55.5600 3361.1200 56.6400 ;
      RECT 2494.8200 55.5600 3305.4200 56.6400 ;
      RECT 2449.0800 55.5600 2492.6200 56.6400 ;
      RECT 2388.9400 55.5600 2446.8800 56.6400 ;
      RECT 2168.7200 55.5600 2386.7400 56.6400 ;
      RECT 1948.5000 55.5600 2166.5200 56.6400 ;
      RECT 1728.2800 55.5600 1946.3000 56.6400 ;
      RECT 1508.0600 55.5600 1726.0800 56.6400 ;
      RECT 1287.9800 55.5600 1505.8600 56.6400 ;
      RECT 1067.7600 55.5600 1285.6400 56.6400 ;
      RECT 9.3000 55.5600 1065.5600 56.6400 ;
      RECT 0.0000 55.5600 5.7000 56.6400 ;
      RECT 0.0000 53.9200 3370.4200 55.5600 ;
      RECT 0.0000 53.7900 1.7000 53.9200 ;
      RECT 1.1000 52.8900 1.7000 53.7900 ;
      RECT 3368.7200 52.8400 3370.4200 53.9200 ;
      RECT 3305.0200 52.8400 3365.1200 53.9200 ;
      RECT 2497.4200 52.8400 3302.8200 53.9200 ;
      RECT 2446.4800 52.8400 2495.2200 53.9200 ;
      RECT 2386.3400 52.8400 2444.2800 53.9200 ;
      RECT 2166.1200 52.8400 2384.1400 53.9200 ;
      RECT 1945.9000 52.8400 2163.9200 53.9200 ;
      RECT 1725.6800 52.8400 1943.7000 53.9200 ;
      RECT 1505.4600 52.8400 1723.4800 53.9200 ;
      RECT 1285.3800 52.8400 1503.2600 53.9200 ;
      RECT 1065.1600 52.8400 1283.0400 53.9200 ;
      RECT 5.3000 52.8400 1062.9600 53.9200 ;
      RECT 0.0000 52.8400 1.7000 52.8900 ;
      RECT 0.0000 51.2000 3370.4200 52.8400 ;
      RECT 3364.7200 50.1200 3370.4200 51.2000 ;
      RECT 3307.6200 50.1200 3361.1200 51.2000 ;
      RECT 2494.8200 50.1200 3305.4200 51.2000 ;
      RECT 2449.0800 50.1200 2492.6200 51.2000 ;
      RECT 2388.9400 50.1200 2446.8800 51.2000 ;
      RECT 2168.7200 50.1200 2386.7400 51.2000 ;
      RECT 1948.5000 50.1200 2166.5200 51.2000 ;
      RECT 1728.2800 50.1200 1946.3000 51.2000 ;
      RECT 1508.0600 50.1200 1726.0800 51.2000 ;
      RECT 1287.9800 50.1200 1505.8600 51.2000 ;
      RECT 1067.7600 50.1200 1285.6400 51.2000 ;
      RECT 9.3000 50.1200 1065.5600 51.2000 ;
      RECT 0.0000 50.1200 5.7000 51.2000 ;
      RECT 0.0000 48.4800 3370.4200 50.1200 ;
      RECT 3368.7200 47.4000 3370.4200 48.4800 ;
      RECT 3305.0200 47.4000 3365.1200 48.4800 ;
      RECT 2497.4200 47.4000 3302.8200 48.4800 ;
      RECT 2446.4800 47.4000 2495.2200 48.4800 ;
      RECT 2386.3400 47.4000 2444.2800 48.4800 ;
      RECT 2166.1200 47.4000 2384.1400 48.4800 ;
      RECT 1945.9000 47.4000 2163.9200 48.4800 ;
      RECT 1725.6800 47.4000 1943.7000 48.4800 ;
      RECT 1505.4600 47.4000 1723.4800 48.4800 ;
      RECT 1285.3800 47.4000 1503.2600 48.4800 ;
      RECT 1065.1600 47.4000 1283.0400 48.4800 ;
      RECT 5.3000 47.4000 1062.9600 48.4800 ;
      RECT 0.0000 47.4000 1.7000 48.4800 ;
      RECT 0.0000 45.7600 3370.4200 47.4000 ;
      RECT 3364.7200 44.6800 3370.4200 45.7600 ;
      RECT 3307.6200 44.6800 3361.1200 45.7600 ;
      RECT 2494.8200 44.6800 3305.4200 45.7600 ;
      RECT 2449.0800 44.6800 2492.6200 45.7600 ;
      RECT 2388.9400 44.6800 2446.8800 45.7600 ;
      RECT 2168.7200 44.6800 2386.7400 45.7600 ;
      RECT 1948.5000 44.6800 2166.5200 45.7600 ;
      RECT 1728.2800 44.6800 1946.3000 45.7600 ;
      RECT 1508.0600 44.6800 1726.0800 45.7600 ;
      RECT 1287.9800 44.6800 1505.8600 45.7600 ;
      RECT 1067.7600 44.6800 1285.6400 45.7600 ;
      RECT 9.3000 44.6800 1065.5600 45.7600 ;
      RECT 0.0000 44.6800 5.7000 45.7600 ;
      RECT 0.0000 43.0400 3370.4200 44.6800 ;
      RECT 0.0000 42.8100 1.7000 43.0400 ;
      RECT 3368.7200 41.9600 3370.4200 43.0400 ;
      RECT 3305.0200 41.9600 3365.1200 43.0400 ;
      RECT 2497.4200 41.9600 3302.8200 43.0400 ;
      RECT 2446.4800 41.9600 2495.2200 43.0400 ;
      RECT 2386.3400 41.9600 2444.2800 43.0400 ;
      RECT 2166.1200 41.9600 2384.1400 43.0400 ;
      RECT 1945.9000 41.9600 2163.9200 43.0400 ;
      RECT 1725.6800 41.9600 1943.7000 43.0400 ;
      RECT 1505.4600 41.9600 1723.4800 43.0400 ;
      RECT 1285.3800 41.9600 1503.2600 43.0400 ;
      RECT 1065.1600 41.9600 1283.0400 43.0400 ;
      RECT 5.3000 41.9600 1062.9600 43.0400 ;
      RECT 1.1000 41.9600 1.7000 42.8100 ;
      RECT 1.1000 41.9100 3370.4200 41.9600 ;
      RECT 0.0000 40.3200 3370.4200 41.9100 ;
      RECT 3364.7200 39.2400 3370.4200 40.3200 ;
      RECT 3307.6200 39.2400 3361.1200 40.3200 ;
      RECT 2494.8200 39.2400 3305.4200 40.3200 ;
      RECT 2449.0800 39.2400 2492.6200 40.3200 ;
      RECT 2388.9400 39.2400 2446.8800 40.3200 ;
      RECT 2168.7200 39.2400 2386.7400 40.3200 ;
      RECT 1948.5000 39.2400 2166.5200 40.3200 ;
      RECT 1728.2800 39.2400 1946.3000 40.3200 ;
      RECT 1508.0600 39.2400 1726.0800 40.3200 ;
      RECT 1287.9800 39.2400 1505.8600 40.3200 ;
      RECT 1067.7600 39.2400 1285.6400 40.3200 ;
      RECT 9.3000 39.2400 1065.5600 40.3200 ;
      RECT 0.0000 39.2400 5.7000 40.3200 ;
      RECT 0.0000 37.6000 3370.4200 39.2400 ;
      RECT 3368.7200 36.5200 3370.4200 37.6000 ;
      RECT 3305.0200 36.5200 3365.1200 37.6000 ;
      RECT 2497.4200 36.5200 3302.8200 37.6000 ;
      RECT 2446.4800 36.5200 2495.2200 37.6000 ;
      RECT 2386.3400 36.5200 2444.2800 37.6000 ;
      RECT 2166.1200 36.5200 2384.1400 37.6000 ;
      RECT 1945.9000 36.5200 2163.9200 37.6000 ;
      RECT 1725.6800 36.5200 1943.7000 37.6000 ;
      RECT 1505.4600 36.5200 1723.4800 37.6000 ;
      RECT 1285.3800 36.5200 1503.2600 37.6000 ;
      RECT 1065.1600 36.5200 1283.0400 37.6000 ;
      RECT 5.3000 36.5200 1062.9600 37.6000 ;
      RECT 0.0000 36.5200 1.7000 37.6000 ;
      RECT 0.0000 34.8800 3370.4200 36.5200 ;
      RECT 3364.7200 33.8000 3370.4200 34.8800 ;
      RECT 3307.6200 33.8000 3361.1200 34.8800 ;
      RECT 2494.8200 33.8000 3305.4200 34.8800 ;
      RECT 2449.0800 33.8000 2492.6200 34.8800 ;
      RECT 2388.9400 33.8000 2446.8800 34.8800 ;
      RECT 2168.7200 33.8000 2386.7400 34.8800 ;
      RECT 1948.5000 33.8000 2166.5200 34.8800 ;
      RECT 1728.2800 33.8000 1946.3000 34.8800 ;
      RECT 1508.0600 33.8000 1726.0800 34.8800 ;
      RECT 1287.9800 33.8000 1505.8600 34.8800 ;
      RECT 1067.7600 33.8000 1285.6400 34.8800 ;
      RECT 9.3000 33.8000 1065.5600 34.8800 ;
      RECT 0.0000 33.8000 5.7000 34.8800 ;
      RECT 0.0000 32.1600 3370.4200 33.8000 ;
      RECT 0.0000 31.8300 1.7000 32.1600 ;
      RECT 3368.7200 31.0800 3370.4200 32.1600 ;
      RECT 3305.0200 31.0800 3365.1200 32.1600 ;
      RECT 2497.4200 31.0800 3302.8200 32.1600 ;
      RECT 2446.4800 31.0800 2495.2200 32.1600 ;
      RECT 2386.3400 31.0800 2444.2800 32.1600 ;
      RECT 2166.1200 31.0800 2384.1400 32.1600 ;
      RECT 1945.9000 31.0800 2163.9200 32.1600 ;
      RECT 1725.6800 31.0800 1943.7000 32.1600 ;
      RECT 1505.4600 31.0800 1723.4800 32.1600 ;
      RECT 1285.3800 31.0800 1503.2600 32.1600 ;
      RECT 1065.1600 31.0800 1283.0400 32.1600 ;
      RECT 5.3000 31.0800 1062.9600 32.1600 ;
      RECT 1.1000 31.0800 1.7000 31.8300 ;
      RECT 1.1000 30.9300 3370.4200 31.0800 ;
      RECT 0.0000 29.4400 3370.4200 30.9300 ;
      RECT 3364.7200 28.3600 3370.4200 29.4400 ;
      RECT 3307.6200 28.3600 3361.1200 29.4400 ;
      RECT 2494.8200 28.3600 3305.4200 29.4400 ;
      RECT 2449.0800 28.3600 2492.6200 29.4400 ;
      RECT 2388.9400 28.3600 2446.8800 29.4400 ;
      RECT 2168.7200 28.3600 2386.7400 29.4400 ;
      RECT 1948.5000 28.3600 2166.5200 29.4400 ;
      RECT 1728.2800 28.3600 1946.3000 29.4400 ;
      RECT 1508.0600 28.3600 1726.0800 29.4400 ;
      RECT 1287.9800 28.3600 1505.8600 29.4400 ;
      RECT 1067.7600 28.3600 1285.6400 29.4400 ;
      RECT 9.3000 28.3600 1065.5600 29.4400 ;
      RECT 0.0000 28.3600 5.7000 29.4400 ;
      RECT 0.0000 26.7200 3370.4200 28.3600 ;
      RECT 3368.7200 25.6400 3370.4200 26.7200 ;
      RECT 3305.0200 25.6400 3365.1200 26.7200 ;
      RECT 2497.4200 25.6400 3302.8200 26.7200 ;
      RECT 2446.4800 25.6400 2495.2200 26.7200 ;
      RECT 2386.3400 25.6400 2444.2800 26.7200 ;
      RECT 2166.1200 25.6400 2384.1400 26.7200 ;
      RECT 1945.9000 25.6400 2163.9200 26.7200 ;
      RECT 1725.6800 25.6400 1943.7000 26.7200 ;
      RECT 1505.4600 25.6400 1723.4800 26.7200 ;
      RECT 1285.3800 25.6400 1503.2600 26.7200 ;
      RECT 1065.1600 25.6400 1283.0400 26.7200 ;
      RECT 5.3000 25.6400 1062.9600 26.7200 ;
      RECT 0.0000 25.6400 1.7000 26.7200 ;
      RECT 0.0000 24.0000 3370.4200 25.6400 ;
      RECT 3364.7200 22.9200 3370.4200 24.0000 ;
      RECT 3307.6200 22.9200 3361.1200 24.0000 ;
      RECT 2494.8200 22.9200 3305.4200 24.0000 ;
      RECT 2449.0800 22.9200 2492.6200 24.0000 ;
      RECT 2388.9400 22.9200 2446.8800 24.0000 ;
      RECT 2168.7200 22.9200 2386.7400 24.0000 ;
      RECT 1948.5000 22.9200 2166.5200 24.0000 ;
      RECT 1728.2800 22.9200 1946.3000 24.0000 ;
      RECT 1508.0600 22.9200 1726.0800 24.0000 ;
      RECT 1287.9800 22.9200 1505.8600 24.0000 ;
      RECT 1067.7600 22.9200 1285.6400 24.0000 ;
      RECT 9.3000 22.9200 1065.5600 24.0000 ;
      RECT 0.0000 22.9200 5.7000 24.0000 ;
      RECT 0.0000 21.2800 3370.4200 22.9200 ;
      RECT 0.0000 20.8500 1.7000 21.2800 ;
      RECT 3368.7200 20.2000 3370.4200 21.2800 ;
      RECT 3305.0200 20.2000 3365.1200 21.2800 ;
      RECT 2497.4200 20.2000 3302.8200 21.2800 ;
      RECT 2446.4800 20.2000 2495.2200 21.2800 ;
      RECT 2386.3400 20.2000 2444.2800 21.2800 ;
      RECT 2166.1200 20.2000 2384.1400 21.2800 ;
      RECT 1945.9000 20.2000 2163.9200 21.2800 ;
      RECT 1725.6800 20.2000 1943.7000 21.2800 ;
      RECT 1505.4600 20.2000 1723.4800 21.2800 ;
      RECT 1285.3800 20.2000 1503.2600 21.2800 ;
      RECT 1065.1600 20.2000 1283.0400 21.2800 ;
      RECT 5.3000 20.2000 1062.9600 21.2800 ;
      RECT 1.1000 20.2000 1.7000 20.8500 ;
      RECT 1.1000 19.9500 3370.4200 20.2000 ;
      RECT 0.0000 18.5600 3370.4200 19.9500 ;
      RECT 3364.7200 17.4800 3370.4200 18.5600 ;
      RECT 3307.6200 17.4800 3361.1200 18.5600 ;
      RECT 2494.8200 17.4800 3305.4200 18.5600 ;
      RECT 2449.0800 17.4800 2492.6200 18.5600 ;
      RECT 2388.9400 17.4800 2446.8800 18.5600 ;
      RECT 2168.7200 17.4800 2386.7400 18.5600 ;
      RECT 1948.5000 17.4800 2166.5200 18.5600 ;
      RECT 1728.2800 17.4800 1946.3000 18.5600 ;
      RECT 1508.0600 17.4800 1726.0800 18.5600 ;
      RECT 1287.9800 17.4800 1505.8600 18.5600 ;
      RECT 1067.7600 17.4800 1285.6400 18.5600 ;
      RECT 9.3000 17.4800 1065.5600 18.5600 ;
      RECT 0.0000 17.4800 5.7000 18.5600 ;
      RECT 0.0000 15.8400 3370.4200 17.4800 ;
      RECT 3368.7200 14.7600 3370.4200 15.8400 ;
      RECT 3305.0200 14.7600 3365.1200 15.8400 ;
      RECT 2497.4200 14.7600 3302.8200 15.8400 ;
      RECT 2446.4800 14.7600 2495.2200 15.8400 ;
      RECT 2386.3400 14.7600 2444.2800 15.8400 ;
      RECT 2166.1200 14.7600 2384.1400 15.8400 ;
      RECT 1945.9000 14.7600 2163.9200 15.8400 ;
      RECT 1725.6800 14.7600 1943.7000 15.8400 ;
      RECT 1505.4600 14.7600 1723.4800 15.8400 ;
      RECT 1285.3800 14.7600 1503.2600 15.8400 ;
      RECT 1065.1600 14.7600 1283.0400 15.8400 ;
      RECT 5.3000 14.7600 1062.9600 15.8400 ;
      RECT 0.0000 14.7600 1.7000 15.8400 ;
      RECT 0.0000 13.1200 3370.4200 14.7600 ;
      RECT 3364.7200 12.0400 3370.4200 13.1200 ;
      RECT 3307.6200 12.0400 3361.1200 13.1200 ;
      RECT 2494.8200 12.0400 3305.4200 13.1200 ;
      RECT 2449.0800 12.0400 2492.6200 13.1200 ;
      RECT 2388.9400 12.0400 2446.8800 13.1200 ;
      RECT 2168.7200 12.0400 2386.7400 13.1200 ;
      RECT 1948.5000 12.0400 2166.5200 13.1200 ;
      RECT 1728.2800 12.0400 1946.3000 13.1200 ;
      RECT 1508.0600 12.0400 1726.0800 13.1200 ;
      RECT 1287.9800 12.0400 1505.8600 13.1200 ;
      RECT 1067.7600 12.0400 1285.6400 13.1200 ;
      RECT 9.3000 12.0400 1065.5600 13.1200 ;
      RECT 0.0000 12.0400 5.7000 13.1200 ;
      RECT 0.0000 11.0000 3370.4200 12.0400 ;
      RECT 1065.0600 10.4000 3370.4200 11.0000 ;
      RECT 0.0000 10.4000 1062.6600 11.0000 ;
      RECT 3368.7200 9.3200 3370.4200 10.4000 ;
      RECT 3305.0200 9.3200 3365.1200 10.4000 ;
      RECT 2497.4200 9.3200 3302.8200 10.4000 ;
      RECT 2446.4800 9.3200 2495.2200 10.4000 ;
      RECT 2386.3400 9.3200 2444.2800 10.4000 ;
      RECT 2166.1200 9.3200 2384.1400 10.4000 ;
      RECT 1945.9000 9.3200 2163.9200 10.4000 ;
      RECT 1725.6800 9.3200 1943.7000 10.4000 ;
      RECT 1505.4600 9.3200 1723.4800 10.4000 ;
      RECT 1285.3800 9.3200 1503.2600 10.4000 ;
      RECT 1065.0600 9.3200 1283.0400 10.4000 ;
      RECT 5.3000 9.3200 1062.6600 10.4000 ;
      RECT 0.0000 9.3200 1.7000 10.4000 ;
      RECT 1065.0600 9.3000 3370.4200 9.3200 ;
      RECT 0.0000 9.3000 1062.6600 9.3200 ;
      RECT 3364.7200 5.7000 3370.4200 9.3000 ;
      RECT 0.0000 5.7000 5.7000 9.3000 ;
      RECT 1065.0600 5.6000 3370.4200 5.7000 ;
      RECT 0.0000 5.6000 1062.6600 5.7000 ;
      RECT 0.0000 5.3000 3370.4200 5.6000 ;
      RECT 3368.7200 1.7000 3370.4200 5.3000 ;
      RECT 0.0000 1.7000 1.7000 5.3000 ;
      RECT 0.0000 0.0000 3370.4200 1.7000 ;
    LAYER met4 ;
      RECT 0.0000 2568.0200 3370.4200 2569.7200 ;
      RECT 3305.0200 2564.0200 3365.1200 2568.0200 ;
      RECT 2446.4800 2564.0200 2495.2200 2568.0200 ;
      RECT 2436.3200 2564.0200 2444.2800 2568.0200 ;
      RECT 2386.3400 2564.0200 2396.7000 2568.0200 ;
      RECT 2376.2800 2564.0200 2384.1400 2568.0200 ;
      RECT 2166.1200 2564.0200 2176.3800 2568.0200 ;
      RECT 2156.0600 2564.0200 2163.9200 2568.0200 ;
      RECT 1945.9000 2564.0200 1956.1600 2568.0200 ;
      RECT 1935.8400 2564.0200 1943.7000 2568.0200 ;
      RECT 1725.6800 2564.0200 1735.9400 2568.0200 ;
      RECT 1715.6200 2564.0200 1723.4800 2568.0200 ;
      RECT 1505.4600 2564.0200 1515.7200 2568.0200 ;
      RECT 1495.4000 2564.0200 1503.2600 2568.0200 ;
      RECT 1285.3800 2564.0200 1295.5000 2568.0200 ;
      RECT 1275.1800 2564.0200 1283.0400 2568.0200 ;
      RECT 1065.1600 2564.0200 1075.2800 2568.0200 ;
      RECT 1055.1000 2564.0200 1062.9600 2568.0200 ;
      RECT 1007.4200 2564.0200 1015.2800 2568.0200 ;
      RECT 5.3000 2564.0200 1005.2200 2568.0200 ;
      RECT 2378.6800 2508.7600 2384.1400 2564.0200 ;
      RECT 2376.2800 2508.7600 2376.4800 2564.0200 ;
      RECT 2178.5800 2508.7600 2374.0800 2568.0200 ;
      RECT 2176.1800 2508.7600 2176.3800 2564.0200 ;
      RECT 2168.7200 2508.7600 2173.9800 2564.0200 ;
      RECT 2158.4600 2508.7600 2163.9200 2564.0200 ;
      RECT 2156.0600 2508.7600 2156.2600 2564.0200 ;
      RECT 1958.3600 2508.7600 2153.8600 2568.0200 ;
      RECT 1955.9600 2508.7600 1956.1600 2564.0200 ;
      RECT 1948.5000 2508.7600 1953.7600 2564.0200 ;
      RECT 1938.2400 2508.7600 1943.7000 2564.0200 ;
      RECT 1935.8400 2508.7600 1936.0400 2564.0200 ;
      RECT 1738.1400 2508.7600 1933.6400 2568.0200 ;
      RECT 1735.7400 2508.7600 1735.9400 2564.0200 ;
      RECT 1728.2800 2508.7600 1733.5400 2564.0200 ;
      RECT 1718.0200 2508.7600 1723.4800 2564.0200 ;
      RECT 1715.6200 2508.7600 1715.8200 2564.0200 ;
      RECT 1517.9200 2508.7600 1713.4200 2568.0200 ;
      RECT 1515.5200 2508.7600 1515.7200 2564.0200 ;
      RECT 1508.0600 2508.7600 1513.3200 2564.0200 ;
      RECT 1497.8000 2508.7600 1503.2600 2564.0200 ;
      RECT 1495.4000 2508.7600 1495.6000 2564.0200 ;
      RECT 1297.7000 2508.7600 1493.2000 2568.0200 ;
      RECT 1295.3000 2508.7600 1295.5000 2564.0200 ;
      RECT 1287.9800 2508.7600 1293.1000 2564.0200 ;
      RECT 1277.5800 2508.7600 1283.0400 2564.0200 ;
      RECT 1275.1800 2508.7600 1275.3800 2564.0200 ;
      RECT 1077.4800 2508.7600 1272.9800 2568.0200 ;
      RECT 1075.0800 2508.7600 1075.2800 2564.0200 ;
      RECT 1067.7600 2508.7600 1072.8800 2564.0200 ;
      RECT 2168.7200 2490.0000 2384.1400 2508.7600 ;
      RECT 1948.5000 2490.0000 2163.9200 2508.7600 ;
      RECT 1728.2800 2490.0000 1943.7000 2508.7600 ;
      RECT 1508.0600 2490.0000 1723.4800 2508.7600 ;
      RECT 1287.9800 2490.0000 1503.2600 2508.7600 ;
      RECT 1067.7600 2490.0000 1283.0400 2508.7600 ;
      RECT 2176.1800 2487.2800 2384.1400 2490.0000 ;
      RECT 1955.9600 2487.2800 2163.9200 2490.0000 ;
      RECT 1735.7400 2487.2800 1943.7000 2490.0000 ;
      RECT 1515.5200 2487.2800 1723.4800 2490.0000 ;
      RECT 1295.3000 2487.2800 1503.2600 2490.0000 ;
      RECT 1075.0800 2487.2800 1283.0400 2490.0000 ;
      RECT 2376.2800 2480.7000 2384.1400 2487.2800 ;
      RECT 2176.1800 2480.7000 2374.0800 2487.2800 ;
      RECT 2156.0600 2480.7000 2163.9200 2487.2800 ;
      RECT 1955.9600 2480.7000 2153.8600 2487.2800 ;
      RECT 1935.8400 2480.7000 1943.7000 2487.2800 ;
      RECT 1735.7400 2480.7000 1933.6400 2487.2800 ;
      RECT 1715.6200 2480.7000 1723.4800 2487.2800 ;
      RECT 1515.5200 2480.7000 1713.4200 2487.2800 ;
      RECT 1495.4000 2480.7000 1503.2600 2487.2800 ;
      RECT 1295.3000 2480.7000 1493.2000 2487.2800 ;
      RECT 1275.1800 2480.7000 1283.0400 2487.2800 ;
      RECT 1075.0800 2480.7000 1272.9800 2487.2800 ;
      RECT 2178.5800 2475.3300 2374.0800 2480.7000 ;
      RECT 1958.3600 2475.3300 2153.8600 2480.7000 ;
      RECT 1738.1400 2475.3300 1933.6400 2480.7000 ;
      RECT 1517.9200 2475.3300 1713.4200 2480.7000 ;
      RECT 1297.7000 2475.3300 1493.2000 2480.7000 ;
      RECT 1275.1800 2475.3300 1275.3800 2480.7000 ;
      RECT 1077.4800 2475.3300 1272.9800 2480.7000 ;
      RECT 2376.2800 2474.7000 2376.4800 2480.7000 ;
      RECT 2176.1800 2474.7000 2176.3800 2480.7000 ;
      RECT 2156.0600 2474.7000 2156.2600 2480.7000 ;
      RECT 1955.9600 2474.7000 1956.1600 2480.7000 ;
      RECT 1935.8400 2474.7000 1936.0400 2480.7000 ;
      RECT 1735.7400 2474.7000 1735.9400 2480.7000 ;
      RECT 1715.6200 2474.7000 1715.8200 2480.7000 ;
      RECT 1515.5200 2474.7000 1515.7200 2480.7000 ;
      RECT 1495.4000 2474.7000 1495.6000 2480.7000 ;
      RECT 1295.3000 2474.7000 1295.5000 2480.7000 ;
      RECT 1077.7200 2474.7000 1272.9800 2475.3300 ;
      RECT 1075.0800 2474.7000 1075.2800 2480.7000 ;
      RECT 2378.6800 2474.3000 2384.1400 2480.7000 ;
      RECT 2178.6800 2474.3000 2373.9800 2475.3300 ;
      RECT 2168.7200 2474.3000 2173.9800 2490.0000 ;
      RECT 2158.4600 2474.3000 2163.9200 2480.7000 ;
      RECT 1948.5000 2474.3000 1953.7600 2490.0000 ;
      RECT 1938.2400 2474.3000 1943.7000 2480.7000 ;
      RECT 1738.2400 2474.3000 1933.5400 2475.3300 ;
      RECT 1728.2800 2474.3000 1733.5400 2490.0000 ;
      RECT 1718.0200 2474.3000 1723.4800 2480.7000 ;
      RECT 1518.0200 2474.3000 1713.3200 2475.3300 ;
      RECT 1508.0600 2474.3000 1513.3200 2490.0000 ;
      RECT 1497.8000 2474.3000 1503.2600 2480.7000 ;
      RECT 1297.8000 2474.3000 1493.1000 2475.3300 ;
      RECT 1287.9800 2474.3000 1293.1000 2490.0000 ;
      RECT 1277.5800 2474.3000 1283.0400 2480.7000 ;
      RECT 1075.0800 2474.3000 1075.5200 2474.7000 ;
      RECT 2376.1800 2473.5200 2376.4800 2474.7000 ;
      RECT 2155.9600 2473.5200 2156.2600 2474.7000 ;
      RECT 1935.7400 2473.5200 1936.0400 2474.7000 ;
      RECT 1715.5200 2473.5200 1715.8200 2474.7000 ;
      RECT 1495.3000 2473.5200 1495.6000 2474.7000 ;
      RECT 1275.2200 2473.5200 1275.3800 2475.3300 ;
      RECT 2183.2400 2472.1000 2373.9800 2474.3000 ;
      RECT 2178.6800 2472.1000 2181.0400 2474.3000 ;
      RECT 2176.1800 2472.1000 2176.4800 2474.7000 ;
      RECT 1955.9600 2472.1000 1956.2600 2474.7000 ;
      RECT 1742.8000 2472.1000 1933.5400 2474.3000 ;
      RECT 1738.2400 2472.1000 1740.6000 2474.3000 ;
      RECT 1735.7400 2472.1000 1736.0400 2474.7000 ;
      RECT 1522.5800 2472.1000 1713.3200 2474.3000 ;
      RECT 1518.0200 2472.1000 1520.3800 2474.3000 ;
      RECT 1515.5200 2472.1000 1515.8200 2474.7000 ;
      RECT 1302.3600 2472.1000 1493.1000 2474.3000 ;
      RECT 1297.8000 2472.1000 1300.1600 2474.3000 ;
      RECT 1295.3000 2472.1000 1295.6000 2474.7000 ;
      RECT 1067.7600 2472.1000 1072.8800 2490.0000 ;
      RECT 2388.9400 2470.4600 2396.7000 2564.0200 ;
      RECT 1277.8200 2469.3000 1283.0400 2474.3000 ;
      RECT 1275.2200 2469.3000 1275.6200 2473.5200 ;
      RECT 1077.7200 2469.3000 1273.0200 2474.7000 ;
      RECT 1075.1200 2469.3000 1075.5200 2474.3000 ;
      RECT 2158.5600 2469.0400 2163.9200 2474.3000 ;
      RECT 2155.9600 2469.0400 2156.3600 2473.5200 ;
      RECT 1958.4600 2469.0400 2153.7600 2475.3300 ;
      RECT 1955.8600 2469.0400 1956.2600 2472.1000 ;
      RECT 1057.5000 2468.7600 1062.9600 2564.0200 ;
      RECT 1055.1000 2468.7600 1055.3000 2564.0200 ;
      RECT 1017.4800 2468.7600 1052.9000 2568.0200 ;
      RECT 1015.0800 2468.7600 1015.2800 2564.0200 ;
      RECT 1007.4200 2468.7600 1012.8800 2564.0200 ;
      RECT 2438.9200 2468.5000 2444.2800 2564.0200 ;
      RECT 2436.3200 2468.5000 2436.7200 2564.0200 ;
      RECT 2398.9000 2468.5000 2434.1200 2568.0200 ;
      RECT 2396.3000 2468.5000 2396.7000 2470.4600 ;
      RECT 2378.7800 2468.5000 2384.1400 2474.3000 ;
      RECT 2376.1800 2468.5000 2376.5800 2473.5200 ;
      RECT 2178.6800 2468.5000 2373.9800 2472.1000 ;
      RECT 2176.0800 2468.5000 2176.4800 2472.1000 ;
      RECT 2168.7200 2468.5000 2173.8800 2474.3000 ;
      RECT 1938.3400 2468.5000 1943.7000 2474.3000 ;
      RECT 1935.7400 2468.5000 1936.1400 2473.5200 ;
      RECT 1738.2400 2468.5000 1933.5400 2472.1000 ;
      RECT 1735.6400 2468.5000 1736.0400 2472.1000 ;
      RECT 1728.2800 2468.5000 1733.4400 2474.3000 ;
      RECT 1718.1200 2468.5000 1723.4800 2474.3000 ;
      RECT 1715.5200 2468.5000 1715.9200 2473.5200 ;
      RECT 1518.0200 2468.5000 1713.3200 2472.1000 ;
      RECT 1515.4200 2468.5000 1515.8200 2472.1000 ;
      RECT 1508.0600 2468.5000 1513.2200 2474.3000 ;
      RECT 1497.9000 2468.5000 1503.2600 2474.3000 ;
      RECT 1495.3000 2468.5000 1495.7000 2473.5200 ;
      RECT 1297.8000 2468.5000 1493.1000 2472.1000 ;
      RECT 1295.2000 2468.5000 1295.6000 2472.1000 ;
      RECT 1287.9800 2468.5000 1293.0000 2474.3000 ;
      RECT 2396.3000 2467.3600 2444.2800 2468.5000 ;
      RECT 2388.9400 2467.3600 2394.1000 2470.4600 ;
      RECT 1007.4200 2466.5500 1062.9600 2468.7600 ;
      RECT 1728.2800 2466.3900 1943.7000 2468.5000 ;
      RECT 1062.4600 2464.3500 1062.9600 2466.5500 ;
      RECT 1007.4200 2464.3500 1060.2600 2466.5500 ;
      RECT 1943.2000 2464.1900 1943.7000 2466.3900 ;
      RECT 1728.2800 2464.1900 1941.0000 2466.3900 ;
      RECT 2168.7200 2463.8250 2384.1400 2468.5000 ;
      RECT 1728.2800 2463.8250 1943.7000 2464.1900 ;
      RECT 1508.0600 2463.8250 1723.4800 2468.5000 ;
      RECT 1287.9800 2463.8250 1503.2600 2468.5000 ;
      RECT 2183.2400 2457.8400 2384.1400 2463.8250 ;
      RECT 2168.7200 2457.8400 2181.0400 2463.8250 ;
      RECT 1742.8000 2457.8400 1943.7000 2463.8250 ;
      RECT 1728.2800 2457.8400 1740.6000 2463.8250 ;
      RECT 1522.5800 2457.8400 1723.4800 2463.8250 ;
      RECT 1508.0600 2457.8400 1520.3800 2463.8250 ;
      RECT 1302.3600 2457.8400 1503.2600 2463.8250 ;
      RECT 1287.9800 2457.8400 1300.1600 2463.8250 ;
      RECT 1075.1200 2456.9400 1283.0400 2469.3000 ;
      RECT 1067.7600 2456.9400 1072.9200 2472.1000 ;
      RECT 1955.8600 2456.6800 2163.9200 2469.0400 ;
      RECT 1948.5000 2456.6800 1953.6600 2474.3000 ;
      RECT 1007.4200 2263.3400 1062.9600 2464.3500 ;
      RECT 2388.9400 2263.0800 2444.2800 2467.3600 ;
      RECT 1007.4200 2260.6200 1055.3000 2263.3400 ;
      RECT 2396.3000 2260.3600 2444.2800 2263.0800 ;
      RECT 2168.7200 2260.3600 2384.1400 2457.8400 ;
      RECT 1728.2800 2260.3600 1943.7000 2457.8400 ;
      RECT 1508.0600 2260.3600 1723.4800 2457.8400 ;
      RECT 1287.9800 2260.3600 1503.2600 2457.8400 ;
      RECT 2178.6800 2252.4550 2384.1400 2260.3600 ;
      RECT 2168.7200 2252.4550 2176.4800 2260.3600 ;
      RECT 1738.2400 2252.4550 1943.7000 2260.3600 ;
      RECT 1728.2800 2252.4550 1736.0400 2260.3600 ;
      RECT 1518.0200 2252.4550 1723.4800 2260.3600 ;
      RECT 1508.0600 2252.4550 1515.8200 2260.3600 ;
      RECT 1297.8000 2252.4550 1503.2600 2260.3600 ;
      RECT 1287.9800 2252.4550 1295.6000 2260.3600 ;
      RECT 1017.4800 2251.3200 1055.3000 2260.6200 ;
      RECT 1007.4200 2251.3200 1015.2800 2260.6200 ;
      RECT 2436.3200 2251.0600 2444.2800 2260.3600 ;
      RECT 2396.3000 2251.0600 2434.1200 2260.3600 ;
      RECT 2168.7200 2251.0600 2384.1400 2252.4550 ;
      RECT 1728.2800 2251.0600 1943.7000 2252.4550 ;
      RECT 1508.0600 2251.0600 1723.4800 2252.4550 ;
      RECT 1287.9800 2251.0600 1503.2600 2252.4550 ;
      RECT 1055.1000 2239.1200 1055.3000 2251.3200 ;
      RECT 1017.4800 2239.1200 1052.9000 2251.3200 ;
      RECT 1015.0800 2239.1200 1015.2800 2251.3200 ;
      RECT 1007.4200 2239.1200 1012.8800 2251.3200 ;
      RECT 2438.9200 2238.8600 2444.2800 2251.0600 ;
      RECT 2436.3200 2238.8600 2436.7200 2251.0600 ;
      RECT 2398.9000 2238.8600 2434.1200 2251.0600 ;
      RECT 2396.3000 2238.8600 2396.7000 2251.0600 ;
      RECT 2378.7800 2238.8600 2384.1400 2251.0600 ;
      RECT 2376.1800 2238.8600 2376.5800 2251.0600 ;
      RECT 2178.6800 2238.8600 2373.9800 2251.0600 ;
      RECT 2176.0800 2238.8600 2176.4800 2251.0600 ;
      RECT 1938.3400 2238.8600 1943.7000 2251.0600 ;
      RECT 1935.7400 2238.8600 1936.1400 2251.0600 ;
      RECT 1738.2400 2238.8600 1933.5400 2251.0600 ;
      RECT 1735.6400 2238.8600 1736.0400 2251.0600 ;
      RECT 1718.1200 2238.8600 1723.4800 2251.0600 ;
      RECT 1715.5200 2238.8600 1715.9200 2251.0600 ;
      RECT 1518.0200 2238.8600 1713.3200 2251.0600 ;
      RECT 1515.4200 2238.8600 1515.8200 2251.0600 ;
      RECT 1497.9000 2238.8600 1503.2600 2251.0600 ;
      RECT 1495.3000 2238.8600 1495.7000 2251.0600 ;
      RECT 1297.8000 2238.8600 1493.1000 2251.0600 ;
      RECT 1295.2000 2238.8600 1295.6000 2251.0600 ;
      RECT 1057.5000 2228.4600 1062.9600 2263.3400 ;
      RECT 1007.4200 2228.4600 1055.3000 2239.1200 ;
      RECT 2396.3000 2228.2000 2444.2800 2238.8600 ;
      RECT 2388.9400 2228.2000 2394.1000 2263.0800 ;
      RECT 2176.0800 2228.2000 2384.1400 2238.8600 ;
      RECT 2168.7200 2228.2000 2173.8800 2251.0600 ;
      RECT 1735.6400 2228.2000 1943.7000 2238.8600 ;
      RECT 1728.2800 2228.2000 1733.4400 2251.0600 ;
      RECT 1515.4200 2228.2000 1723.4800 2238.8600 ;
      RECT 1508.0600 2228.2000 1513.2200 2251.0600 ;
      RECT 1295.2000 2228.2000 1503.2600 2238.8600 ;
      RECT 1287.9800 2228.2000 1293.0000 2251.0600 ;
      RECT 1067.7600 2030.9800 1283.0400 2456.9400 ;
      RECT 1007.4200 2030.9800 1062.9600 2228.4600 ;
      RECT 2388.9400 2030.7200 2444.2800 2228.2000 ;
      RECT 2168.7200 2030.7200 2384.1400 2228.2000 ;
      RECT 1948.5000 2030.7200 2163.9200 2456.6800 ;
      RECT 1728.2800 2030.7200 1943.7000 2228.2000 ;
      RECT 1508.0600 2030.7200 1723.4800 2228.2000 ;
      RECT 1287.9800 2030.7200 1503.2600 2228.2000 ;
      RECT 9.3000 2025.9200 1002.6200 2564.0200 ;
      RECT 9.3000 2024.8400 1001.0300 2025.9200 ;
      RECT 1077.7200 2023.0750 1283.0400 2030.9800 ;
      RECT 1067.7600 2023.0750 1075.5200 2030.9800 ;
      RECT 2178.6800 2022.8150 2384.1400 2030.7200 ;
      RECT 2168.7200 2022.8150 2176.4800 2030.7200 ;
      RECT 1958.4600 2022.8150 2163.9200 2030.7200 ;
      RECT 1948.5000 2022.8150 1956.2600 2030.7200 ;
      RECT 1738.2400 2022.8150 1943.7000 2030.7200 ;
      RECT 1728.2800 2022.8150 1736.0400 2030.7200 ;
      RECT 1518.0200 2022.8150 1723.4800 2030.7200 ;
      RECT 1508.0600 2022.8150 1515.8200 2030.7200 ;
      RECT 1297.8000 2022.8150 1503.2600 2030.7200 ;
      RECT 1287.9800 2022.8150 1295.6000 2030.7200 ;
      RECT 1067.7600 2021.6800 1283.0400 2023.0750 ;
      RECT 1017.4800 2021.6800 1062.9600 2030.9800 ;
      RECT 1007.4200 2021.6800 1015.2800 2030.9800 ;
      RECT 2436.3200 2021.4200 2444.2800 2030.7200 ;
      RECT 2388.9400 2021.4200 2434.1200 2030.7200 ;
      RECT 2168.7200 2021.4200 2384.1400 2022.8150 ;
      RECT 1948.5000 2021.4200 2163.9200 2022.8150 ;
      RECT 1728.2800 2021.4200 1943.7000 2022.8150 ;
      RECT 1508.0600 2021.4200 1723.4800 2022.8150 ;
      RECT 1287.9800 2021.4200 1503.2600 2022.8150 ;
      RECT 9.3000 2017.8800 1002.6200 2024.8400 ;
      RECT 965.0200 2015.2800 1002.6200 2017.8800 ;
      RECT 9.3000 2015.2800 155.2200 2017.8800 ;
      RECT 1277.8200 2010.0200 1283.0400 2021.6800 ;
      RECT 1275.2200 2010.0200 1275.6200 2021.6800 ;
      RECT 1077.7200 2010.0200 1273.0200 2021.6800 ;
      RECT 1075.1200 2010.0200 1075.5200 2021.6800 ;
      RECT 2158.5600 2009.7600 2163.9200 2021.4200 ;
      RECT 2155.9600 2009.7600 2156.3600 2021.4200 ;
      RECT 1958.4600 2009.7600 2153.7600 2021.4200 ;
      RECT 1955.8600 2009.7600 1956.2600 2021.4200 ;
      RECT 1055.1000 2009.4800 1055.3000 2021.6800 ;
      RECT 1017.4800 2009.4800 1052.9000 2021.6800 ;
      RECT 1015.0800 2009.4800 1015.2800 2021.6800 ;
      RECT 1007.4200 2009.4800 1012.8800 2021.6800 ;
      RECT 2438.9200 2009.2200 2444.2800 2021.4200 ;
      RECT 2436.3200 2009.2200 2436.7200 2021.4200 ;
      RECT 2398.9000 2009.2200 2434.1200 2021.4200 ;
      RECT 2396.3000 2009.2200 2396.7000 2021.4200 ;
      RECT 2378.7800 2009.2200 2384.1400 2021.4200 ;
      RECT 2376.1800 2009.2200 2376.5800 2021.4200 ;
      RECT 2178.6800 2009.2200 2373.9800 2021.4200 ;
      RECT 2176.0800 2009.2200 2176.4800 2021.4200 ;
      RECT 1938.3400 2009.2200 1943.7000 2021.4200 ;
      RECT 1935.7400 2009.2200 1936.1400 2021.4200 ;
      RECT 1738.2400 2009.2200 1933.5400 2021.4200 ;
      RECT 1735.6400 2009.2200 1736.0400 2021.4200 ;
      RECT 1718.1200 2009.2200 1723.4800 2021.4200 ;
      RECT 1715.5200 2009.2200 1715.9200 2021.4200 ;
      RECT 1518.0200 2009.2200 1713.3200 2021.4200 ;
      RECT 1515.4200 2009.2200 1515.8200 2021.4200 ;
      RECT 1497.9000 2009.2200 1503.2600 2021.4200 ;
      RECT 1495.3000 2009.2200 1495.7000 2021.4200 ;
      RECT 1297.8000 2009.2200 1493.1000 2021.4200 ;
      RECT 1295.2000 2009.2200 1295.6000 2021.4200 ;
      RECT 1057.5000 2007.2700 1062.9600 2021.6800 ;
      RECT 1735.6400 2007.1100 1943.7000 2009.2200 ;
      RECT 1062.4600 2005.0700 1062.9600 2007.2700 ;
      RECT 1057.5000 2005.0700 1060.2600 2007.2700 ;
      RECT 1943.2000 2004.9100 1943.7000 2007.1100 ;
      RECT 1735.6400 2004.9100 1941.0000 2007.1100 ;
      RECT 1057.5000 1998.8200 1062.9600 2005.0700 ;
      RECT 1007.4200 1998.8200 1055.3000 2009.4800 ;
      RECT 2396.3000 1998.5600 2444.2800 2009.2200 ;
      RECT 2388.9400 1998.5600 2394.1000 2021.4200 ;
      RECT 2176.0800 1998.5600 2384.1400 2009.2200 ;
      RECT 2168.7200 1998.5600 2173.8800 2021.4200 ;
      RECT 1735.6400 1998.5600 1943.7000 2004.9100 ;
      RECT 1728.2800 1998.5600 1733.4400 2021.4200 ;
      RECT 1515.4200 1998.5600 1723.4800 2009.2200 ;
      RECT 1508.0600 1998.5600 1513.2200 2021.4200 ;
      RECT 1295.2000 1998.5600 1503.2600 2009.2200 ;
      RECT 1287.9800 1998.5600 1293.0000 2021.4200 ;
      RECT 1075.1200 1997.6600 1283.0400 2010.0200 ;
      RECT 1067.7600 1997.6600 1072.9200 2021.6800 ;
      RECT 1955.8600 1997.4000 2163.9200 2009.7600 ;
      RECT 1948.5000 1997.4000 1953.6600 2021.4200 ;
      RECT 2497.4200 1932.8000 3302.8200 2568.0200 ;
      RECT 157.4200 1932.8000 962.8200 2017.8800 ;
      RECT 3289.7800 1930.6000 3302.8200 1932.8000 ;
      RECT 2497.4200 1930.6000 3287.5800 1932.8000 ;
      RECT 949.7800 1930.6000 962.8200 1932.8000 ;
      RECT 157.4200 1930.6000 947.5800 1932.8000 ;
      RECT 2497.4200 1907.8000 3302.8200 1930.6000 ;
      RECT 157.4200 1907.8000 962.8200 1930.6000 ;
      RECT 3289.7800 1905.6000 3302.8200 1907.8000 ;
      RECT 2497.4200 1905.6000 3287.5800 1907.8000 ;
      RECT 949.7800 1905.6000 962.8200 1907.8000 ;
      RECT 157.4200 1905.6000 947.5800 1907.8000 ;
      RECT 1007.4200 1801.3400 1062.9600 1998.8200 ;
      RECT 2388.9400 1801.0800 2444.2800 1998.5600 ;
      RECT 2168.7200 1801.0800 2384.1400 1998.5600 ;
      RECT 1728.2800 1801.0800 1943.7000 1998.5600 ;
      RECT 1508.0600 1801.0800 1723.4800 1998.5600 ;
      RECT 1287.9800 1801.0800 1503.2600 1998.5600 ;
      RECT 2178.6800 1793.1750 2384.1400 1801.0800 ;
      RECT 2168.7200 1793.1750 2176.4800 1801.0800 ;
      RECT 1738.2400 1793.1750 1943.7000 1801.0800 ;
      RECT 1728.2800 1793.1750 1736.0400 1801.0800 ;
      RECT 1518.0200 1793.1750 1723.4800 1801.0800 ;
      RECT 1508.0600 1793.1750 1515.8200 1801.0800 ;
      RECT 1297.8000 1793.1750 1503.2600 1801.0800 ;
      RECT 1287.9800 1793.1750 1295.6000 1801.0800 ;
      RECT 1017.4800 1792.0400 1062.9600 1801.3400 ;
      RECT 1007.4200 1792.0400 1015.2800 1801.3400 ;
      RECT 2436.3200 1791.7800 2444.2800 1801.0800 ;
      RECT 2388.9400 1791.7800 2434.1200 1801.0800 ;
      RECT 2168.7200 1791.7800 2384.1400 1793.1750 ;
      RECT 1728.2800 1791.7800 1943.7000 1793.1750 ;
      RECT 1508.0600 1791.7800 1723.4800 1793.1750 ;
      RECT 1287.9800 1791.7800 1503.2600 1793.1750 ;
      RECT 1057.5000 1779.8400 1062.9600 1792.0400 ;
      RECT 1055.1000 1779.8400 1055.3000 1792.0400 ;
      RECT 1017.4800 1779.8400 1052.9000 1792.0400 ;
      RECT 1015.0800 1779.8400 1015.2800 1792.0400 ;
      RECT 2438.9200 1779.5800 2444.2800 1791.7800 ;
      RECT 2436.3200 1779.5800 2436.7200 1791.7800 ;
      RECT 2398.9000 1779.5800 2434.1200 1791.7800 ;
      RECT 2396.3000 1779.5800 2396.7000 1791.7800 ;
      RECT 2378.7800 1779.5800 2384.1400 1791.7800 ;
      RECT 2376.1800 1779.5800 2376.5800 1791.7800 ;
      RECT 2178.6800 1779.5800 2373.9800 1791.7800 ;
      RECT 2176.0800 1779.5800 2176.4800 1791.7800 ;
      RECT 1938.3400 1779.5800 1943.7000 1791.7800 ;
      RECT 1935.7400 1779.5800 1936.1400 1791.7800 ;
      RECT 1738.2400 1779.5800 1933.5400 1791.7800 ;
      RECT 1735.6400 1779.5800 1736.0400 1791.7800 ;
      RECT 1718.1200 1779.5800 1723.4800 1791.7800 ;
      RECT 1715.5200 1779.5800 1715.9200 1791.7800 ;
      RECT 1518.0200 1779.5800 1713.3200 1791.7800 ;
      RECT 1515.4200 1779.5800 1515.8200 1791.7800 ;
      RECT 1497.9000 1779.5800 1503.2600 1791.7800 ;
      RECT 1495.3000 1779.5800 1495.7000 1791.7800 ;
      RECT 1297.8000 1779.5800 1493.1000 1791.7800 ;
      RECT 1295.2000 1779.5800 1295.6000 1791.7800 ;
      RECT 1015.0800 1769.1800 1062.9600 1779.8400 ;
      RECT 1007.4200 1769.1800 1012.8800 1792.0400 ;
      RECT 2396.3000 1768.9200 2444.2800 1779.5800 ;
      RECT 2388.9400 1768.9200 2394.1000 1791.7800 ;
      RECT 2176.0800 1768.9200 2384.1400 1779.5800 ;
      RECT 2168.7200 1768.9200 2173.8800 1791.7800 ;
      RECT 1735.6400 1768.9200 1943.7000 1779.5800 ;
      RECT 1728.2800 1768.9200 1733.4400 1791.7800 ;
      RECT 1515.4200 1768.9200 1723.4800 1779.5800 ;
      RECT 1508.0600 1768.9200 1513.2200 1791.7800 ;
      RECT 1295.2000 1768.9200 1503.2600 1779.5800 ;
      RECT 1287.9800 1768.9200 1293.0000 1791.7800 ;
      RECT 1067.7600 1571.7000 1283.0400 1997.6600 ;
      RECT 1007.4200 1571.7000 1062.9600 1769.1800 ;
      RECT 2388.9400 1571.4400 2444.2800 1768.9200 ;
      RECT 2168.7200 1571.4400 2384.1400 1768.9200 ;
      RECT 1948.5000 1571.4400 2163.9200 1997.4000 ;
      RECT 1728.2800 1571.4400 1943.7000 1768.9200 ;
      RECT 1508.0600 1571.4400 1723.4800 1768.9200 ;
      RECT 1287.9800 1571.4400 1503.2600 1768.9200 ;
      RECT 1077.7200 1563.7950 1283.0400 1571.7000 ;
      RECT 1067.7600 1563.7950 1075.5200 1571.7000 ;
      RECT 2178.6800 1563.5350 2384.1400 1571.4400 ;
      RECT 2168.7200 1563.5350 2176.4800 1571.4400 ;
      RECT 1958.4600 1563.5350 2163.9200 1571.4400 ;
      RECT 1948.5000 1563.5350 1956.2600 1571.4400 ;
      RECT 1738.2400 1563.5350 1943.7000 1571.4400 ;
      RECT 1728.2800 1563.5350 1736.0400 1571.4400 ;
      RECT 1518.0200 1563.5350 1723.4800 1571.4400 ;
      RECT 1508.0600 1563.5350 1515.8200 1571.4400 ;
      RECT 1297.8000 1563.5350 1503.2600 1571.4400 ;
      RECT 1287.9800 1563.5350 1295.6000 1571.4400 ;
      RECT 1067.7600 1562.4000 1283.0400 1563.7950 ;
      RECT 1017.4800 1562.4000 1062.9600 1571.7000 ;
      RECT 1007.4200 1562.4000 1015.2800 1571.7000 ;
      RECT 2436.3200 1562.1400 2444.2800 1571.4400 ;
      RECT 2388.9400 1562.1400 2434.1200 1571.4400 ;
      RECT 2168.7200 1562.1400 2384.1400 1563.5350 ;
      RECT 1948.5000 1562.1400 2163.9200 1563.5350 ;
      RECT 1728.2800 1562.1400 1943.7000 1563.5350 ;
      RECT 1508.0600 1562.1400 1723.4800 1563.5350 ;
      RECT 1287.9800 1562.1400 1503.2600 1563.5350 ;
      RECT 1277.8200 1550.7400 1283.0400 1562.4000 ;
      RECT 1275.2200 1550.7400 1275.6200 1562.4000 ;
      RECT 1077.7200 1550.7400 1273.0200 1562.4000 ;
      RECT 1075.1200 1550.7400 1075.5200 1562.4000 ;
      RECT 2158.5600 1550.4800 2163.9200 1562.1400 ;
      RECT 2155.9600 1550.4800 2156.3600 1562.1400 ;
      RECT 1958.4600 1550.4800 2153.7600 1562.1400 ;
      RECT 1955.8600 1550.4800 1956.2600 1562.1400 ;
      RECT 1055.1000 1550.2000 1055.3000 1562.4000 ;
      RECT 1017.4800 1550.2000 1052.9000 1562.4000 ;
      RECT 1015.0800 1550.2000 1015.2800 1562.4000 ;
      RECT 1007.4200 1550.2000 1012.8800 1562.4000 ;
      RECT 2438.9200 1549.9400 2444.2800 1562.1400 ;
      RECT 2436.3200 1549.9400 2436.7200 1562.1400 ;
      RECT 2398.9000 1549.9400 2434.1200 1562.1400 ;
      RECT 2396.3000 1549.9400 2396.7000 1562.1400 ;
      RECT 2378.7800 1549.9400 2384.1400 1562.1400 ;
      RECT 2376.1800 1549.9400 2376.5800 1562.1400 ;
      RECT 2178.6800 1549.9400 2373.9800 1562.1400 ;
      RECT 2176.0800 1549.9400 2176.4800 1562.1400 ;
      RECT 1938.3400 1549.9400 1943.7000 1562.1400 ;
      RECT 1935.7400 1549.9400 1936.1400 1562.1400 ;
      RECT 1738.2400 1549.9400 1933.5400 1562.1400 ;
      RECT 1735.6400 1549.9400 1736.0400 1562.1400 ;
      RECT 1718.1200 1549.9400 1723.4800 1562.1400 ;
      RECT 1715.5200 1549.9400 1715.9200 1562.1400 ;
      RECT 1518.0200 1549.9400 1713.3200 1562.1400 ;
      RECT 1515.4200 1549.9400 1515.8200 1562.1400 ;
      RECT 1497.9000 1549.9400 1503.2600 1562.1400 ;
      RECT 1495.3000 1549.9400 1495.7000 1562.1400 ;
      RECT 1297.8000 1549.9400 1493.1000 1562.1400 ;
      RECT 1295.2000 1549.9400 1295.6000 1562.1400 ;
      RECT 1057.5000 1547.9900 1062.9600 1562.4000 ;
      RECT 1735.6400 1547.8300 1943.7000 1549.9400 ;
      RECT 1062.4600 1545.7900 1062.9600 1547.9900 ;
      RECT 1057.5000 1545.7900 1060.2600 1547.9900 ;
      RECT 1943.2000 1545.6300 1943.7000 1547.8300 ;
      RECT 1735.6400 1545.6300 1941.0000 1547.8300 ;
      RECT 1057.5000 1539.5400 1062.9600 1545.7900 ;
      RECT 1007.4200 1539.5400 1055.3000 1550.2000 ;
      RECT 2396.3000 1539.2800 2444.2800 1549.9400 ;
      RECT 2388.9400 1539.2800 2394.1000 1562.1400 ;
      RECT 2176.0800 1539.2800 2384.1400 1549.9400 ;
      RECT 2168.7200 1539.2800 2173.8800 1562.1400 ;
      RECT 1735.6400 1539.2800 1943.7000 1545.6300 ;
      RECT 1728.2800 1539.2800 1733.4400 1562.1400 ;
      RECT 1515.4200 1539.2800 1723.4800 1549.9400 ;
      RECT 1508.0600 1539.2800 1513.2200 1562.1400 ;
      RECT 1295.2000 1539.2800 1503.2600 1549.9400 ;
      RECT 1287.9800 1539.2800 1293.0000 1562.1400 ;
      RECT 1075.1200 1538.3800 1283.0400 1550.7400 ;
      RECT 1067.7600 1538.3800 1072.9200 1562.4000 ;
      RECT 1955.8600 1538.1200 2163.9200 1550.4800 ;
      RECT 1948.5000 1538.1200 1953.6600 1562.1400 ;
      RECT 1007.4200 1342.0600 1062.9600 1539.5400 ;
      RECT 2388.9400 1341.8000 2444.2800 1539.2800 ;
      RECT 2168.7200 1341.8000 2384.1400 1539.2800 ;
      RECT 1728.2800 1341.8000 1943.7000 1539.2800 ;
      RECT 1508.0600 1341.8000 1723.4800 1539.2800 ;
      RECT 1287.9800 1341.8000 1503.2600 1539.2800 ;
      RECT 2178.6800 1333.8950 2384.1400 1341.8000 ;
      RECT 2168.7200 1333.8950 2176.4800 1341.8000 ;
      RECT 1738.2400 1333.8950 1943.7000 1341.8000 ;
      RECT 1728.2800 1333.8950 1736.0400 1341.8000 ;
      RECT 1518.0200 1333.8950 1723.4800 1341.8000 ;
      RECT 1508.0600 1333.8950 1515.8200 1341.8000 ;
      RECT 1297.8000 1333.8950 1503.2600 1341.8000 ;
      RECT 1287.9800 1333.8950 1295.6000 1341.8000 ;
      RECT 1017.4800 1332.7600 1062.9600 1342.0600 ;
      RECT 1007.4200 1332.7600 1015.2800 1342.0600 ;
      RECT 2436.3200 1332.5000 2444.2800 1341.8000 ;
      RECT 2388.9400 1332.5000 2434.1200 1341.8000 ;
      RECT 2168.7200 1332.5000 2384.1400 1333.8950 ;
      RECT 1728.2800 1332.5000 1943.7000 1333.8950 ;
      RECT 1508.0600 1332.5000 1723.4800 1333.8950 ;
      RECT 1287.9800 1332.5000 1503.2600 1333.8950 ;
      RECT 1057.5000 1320.5600 1062.9600 1332.7600 ;
      RECT 1055.1000 1320.5600 1055.3000 1332.7600 ;
      RECT 1017.4800 1320.5600 1052.9000 1332.7600 ;
      RECT 1015.0800 1320.5600 1015.2800 1332.7600 ;
      RECT 2438.9200 1320.3000 2444.2800 1332.5000 ;
      RECT 2436.3200 1320.3000 2436.7200 1332.5000 ;
      RECT 2398.9000 1320.3000 2434.1200 1332.5000 ;
      RECT 2396.3000 1320.3000 2396.7000 1332.5000 ;
      RECT 2378.7800 1320.3000 2384.1400 1332.5000 ;
      RECT 2376.1800 1320.3000 2376.5800 1332.5000 ;
      RECT 2178.6800 1320.3000 2373.9800 1332.5000 ;
      RECT 2176.0800 1320.3000 2176.4800 1332.5000 ;
      RECT 1938.3400 1320.3000 1943.7000 1332.5000 ;
      RECT 1935.7400 1320.3000 1936.1400 1332.5000 ;
      RECT 1738.2400 1320.3000 1933.5400 1332.5000 ;
      RECT 1735.6400 1320.3000 1736.0400 1332.5000 ;
      RECT 1718.1200 1320.3000 1723.4800 1332.5000 ;
      RECT 1715.5200 1320.3000 1715.9200 1332.5000 ;
      RECT 1518.0200 1320.3000 1713.3200 1332.5000 ;
      RECT 1515.4200 1320.3000 1515.8200 1332.5000 ;
      RECT 1497.9000 1320.3000 1503.2600 1332.5000 ;
      RECT 1495.3000 1320.3000 1495.7000 1332.5000 ;
      RECT 1297.8000 1320.3000 1493.1000 1332.5000 ;
      RECT 1295.2000 1320.3000 1295.6000 1332.5000 ;
      RECT 1015.0800 1309.9000 1062.9600 1320.5600 ;
      RECT 1007.4200 1309.9000 1012.8800 1332.7600 ;
      RECT 2396.3000 1309.6400 2444.2800 1320.3000 ;
      RECT 2388.9400 1309.6400 2394.1000 1332.5000 ;
      RECT 2176.0800 1309.6400 2384.1400 1320.3000 ;
      RECT 2168.7200 1309.6400 2173.8800 1332.5000 ;
      RECT 1735.6400 1309.6400 1943.7000 1320.3000 ;
      RECT 1728.2800 1309.6400 1733.4400 1332.5000 ;
      RECT 1515.4200 1309.6400 1723.4800 1320.3000 ;
      RECT 1508.0600 1309.6400 1513.2200 1332.5000 ;
      RECT 1295.2000 1309.6400 1503.2600 1320.3000 ;
      RECT 1287.9800 1309.6400 1293.0000 1332.5000 ;
      RECT 1067.7600 1112.4200 1283.0400 1538.3800 ;
      RECT 1007.4200 1112.4200 1062.9600 1309.9000 ;
      RECT 2388.9400 1112.1600 2444.2800 1309.6400 ;
      RECT 2168.7200 1112.1600 2384.1400 1309.6400 ;
      RECT 1948.5000 1112.1600 2163.9200 1538.1200 ;
      RECT 1728.2800 1112.1600 1943.7000 1309.6400 ;
      RECT 1508.0600 1112.1600 1723.4800 1309.6400 ;
      RECT 1287.9800 1112.1600 1503.2600 1309.6400 ;
      RECT 1077.7200 1104.5150 1283.0400 1112.4200 ;
      RECT 1067.7600 1104.5150 1075.5200 1112.4200 ;
      RECT 2178.6800 1104.2550 2384.1400 1112.1600 ;
      RECT 2168.7200 1104.2550 2176.4800 1112.1600 ;
      RECT 1958.4600 1104.2550 2163.9200 1112.1600 ;
      RECT 1948.5000 1104.2550 1956.2600 1112.1600 ;
      RECT 1738.2400 1104.2550 1943.7000 1112.1600 ;
      RECT 1728.2800 1104.2550 1736.0400 1112.1600 ;
      RECT 1518.0200 1104.2550 1723.4800 1112.1600 ;
      RECT 1508.0600 1104.2550 1515.8200 1112.1600 ;
      RECT 1297.8000 1104.2550 1503.2600 1112.1600 ;
      RECT 1287.9800 1104.2550 1295.6000 1112.1600 ;
      RECT 1067.7600 1103.1200 1283.0400 1104.5150 ;
      RECT 1017.4800 1103.1200 1062.9600 1112.4200 ;
      RECT 1007.4200 1103.1200 1015.2800 1112.4200 ;
      RECT 2436.3200 1102.8600 2444.2800 1112.1600 ;
      RECT 2388.9400 1102.8600 2434.1200 1112.1600 ;
      RECT 2168.7200 1102.8600 2384.1400 1104.2550 ;
      RECT 1948.5000 1102.8600 2163.9200 1104.2550 ;
      RECT 1728.2800 1102.8600 1943.7000 1104.2550 ;
      RECT 1508.0600 1102.8600 1723.4800 1104.2550 ;
      RECT 1287.9800 1102.8600 1503.2600 1104.2550 ;
      RECT 1277.8200 1091.4600 1283.0400 1103.1200 ;
      RECT 1275.2200 1091.4600 1275.6200 1103.1200 ;
      RECT 1077.7200 1091.4600 1273.0200 1103.1200 ;
      RECT 1075.1200 1091.4600 1075.5200 1103.1200 ;
      RECT 2158.5600 1091.2000 2163.9200 1102.8600 ;
      RECT 2155.9600 1091.2000 2156.3600 1102.8600 ;
      RECT 1958.4600 1091.2000 2153.7600 1102.8600 ;
      RECT 1955.8600 1091.2000 1956.2600 1102.8600 ;
      RECT 1055.1000 1090.9200 1055.3000 1103.1200 ;
      RECT 1017.4800 1090.9200 1052.9000 1103.1200 ;
      RECT 1015.0800 1090.9200 1015.2800 1103.1200 ;
      RECT 1007.4200 1090.9200 1012.8800 1103.1200 ;
      RECT 2438.9200 1090.6600 2444.2800 1102.8600 ;
      RECT 2436.3200 1090.6600 2436.7200 1102.8600 ;
      RECT 2398.9000 1090.6600 2434.1200 1102.8600 ;
      RECT 2396.3000 1090.6600 2396.7000 1102.8600 ;
      RECT 2378.7800 1090.6600 2384.1400 1102.8600 ;
      RECT 2376.1800 1090.6600 2376.5800 1102.8600 ;
      RECT 2178.6800 1090.6600 2373.9800 1102.8600 ;
      RECT 2176.0800 1090.6600 2176.4800 1102.8600 ;
      RECT 1938.3400 1090.6600 1943.7000 1102.8600 ;
      RECT 1935.7400 1090.6600 1936.1400 1102.8600 ;
      RECT 1738.2400 1090.6600 1933.5400 1102.8600 ;
      RECT 1735.6400 1090.6600 1736.0400 1102.8600 ;
      RECT 1718.1200 1090.6600 1723.4800 1102.8600 ;
      RECT 1715.5200 1090.6600 1715.9200 1102.8600 ;
      RECT 1518.0200 1090.6600 1713.3200 1102.8600 ;
      RECT 1515.4200 1090.6600 1515.8200 1102.8600 ;
      RECT 1497.9000 1090.6600 1503.2600 1102.8600 ;
      RECT 1495.3000 1090.6600 1495.7000 1102.8600 ;
      RECT 1297.8000 1090.6600 1493.1000 1102.8600 ;
      RECT 1295.2000 1090.6600 1295.6000 1102.8600 ;
      RECT 1057.5000 1088.7100 1062.9600 1103.1200 ;
      RECT 1735.6400 1088.5500 1943.7000 1090.6600 ;
      RECT 1062.4600 1086.5100 1062.9600 1088.7100 ;
      RECT 1057.5000 1086.5100 1060.2600 1088.7100 ;
      RECT 1943.2000 1086.3500 1943.7000 1088.5500 ;
      RECT 1735.6400 1086.3500 1941.0000 1088.5500 ;
      RECT 1057.5000 1080.2600 1062.9600 1086.5100 ;
      RECT 1007.4200 1080.2600 1055.3000 1090.9200 ;
      RECT 2396.3000 1080.0000 2444.2800 1090.6600 ;
      RECT 2388.9400 1080.0000 2394.1000 1102.8600 ;
      RECT 2176.0800 1080.0000 2384.1400 1090.6600 ;
      RECT 2168.7200 1080.0000 2173.8800 1102.8600 ;
      RECT 1735.6400 1080.0000 1943.7000 1086.3500 ;
      RECT 1728.2800 1080.0000 1733.4400 1102.8600 ;
      RECT 1515.4200 1080.0000 1723.4800 1090.6600 ;
      RECT 1508.0600 1080.0000 1513.2200 1102.8600 ;
      RECT 1295.2000 1080.0000 1503.2600 1090.6600 ;
      RECT 1287.9800 1080.0000 1293.0000 1102.8600 ;
      RECT 1075.1200 1079.1000 1283.0400 1091.4600 ;
      RECT 1067.7600 1079.1000 1072.9200 1103.1200 ;
      RECT 1955.8600 1078.8400 2163.9200 1091.2000 ;
      RECT 1948.5000 1078.8400 1953.6600 1102.8600 ;
      RECT 1007.4200 882.7800 1062.9600 1080.2600 ;
      RECT 2388.9400 882.5200 2444.2800 1080.0000 ;
      RECT 2168.7200 882.5200 2384.1400 1080.0000 ;
      RECT 1728.2800 882.5200 1943.7000 1080.0000 ;
      RECT 1508.0600 882.5200 1723.4800 1080.0000 ;
      RECT 1287.9800 882.5200 1503.2600 1080.0000 ;
      RECT 2178.6800 874.6150 2384.1400 882.5200 ;
      RECT 2168.7200 874.6150 2176.4800 882.5200 ;
      RECT 1738.2400 874.6150 1943.7000 882.5200 ;
      RECT 1728.2800 874.6150 1736.0400 882.5200 ;
      RECT 1518.0200 874.6150 1723.4800 882.5200 ;
      RECT 1508.0600 874.6150 1515.8200 882.5200 ;
      RECT 1297.8000 874.6150 1503.2600 882.5200 ;
      RECT 1287.9800 874.6150 1295.6000 882.5200 ;
      RECT 1017.4800 873.4800 1062.9600 882.7800 ;
      RECT 1007.4200 873.4800 1015.2800 882.7800 ;
      RECT 2436.3200 873.2200 2444.2800 882.5200 ;
      RECT 2388.9400 873.2200 2434.1200 882.5200 ;
      RECT 2168.7200 873.2200 2384.1400 874.6150 ;
      RECT 1728.2800 873.2200 1943.7000 874.6150 ;
      RECT 1508.0600 873.2200 1723.4800 874.6150 ;
      RECT 1287.9800 873.2200 1503.2600 874.6150 ;
      RECT 1057.5000 861.2800 1062.9600 873.4800 ;
      RECT 1055.1000 861.2800 1055.3000 873.4800 ;
      RECT 1017.4800 861.2800 1052.9000 873.4800 ;
      RECT 1015.0800 861.2800 1015.2800 873.4800 ;
      RECT 2438.9200 861.0200 2444.2800 873.2200 ;
      RECT 2436.3200 861.0200 2436.7200 873.2200 ;
      RECT 2398.9000 861.0200 2434.1200 873.2200 ;
      RECT 2396.3000 861.0200 2396.7000 873.2200 ;
      RECT 2378.7800 861.0200 2384.1400 873.2200 ;
      RECT 2376.1800 861.0200 2376.5800 873.2200 ;
      RECT 2178.6800 861.0200 2373.9800 873.2200 ;
      RECT 2176.0800 861.0200 2176.4800 873.2200 ;
      RECT 1938.3400 861.0200 1943.7000 873.2200 ;
      RECT 1935.7400 861.0200 1936.1400 873.2200 ;
      RECT 1738.2400 861.0200 1933.5400 873.2200 ;
      RECT 1735.6400 861.0200 1736.0400 873.2200 ;
      RECT 1718.1200 861.0200 1723.4800 873.2200 ;
      RECT 1715.5200 861.0200 1715.9200 873.2200 ;
      RECT 1518.0200 861.0200 1713.3200 873.2200 ;
      RECT 1515.4200 861.0200 1515.8200 873.2200 ;
      RECT 1497.9000 861.0200 1503.2600 873.2200 ;
      RECT 1495.3000 861.0200 1495.7000 873.2200 ;
      RECT 1297.8000 861.0200 1493.1000 873.2200 ;
      RECT 1295.2000 861.0200 1295.6000 873.2200 ;
      RECT 1015.0800 850.6200 1062.9600 861.2800 ;
      RECT 1007.4200 850.6200 1012.8800 873.4800 ;
      RECT 2396.3000 850.3600 2444.2800 861.0200 ;
      RECT 2388.9400 850.3600 2394.1000 873.2200 ;
      RECT 2176.0800 850.3600 2384.1400 861.0200 ;
      RECT 2168.7200 850.3600 2173.8800 873.2200 ;
      RECT 1735.6400 850.3600 1943.7000 861.0200 ;
      RECT 1728.2800 850.3600 1733.4400 873.2200 ;
      RECT 1515.4200 850.3600 1723.4800 861.0200 ;
      RECT 1508.0600 850.3600 1513.2200 873.2200 ;
      RECT 1295.2000 850.3600 1503.2600 861.0200 ;
      RECT 1287.9800 850.3600 1293.0000 873.2200 ;
      RECT 1067.7600 653.1400 1283.0400 1079.1000 ;
      RECT 1007.4200 653.1400 1062.9600 850.6200 ;
      RECT 2388.9400 652.8800 2444.2800 850.3600 ;
      RECT 2168.7200 652.8800 2384.1400 850.3600 ;
      RECT 1948.5000 652.8800 2163.9200 1078.8400 ;
      RECT 1728.2800 652.8800 1943.7000 850.3600 ;
      RECT 1508.0600 652.8800 1723.4800 850.3600 ;
      RECT 1287.9800 652.8800 1503.2600 850.3600 ;
      RECT 1077.7200 645.2350 1283.0400 653.1400 ;
      RECT 1067.7600 645.2350 1075.5200 653.1400 ;
      RECT 2178.6800 644.9750 2384.1400 652.8800 ;
      RECT 2168.7200 644.9750 2176.4800 652.8800 ;
      RECT 1958.4600 644.9750 2163.9200 652.8800 ;
      RECT 1948.5000 644.9750 1956.2600 652.8800 ;
      RECT 1738.2400 644.9750 1943.7000 652.8800 ;
      RECT 1728.2800 644.9750 1736.0400 652.8800 ;
      RECT 1518.0200 644.9750 1723.4800 652.8800 ;
      RECT 1508.0600 644.9750 1515.8200 652.8800 ;
      RECT 1297.8000 644.9750 1503.2600 652.8800 ;
      RECT 1287.9800 644.9750 1295.6000 652.8800 ;
      RECT 1067.7600 643.8400 1283.0400 645.2350 ;
      RECT 1017.4800 643.8400 1062.9600 653.1400 ;
      RECT 1007.4200 643.8400 1015.2800 653.1400 ;
      RECT 2436.3200 643.5800 2444.2800 652.8800 ;
      RECT 2388.9400 643.5800 2434.1200 652.8800 ;
      RECT 2168.7200 643.5800 2384.1400 644.9750 ;
      RECT 1948.5000 643.5800 2163.9200 644.9750 ;
      RECT 1728.2800 643.5800 1943.7000 644.9750 ;
      RECT 1508.0600 643.5800 1723.4800 644.9750 ;
      RECT 1287.9800 643.5800 1503.2600 644.9750 ;
      RECT 157.4200 640.0400 962.8200 1905.6000 ;
      RECT 965.0200 637.8400 965.4200 2015.2800 ;
      RECT 665.0200 637.8400 962.8200 640.0400 ;
      RECT 157.4200 637.8400 505.2200 640.0400 ;
      RECT 154.8200 637.8400 155.2200 2015.2800 ;
      RECT 665.0200 637.4400 965.4200 637.8400 ;
      RECT 154.8200 637.4400 505.2200 637.8400 ;
      RECT 967.6200 635.2400 1002.6200 2015.2800 ;
      RECT 667.6200 635.2400 965.4200 637.4400 ;
      RECT 154.8200 635.2400 502.6200 637.4400 ;
      RECT 9.3000 635.2400 152.6200 2015.2800 ;
      RECT 1277.8200 632.1800 1283.0400 643.8400 ;
      RECT 1275.2200 632.1800 1275.6200 643.8400 ;
      RECT 1077.7200 632.1800 1273.0200 643.8400 ;
      RECT 1075.1200 632.1800 1075.5200 643.8400 ;
      RECT 2158.5600 631.9200 2163.9200 643.5800 ;
      RECT 2155.9600 631.9200 2156.3600 643.5800 ;
      RECT 1958.4600 631.9200 2153.7600 643.5800 ;
      RECT 1955.8600 631.9200 1956.2600 643.5800 ;
      RECT 1055.1000 631.6400 1055.3000 643.8400 ;
      RECT 1017.4800 631.6400 1052.9000 643.8400 ;
      RECT 1015.0800 631.6400 1015.2800 643.8400 ;
      RECT 1007.4200 631.6400 1012.8800 643.8400 ;
      RECT 2438.9200 631.3800 2444.2800 643.5800 ;
      RECT 2436.3200 631.3800 2436.7200 643.5800 ;
      RECT 2398.9000 631.3800 2434.1200 643.5800 ;
      RECT 2396.3000 631.3800 2396.7000 643.5800 ;
      RECT 2378.7800 631.3800 2384.1400 643.5800 ;
      RECT 2376.1800 631.3800 2376.5800 643.5800 ;
      RECT 2178.6800 631.3800 2373.9800 643.5800 ;
      RECT 2176.0800 631.3800 2176.4800 643.5800 ;
      RECT 1938.3400 631.3800 1943.7000 643.5800 ;
      RECT 1935.7400 631.3800 1936.1400 643.5800 ;
      RECT 1738.2400 631.3800 1933.5400 643.5800 ;
      RECT 1735.6400 631.3800 1736.0400 643.5800 ;
      RECT 1718.1200 631.3800 1723.4800 643.5800 ;
      RECT 1715.5200 631.3800 1715.9200 643.5800 ;
      RECT 1518.0200 631.3800 1713.3200 643.5800 ;
      RECT 1515.4200 631.3800 1515.8200 643.5800 ;
      RECT 1497.9000 631.3800 1503.2600 643.5800 ;
      RECT 1495.3000 631.3800 1495.7000 643.5800 ;
      RECT 1297.8000 631.3800 1493.1000 643.5800 ;
      RECT 1295.2000 631.3800 1295.6000 643.5800 ;
      RECT 1057.5000 629.4300 1062.9600 643.8400 ;
      RECT 1735.6400 629.2700 1943.7000 631.3800 ;
      RECT 1062.4600 627.2300 1062.9600 629.4300 ;
      RECT 1057.5000 627.2300 1060.2600 629.4300 ;
      RECT 1943.2000 627.0700 1943.7000 629.2700 ;
      RECT 1735.6400 627.0700 1941.0000 629.2700 ;
      RECT 1057.5000 620.9800 1062.9600 627.2300 ;
      RECT 1007.4200 620.9800 1055.3000 631.6400 ;
      RECT 2396.3000 620.7200 2444.2800 631.3800 ;
      RECT 2388.9400 620.7200 2394.1000 643.5800 ;
      RECT 2176.0800 620.7200 2384.1400 631.3800 ;
      RECT 2168.7200 620.7200 2173.8800 643.5800 ;
      RECT 1735.6400 620.7200 1943.7000 627.0700 ;
      RECT 1728.2800 620.7200 1733.4400 643.5800 ;
      RECT 1515.4200 620.7200 1723.4800 631.3800 ;
      RECT 1508.0600 620.7200 1513.2200 643.5800 ;
      RECT 1295.2000 620.7200 1503.2600 631.3800 ;
      RECT 1287.9800 620.7200 1293.0000 643.5800 ;
      RECT 1075.1200 619.8200 1283.0400 632.1800 ;
      RECT 1067.7600 619.8200 1072.9200 643.8400 ;
      RECT 1955.8600 619.5600 2163.9200 631.9200 ;
      RECT 1948.5000 619.5600 1953.6600 643.5800 ;
      RECT 507.4200 507.2800 662.8200 640.0400 ;
      RECT 649.7800 505.0800 662.8200 507.2800 ;
      RECT 507.4200 505.0800 647.5800 507.2800 ;
      RECT 507.4200 459.1200 662.8200 505.0800 ;
      RECT 649.7800 456.9200 662.8200 459.1200 ;
      RECT 507.4200 456.9200 647.5800 459.1200 ;
      RECT 1007.4200 423.5000 1062.9600 620.9800 ;
      RECT 2388.9400 423.2400 2444.2800 620.7200 ;
      RECT 2168.7200 423.2400 2384.1400 620.7200 ;
      RECT 1728.2800 423.2400 1943.7000 620.7200 ;
      RECT 1508.0600 423.2400 1723.4800 620.7200 ;
      RECT 1287.9800 423.2400 1503.2600 620.7200 ;
      RECT 2449.0800 415.6800 2492.6200 2564.0200 ;
      RECT 2178.6800 415.3350 2384.1400 423.2400 ;
      RECT 2168.7200 415.3350 2176.4800 423.2400 ;
      RECT 1738.2400 415.3350 1943.7000 423.2400 ;
      RECT 1728.2800 415.3350 1736.0400 423.2400 ;
      RECT 1518.0200 415.3350 1723.4800 423.2400 ;
      RECT 1508.0600 415.3350 1515.8200 423.2400 ;
      RECT 1297.8000 415.3350 1503.2600 423.2400 ;
      RECT 1287.9800 415.3350 1295.6000 423.2400 ;
      RECT 2450.4400 414.6000 2492.6200 415.6800 ;
      RECT 1017.4800 414.2000 1062.9600 423.5000 ;
      RECT 1007.4200 414.2000 1015.2800 423.5000 ;
      RECT 2436.3200 413.9400 2444.2800 423.2400 ;
      RECT 2388.9400 413.9400 2434.1200 423.2400 ;
      RECT 2168.7200 413.9400 2384.1400 415.3350 ;
      RECT 1728.2800 413.9400 1943.7000 415.3350 ;
      RECT 1508.0600 413.9400 1723.4800 415.3350 ;
      RECT 1287.9800 413.9400 1503.2600 415.3350 ;
      RECT 1057.5000 402.0000 1062.9600 414.2000 ;
      RECT 1055.1000 402.0000 1055.3000 414.2000 ;
      RECT 1017.4800 402.0000 1052.9000 414.2000 ;
      RECT 1015.0800 402.0000 1015.2800 414.2000 ;
      RECT 2438.9200 401.7400 2444.2800 413.9400 ;
      RECT 2436.3200 401.7400 2436.7200 413.9400 ;
      RECT 2398.9000 401.7400 2434.1200 413.9400 ;
      RECT 2396.3000 401.7400 2396.7000 413.9400 ;
      RECT 2378.7800 401.7400 2384.1400 413.9400 ;
      RECT 2376.1800 401.7400 2376.5800 413.9400 ;
      RECT 2178.6800 401.7400 2373.9800 413.9400 ;
      RECT 2176.0800 401.7400 2176.4800 413.9400 ;
      RECT 1938.3400 401.7400 1943.7000 413.9400 ;
      RECT 1935.7400 401.7400 1936.1400 413.9400 ;
      RECT 1738.2400 401.7400 1933.5400 413.9400 ;
      RECT 1735.6400 401.7400 1736.0400 413.9400 ;
      RECT 1718.1200 401.7400 1723.4800 413.9400 ;
      RECT 1715.5200 401.7400 1715.9200 413.9400 ;
      RECT 1518.0200 401.7400 1713.3200 413.9400 ;
      RECT 1515.4200 401.7400 1515.8200 413.9400 ;
      RECT 1497.9000 401.7400 1503.2600 413.9400 ;
      RECT 1495.3000 401.7400 1495.7000 413.9400 ;
      RECT 1297.8000 401.7400 1493.1000 413.9400 ;
      RECT 1295.2000 401.7400 1295.6000 413.9400 ;
      RECT 1015.0800 391.3400 1062.9600 402.0000 ;
      RECT 1007.4200 391.3400 1012.8800 414.2000 ;
      RECT 2396.3000 391.0800 2444.2800 401.7400 ;
      RECT 2388.9400 391.0800 2394.1000 413.9400 ;
      RECT 2176.0800 391.0800 2384.1400 401.7400 ;
      RECT 2168.7200 391.0800 2173.8800 413.9400 ;
      RECT 1735.6400 391.0800 1943.7000 401.7400 ;
      RECT 1728.2800 391.0800 1733.4400 413.9400 ;
      RECT 1515.4200 391.0800 1723.4800 401.7400 ;
      RECT 1508.0600 391.0800 1513.2200 413.9400 ;
      RECT 1295.2000 391.0800 1503.2600 401.7400 ;
      RECT 1287.9800 391.0800 1293.0000 413.9400 ;
      RECT 1067.7600 193.8600 1283.0400 619.8200 ;
      RECT 1007.4200 193.8600 1062.9600 391.3400 ;
      RECT 2388.9400 193.6000 2444.2800 391.0800 ;
      RECT 2168.7200 193.6000 2384.1400 391.0800 ;
      RECT 1948.5000 193.6000 2163.9200 619.5600 ;
      RECT 1728.2800 193.6000 1943.7000 391.0800 ;
      RECT 1508.0600 193.6000 1723.4800 391.0800 ;
      RECT 1287.9800 193.6000 1503.2600 391.0800 ;
      RECT 1077.7200 185.9550 1283.0400 193.8600 ;
      RECT 1067.7600 185.9550 1075.5200 193.8600 ;
      RECT 2178.6800 185.6950 2384.1400 193.6000 ;
      RECT 2168.7200 185.6950 2176.4800 193.6000 ;
      RECT 1958.4600 185.6950 2163.9200 193.6000 ;
      RECT 1948.5000 185.6950 1956.2600 193.6000 ;
      RECT 1738.2400 185.6950 1943.7000 193.6000 ;
      RECT 1728.2800 185.6950 1736.0400 193.6000 ;
      RECT 1518.0200 185.6950 1723.4800 193.6000 ;
      RECT 1508.0600 185.6950 1515.8200 193.6000 ;
      RECT 1297.8000 185.6950 1503.2600 193.6000 ;
      RECT 1287.9800 185.6950 1295.6000 193.6000 ;
      RECT 1067.7600 184.5600 1283.0400 185.9550 ;
      RECT 1017.4800 184.5600 1062.9600 193.8600 ;
      RECT 1007.4200 184.5600 1015.2800 193.8600 ;
      RECT 2436.3200 184.3000 2444.2800 193.6000 ;
      RECT 2388.9400 184.3000 2434.1200 193.6000 ;
      RECT 2168.7200 184.3000 2384.1400 185.6950 ;
      RECT 1948.5000 184.3000 2163.9200 185.6950 ;
      RECT 1728.2800 184.3000 1943.7000 185.6950 ;
      RECT 1508.0600 184.3000 1723.4800 185.6950 ;
      RECT 1287.9800 184.3000 1503.2600 185.6950 ;
      RECT 1275.2200 179.3000 1275.6200 184.5600 ;
      RECT 1075.1200 179.3000 1075.5200 184.5600 ;
      RECT 2376.1800 178.9700 2376.5800 184.3000 ;
      RECT 2176.0800 178.9700 2176.4800 184.3000 ;
      RECT 2155.9600 178.9700 2156.3600 184.3000 ;
      RECT 1955.8600 178.9700 1956.2600 184.3000 ;
      RECT 1935.7400 178.9700 1936.1400 184.3000 ;
      RECT 1735.6400 178.9700 1736.0400 184.3000 ;
      RECT 1715.5200 178.9700 1715.9200 184.3000 ;
      RECT 1515.4200 178.9700 1515.8200 184.3000 ;
      RECT 1495.3000 178.9700 1495.7000 184.3000 ;
      RECT 1295.2000 178.9700 1295.6000 184.3000 ;
      RECT 1077.7200 178.5600 1273.0200 184.5600 ;
      RECT 1055.1000 178.5600 1055.3000 184.5600 ;
      RECT 1017.4800 178.5600 1052.9000 184.5600 ;
      RECT 1015.0800 178.5600 1015.2800 184.5600 ;
      RECT 1007.4200 178.5600 1012.8800 184.5600 ;
      RECT 1004.8200 178.5600 1005.2200 2564.0200 ;
      RECT 665.0200 178.5600 665.4200 637.4400 ;
      RECT 507.4200 178.5600 662.8200 456.9200 ;
      RECT 504.8200 178.5600 505.2200 637.4400 ;
      RECT 2436.3200 178.3000 2436.7200 184.3000 ;
      RECT 2398.9000 178.3000 2434.1200 184.3000 ;
      RECT 2396.3000 178.3000 2396.7000 184.3000 ;
      RECT 2178.6800 178.3000 2373.9800 184.3000 ;
      RECT 1958.4600 178.3000 2153.7600 184.3000 ;
      RECT 1738.2400 178.3000 1933.5400 184.3000 ;
      RECT 1518.0200 178.3000 1713.3200 184.3000 ;
      RECT 1297.8000 178.3000 1493.1000 184.3000 ;
      RECT 1275.3200 178.1600 1275.6200 179.3000 ;
      RECT 1075.1200 178.1600 1075.4200 179.3000 ;
      RECT 2376.2800 177.9000 2376.5800 178.9700 ;
      RECT 2176.0800 177.9000 2176.3800 178.9700 ;
      RECT 2156.0600 177.9000 2156.3600 178.9700 ;
      RECT 1955.8600 177.9000 1956.1600 178.9700 ;
      RECT 1935.8400 177.9000 1936.1400 178.9700 ;
      RECT 1735.6400 177.9000 1735.9400 178.9700 ;
      RECT 1715.6200 177.9000 1715.9200 178.9700 ;
      RECT 1515.4200 177.9000 1515.7200 178.9700 ;
      RECT 1495.4000 177.9000 1495.7000 178.9700 ;
      RECT 1295.2000 177.9000 1295.5000 178.9700 ;
      RECT 1277.8200 177.4800 1283.0400 184.5600 ;
      RECT 1067.7600 177.4800 1072.9200 184.5600 ;
      RECT 2378.7800 177.0100 2384.1400 184.3000 ;
      RECT 2168.7200 177.0100 2173.8800 184.3000 ;
      RECT 2158.5600 177.0100 2163.9200 184.3000 ;
      RECT 1948.5000 177.0100 1953.6600 184.3000 ;
      RECT 1938.3400 177.0100 1943.7000 184.3000 ;
      RECT 1728.2800 177.0100 1733.4400 184.3000 ;
      RECT 1718.1200 177.0100 1723.4800 184.3000 ;
      RECT 1508.0600 177.0100 1513.2200 184.3000 ;
      RECT 1497.9000 177.0100 1503.2600 184.3000 ;
      RECT 1287.9800 177.0100 1293.0000 184.3000 ;
      RECT 1057.5000 175.9600 1062.9600 184.5600 ;
      RECT 1015.0800 175.9600 1055.3000 178.5600 ;
      RECT 1004.8200 175.9600 1012.8800 178.5600 ;
      RECT 667.6200 175.9600 1002.6200 635.2400 ;
      RECT 504.8200 175.9600 665.4200 178.5600 ;
      RECT 9.3000 175.9600 502.6200 635.2400 ;
      RECT 2438.9200 175.7000 2444.2800 184.3000 ;
      RECT 2396.3000 175.7000 2436.7200 178.3000 ;
      RECT 2388.9400 175.7000 2394.1000 184.3000 ;
      RECT 1277.7200 172.3600 1283.0400 177.4800 ;
      RECT 1275.3200 172.3600 1275.5200 178.1600 ;
      RECT 1077.6200 172.3600 1273.1200 178.5600 ;
      RECT 1075.2200 172.3600 1075.4200 178.1600 ;
      RECT 2378.6800 172.1000 2384.1400 177.0100 ;
      RECT 2376.2800 172.1000 2376.4800 177.9000 ;
      RECT 2178.5800 172.1000 2374.0800 178.3000 ;
      RECT 2176.1800 172.1000 2176.3800 177.9000 ;
      RECT 2158.4600 172.1000 2163.9200 177.0100 ;
      RECT 2156.0600 172.1000 2156.2600 177.9000 ;
      RECT 1958.3600 172.1000 2153.8600 178.3000 ;
      RECT 1955.9600 172.1000 1956.1600 177.9000 ;
      RECT 1938.2400 172.1000 1943.7000 177.0100 ;
      RECT 1935.8400 172.1000 1936.0400 177.9000 ;
      RECT 1738.1400 172.1000 1933.6400 178.3000 ;
      RECT 1735.7400 172.1000 1735.9400 177.9000 ;
      RECT 1718.0200 172.1000 1723.4800 177.0100 ;
      RECT 1715.6200 172.1000 1715.8200 177.9000 ;
      RECT 1517.9200 172.1000 1713.4200 178.3000 ;
      RECT 1515.5200 172.1000 1515.7200 177.9000 ;
      RECT 1497.8000 172.1000 1503.2600 177.0100 ;
      RECT 1495.4000 172.1000 1495.6000 177.9000 ;
      RECT 1297.7000 172.1000 1493.2000 178.3000 ;
      RECT 1295.3000 172.1000 1295.5000 177.9000 ;
      RECT 1075.2200 163.4000 1283.0400 172.3600 ;
      RECT 1067.7600 163.4000 1073.0200 177.4800 ;
      RECT 2176.1800 163.1400 2384.1400 172.1000 ;
      RECT 2168.7200 163.1400 2173.9800 177.0100 ;
      RECT 1955.9600 163.1400 2163.9200 172.1000 ;
      RECT 1948.5000 163.1400 1953.7600 177.0100 ;
      RECT 1735.7400 163.1400 1943.7000 172.1000 ;
      RECT 1728.2800 163.1400 1733.5400 177.0100 ;
      RECT 1515.5200 163.1400 1723.4800 172.1000 ;
      RECT 1508.0600 163.1400 1513.3200 177.0100 ;
      RECT 1295.3000 163.1400 1503.2600 172.1000 ;
      RECT 1287.9800 163.1400 1293.1000 177.0100 ;
      RECT 1067.7600 150.8800 1283.0400 163.4000 ;
      RECT 2168.7200 150.6200 2384.1400 163.1400 ;
      RECT 1948.5000 150.6200 2163.9200 163.1400 ;
      RECT 1728.2800 150.6200 1943.7000 163.1400 ;
      RECT 1508.0600 150.6200 1723.4800 163.1400 ;
      RECT 1287.9800 150.6200 1503.2600 163.1400 ;
      RECT 1275.3200 144.3000 1283.0400 150.8800 ;
      RECT 1067.7600 144.3000 1273.1200 150.8800 ;
      RECT 2376.2800 144.0400 2384.1400 150.6200 ;
      RECT 2168.7200 144.0400 2374.0800 150.6200 ;
      RECT 2156.0600 144.0400 2163.9200 150.6200 ;
      RECT 1948.5000 144.0400 2153.8600 150.6200 ;
      RECT 1935.8400 144.0400 1943.7000 150.6200 ;
      RECT 1728.2800 144.0400 1933.6400 150.6200 ;
      RECT 1715.6200 144.0400 1723.4800 150.6200 ;
      RECT 1508.0600 144.0400 1713.4200 150.6200 ;
      RECT 1495.4000 144.0400 1503.2600 150.6200 ;
      RECT 1287.9800 144.0400 1493.2000 150.6200 ;
      RECT 1275.3200 138.3000 1275.5200 144.3000 ;
      RECT 1077.6200 138.3000 1273.1200 144.3000 ;
      RECT 1075.2200 138.3000 1075.4200 144.3000 ;
      RECT 2388.9400 138.2400 2444.2800 175.7000 ;
      RECT 2376.2800 138.0400 2376.4800 144.0400 ;
      RECT 2178.5800 138.0400 2374.0800 144.0400 ;
      RECT 2176.1800 138.0400 2176.3800 144.0400 ;
      RECT 2156.0600 138.0400 2156.2600 144.0400 ;
      RECT 1958.3600 138.0400 2153.8600 144.0400 ;
      RECT 1955.9600 138.0400 1956.1600 144.0400 ;
      RECT 1935.8400 138.0400 1936.0400 144.0400 ;
      RECT 1738.1400 138.0400 1933.6400 144.0400 ;
      RECT 1735.7400 138.0400 1735.9400 144.0400 ;
      RECT 1715.6200 138.0400 1715.8200 144.0400 ;
      RECT 1517.9200 138.0400 1713.4200 144.0400 ;
      RECT 1515.5200 138.0400 1515.7200 144.0400 ;
      RECT 1495.4000 138.0400 1495.6000 144.0400 ;
      RECT 1297.7000 138.0400 1493.2000 144.0400 ;
      RECT 1295.3000 138.0400 1295.5000 144.0400 ;
      RECT 2390.3000 137.1600 2444.2800 138.2400 ;
      RECT 1277.7200 135.7000 1283.0400 144.3000 ;
      RECT 1075.2200 135.7000 1275.5200 138.3000 ;
      RECT 1067.7600 135.7000 1073.0200 144.3000 ;
      RECT 2378.6800 135.4400 2384.1400 144.0400 ;
      RECT 2176.1800 135.4400 2376.4800 138.0400 ;
      RECT 2168.7200 135.4400 2173.9800 144.0400 ;
      RECT 2158.4600 135.4400 2163.9200 144.0400 ;
      RECT 1955.9600 135.4400 2156.2600 138.0400 ;
      RECT 1948.5000 135.4400 1953.7600 144.0400 ;
      RECT 1938.2400 135.4400 1943.7000 144.0400 ;
      RECT 1735.7400 135.4400 1936.0400 138.0400 ;
      RECT 1728.2800 135.4400 1733.5400 144.0400 ;
      RECT 1718.0200 135.4400 1723.4800 144.0400 ;
      RECT 1515.5200 135.4400 1715.8200 138.0400 ;
      RECT 1508.0600 135.4400 1513.3200 144.0400 ;
      RECT 1497.8000 135.4400 1503.2600 144.0400 ;
      RECT 1295.3000 135.4400 1495.6000 138.0400 ;
      RECT 1287.9800 135.4400 1293.1000 144.0400 ;
      RECT 3364.7200 5.7000 3365.1200 2564.0200 ;
      RECT 3307.6200 5.7000 3361.1200 2564.0200 ;
      RECT 3305.0200 5.7000 3305.4200 2564.0200 ;
      RECT 2494.8200 5.7000 2495.2200 2564.0200 ;
      RECT 2449.0800 5.7000 2492.6200 414.6000 ;
      RECT 2446.4800 5.7000 2446.8800 2564.0200 ;
      RECT 2388.9400 5.7000 2444.2800 137.1600 ;
      RECT 2386.3400 5.7000 2386.7400 2564.0200 ;
      RECT 2168.7200 5.7000 2384.1400 135.4400 ;
      RECT 2166.1200 5.7000 2166.5200 2564.0200 ;
      RECT 1948.5000 5.7000 2163.9200 135.4400 ;
      RECT 1945.9000 5.7000 1946.3000 2564.0200 ;
      RECT 1728.2800 5.7000 1943.7000 135.4400 ;
      RECT 1725.6800 5.7000 1726.0800 2564.0200 ;
      RECT 1508.0600 5.7000 1723.4800 135.4400 ;
      RECT 1505.4600 5.7000 1505.8600 2564.0200 ;
      RECT 1287.9800 5.7000 1503.2600 135.4400 ;
      RECT 1285.3800 5.7000 1285.6400 2564.0200 ;
      RECT 1067.7600 5.7000 1283.0400 135.7000 ;
      RECT 1065.1600 5.7000 1065.5600 2564.0200 ;
      RECT 9.3000 5.7000 1062.9600 175.9600 ;
      RECT 5.3000 5.7000 5.7000 2564.0200 ;
      RECT 3368.7200 1.7000 3370.4200 2568.0200 ;
      RECT 3305.0200 1.7000 3365.1200 5.7000 ;
      RECT 2497.4200 1.7000 3302.8200 1905.6000 ;
      RECT 2446.4800 1.7000 2495.2200 5.7000 ;
      RECT 2386.3400 1.7000 2444.2800 5.7000 ;
      RECT 2166.1200 1.7000 2384.1400 5.7000 ;
      RECT 1945.9000 1.7000 2163.9200 5.7000 ;
      RECT 1725.6800 1.7000 1943.7000 5.7000 ;
      RECT 1505.4600 1.7000 1723.4800 5.7000 ;
      RECT 1285.3800 1.7000 1503.2600 5.7000 ;
      RECT 1065.1600 1.7000 1283.0400 5.7000 ;
      RECT 5.3000 1.7000 1062.9600 5.7000 ;
      RECT 0.0000 1.7000 1.7000 2568.0200 ;
      RECT 0.0000 1.1000 3370.4200 1.7000 ;
      RECT 649.0500 0.0000 3370.4200 1.1000 ;
      RECT 0.0000 0.0000 648.1500 1.1000 ;
  END
END eFPGA_CPU_top

END LIBRARY
