VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.920 900.000 300.520 ;
    END
  END clk
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.130 0.000 862.410 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 0.000 187.590 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 0.000 787.430 4.000 ;
    END
  END la_data_out[9]
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 4.000 ;
    END
  END wb_rst_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 587.520 ;
    END
  END vssa2
  OBS
      LAYER nwell ;
        RECT 5.330 586.105 894.430 587.710 ;
        RECT 5.330 580.665 894.430 583.495 ;
        RECT 5.330 575.225 894.430 578.055 ;
        RECT 5.330 569.785 894.430 572.615 ;
        RECT 5.330 564.345 894.430 567.175 ;
        RECT 5.330 558.905 894.430 561.735 ;
        RECT 5.330 553.465 894.430 556.295 ;
        RECT 5.330 548.025 894.430 550.855 ;
        RECT 5.330 542.585 894.430 545.415 ;
        RECT 5.330 537.145 894.430 539.975 ;
        RECT 5.330 531.705 894.430 534.535 ;
        RECT 5.330 526.265 894.430 529.095 ;
        RECT 5.330 520.825 894.430 523.655 ;
        RECT 5.330 515.385 894.430 518.215 ;
        RECT 5.330 509.945 894.430 512.775 ;
        RECT 5.330 504.505 894.430 507.335 ;
        RECT 5.330 499.065 894.430 501.895 ;
        RECT 5.330 493.625 894.430 496.455 ;
        RECT 5.330 488.185 894.430 491.015 ;
        RECT 5.330 482.745 894.430 485.575 ;
        RECT 5.330 477.305 894.430 480.135 ;
        RECT 5.330 471.865 894.430 474.695 ;
        RECT 5.330 466.425 894.430 469.255 ;
        RECT 5.330 460.985 894.430 463.815 ;
        RECT 5.330 455.545 894.430 458.375 ;
        RECT 5.330 450.105 894.430 452.935 ;
        RECT 5.330 444.665 894.430 447.495 ;
        RECT 5.330 439.225 894.430 442.055 ;
        RECT 5.330 433.785 894.430 436.615 ;
        RECT 5.330 428.345 894.430 431.175 ;
        RECT 5.330 422.905 894.430 425.735 ;
        RECT 5.330 417.465 894.430 420.295 ;
        RECT 5.330 412.025 894.430 414.855 ;
        RECT 5.330 406.585 894.430 409.415 ;
        RECT 5.330 401.145 894.430 403.975 ;
        RECT 5.330 395.705 894.430 398.535 ;
        RECT 5.330 390.265 894.430 393.095 ;
        RECT 5.330 384.825 894.430 387.655 ;
        RECT 5.330 379.385 894.430 382.215 ;
        RECT 5.330 373.945 894.430 376.775 ;
        RECT 5.330 368.505 894.430 371.335 ;
        RECT 5.330 363.065 894.430 365.895 ;
        RECT 5.330 357.625 894.430 360.455 ;
        RECT 5.330 352.185 894.430 355.015 ;
        RECT 5.330 346.745 894.430 349.575 ;
        RECT 5.330 341.305 894.430 344.135 ;
        RECT 5.330 335.865 894.430 338.695 ;
        RECT 5.330 330.425 894.430 333.255 ;
        RECT 5.330 324.985 894.430 327.815 ;
        RECT 5.330 319.545 894.430 322.375 ;
        RECT 5.330 314.105 894.430 316.935 ;
        RECT 5.330 308.665 894.430 311.495 ;
        RECT 5.330 303.225 894.430 306.055 ;
        RECT 5.330 297.785 894.430 300.615 ;
        RECT 5.330 292.345 894.430 295.175 ;
        RECT 5.330 286.905 894.430 289.735 ;
        RECT 5.330 281.465 894.430 284.295 ;
        RECT 5.330 276.025 894.430 278.855 ;
        RECT 5.330 270.585 894.430 273.415 ;
        RECT 5.330 265.145 894.430 267.975 ;
        RECT 5.330 259.705 894.430 262.535 ;
        RECT 5.330 254.265 894.430 257.095 ;
        RECT 5.330 248.825 894.430 251.655 ;
        RECT 5.330 243.385 894.430 246.215 ;
        RECT 5.330 237.945 894.430 240.775 ;
        RECT 5.330 232.505 894.430 235.335 ;
        RECT 5.330 227.065 894.430 229.895 ;
        RECT 5.330 221.625 894.430 224.455 ;
        RECT 5.330 216.185 894.430 219.015 ;
        RECT 5.330 210.745 894.430 213.575 ;
        RECT 5.330 205.305 894.430 208.135 ;
        RECT 5.330 199.865 894.430 202.695 ;
        RECT 5.330 194.425 894.430 197.255 ;
        RECT 5.330 188.985 894.430 191.815 ;
        RECT 5.330 183.545 894.430 186.375 ;
        RECT 5.330 178.105 894.430 180.935 ;
        RECT 5.330 172.665 894.430 175.495 ;
        RECT 5.330 167.225 894.430 170.055 ;
        RECT 5.330 161.785 894.430 164.615 ;
        RECT 5.330 156.345 894.430 159.175 ;
        RECT 5.330 150.905 894.430 153.735 ;
        RECT 5.330 145.465 894.430 148.295 ;
        RECT 5.330 140.025 894.430 142.855 ;
        RECT 5.330 134.585 894.430 137.415 ;
        RECT 5.330 129.145 894.430 131.975 ;
        RECT 5.330 123.705 894.430 126.535 ;
        RECT 5.330 118.265 894.430 121.095 ;
        RECT 5.330 112.825 894.430 115.655 ;
        RECT 5.330 107.385 894.430 110.215 ;
        RECT 5.330 101.945 894.430 104.775 ;
        RECT 5.330 96.505 894.430 99.335 ;
        RECT 5.330 91.065 894.430 93.895 ;
        RECT 5.330 85.625 894.430 88.455 ;
        RECT 5.330 80.185 894.430 83.015 ;
        RECT 5.330 74.745 894.430 77.575 ;
        RECT 5.330 69.305 894.430 72.135 ;
        RECT 5.330 63.865 894.430 66.695 ;
        RECT 5.330 58.425 894.430 61.255 ;
        RECT 5.330 52.985 894.430 55.815 ;
        RECT 5.330 47.545 894.430 50.375 ;
        RECT 5.330 42.105 894.430 44.935 ;
        RECT 5.330 36.665 894.430 39.495 ;
        RECT 5.330 31.225 894.430 34.055 ;
        RECT 5.330 25.785 894.430 28.615 ;
        RECT 5.330 20.345 894.430 23.175 ;
        RECT 5.330 14.905 894.430 17.735 ;
        RECT 5.330 10.690 894.430 12.295 ;
      LAYER li1 ;
        RECT 5.520 10.795 894.240 587.605 ;
      LAYER met1 ;
        RECT 5.520 10.640 894.240 587.760 ;
      LAYER met2 ;
        RECT 21.100 4.280 879.890 587.760 ;
        RECT 21.100 4.000 37.070 4.280 ;
        RECT 37.910 4.000 112.050 4.280 ;
        RECT 112.890 4.000 187.030 4.280 ;
        RECT 187.870 4.000 262.010 4.280 ;
        RECT 262.850 4.000 336.990 4.280 ;
        RECT 337.830 4.000 411.970 4.280 ;
        RECT 412.810 4.000 486.950 4.280 ;
        RECT 487.790 4.000 561.930 4.280 ;
        RECT 562.770 4.000 636.910 4.280 ;
        RECT 637.750 4.000 711.890 4.280 ;
        RECT 712.730 4.000 786.870 4.280 ;
        RECT 787.710 4.000 861.850 4.280 ;
        RECT 862.690 4.000 879.890 4.280 ;
      LAYER met3 ;
        RECT 21.040 300.920 896.000 587.685 ;
        RECT 21.040 299.520 895.600 300.920 ;
        RECT 21.040 10.715 896.000 299.520 ;
      LAYER met4 ;
        RECT 286.415 50.495 327.840 238.505 ;
        RECT 330.240 50.495 331.140 238.505 ;
        RECT 333.540 50.495 334.440 238.505 ;
        RECT 336.840 50.495 337.740 238.505 ;
        RECT 340.140 50.495 404.640 238.505 ;
        RECT 407.040 50.495 407.940 238.505 ;
        RECT 410.340 50.495 411.240 238.505 ;
        RECT 413.640 50.495 414.540 238.505 ;
        RECT 416.940 50.495 433.945 238.505 ;
  END
END user_proj_example
END LIBRARY

