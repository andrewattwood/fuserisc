// SPDX-FileCopyrightText: 2020 Nguyen Dao
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0


	//External IO ports exported directly from the corresponding tiles
module eFPGA (Tile_X0Y1_OPA_I0, Tile_X0Y1_OPA_I1, Tile_X0Y1_OPA_I2, Tile_X0Y1_OPA_I3, UserCLK, Tile_X0Y1_OPB_I0, Tile_X0Y1_OPB_I1, Tile_X0Y1_OPB_I2, Tile_X0Y1_OPB_I3, Tile_X0Y1_RES0_O0, Tile_X0Y1_RES0_O1, Tile_X0Y1_RES0_O2, Tile_X0Y1_RES0_O3, Tile_X0Y1_RES1_O0, Tile_X0Y1_RES1_O1, Tile_X0Y1_RES1_O2, Tile_X0Y1_RES1_O3, Tile_X0Y1_RES2_O0, Tile_X0Y1_RES2_O1, Tile_X0Y1_RES2_O2, Tile_X0Y1_RES2_O3, Tile_X7Y1_OPA_I0, Tile_X7Y1_OPA_I1, Tile_X7Y1_OPA_I2, Tile_X7Y1_OPA_I3, Tile_X7Y1_OPB_I0, Tile_X7Y1_OPB_I1, Tile_X7Y1_OPB_I2, Tile_X7Y1_OPB_I3, Tile_X7Y1_RES0_O0, Tile_X7Y1_RES0_O1, Tile_X7Y1_RES0_O2, Tile_X7Y1_RES0_O3, Tile_X7Y1_RES1_O0, Tile_X7Y1_RES1_O1, Tile_X7Y1_RES1_O2, Tile_X7Y1_RES1_O3, Tile_X7Y1_RES2_O0, Tile_X7Y1_RES2_O1, Tile_X7Y1_RES2_O2, Tile_X7Y1_RES2_O3, Tile_X0Y2_OPA_I0, Tile_X0Y2_OPA_I1, Tile_X0Y2_OPA_I2, Tile_X0Y2_OPA_I3, Tile_X0Y2_OPB_I0, Tile_X0Y2_OPB_I1, Tile_X0Y2_OPB_I2, Tile_X0Y2_OPB_I3, Tile_X0Y2_RES0_O0, Tile_X0Y2_RES0_O1, Tile_X0Y2_RES0_O2, Tile_X0Y2_RES0_O3, Tile_X0Y2_RES1_O0, Tile_X0Y2_RES1_O1, Tile_X0Y2_RES1_O2, Tile_X0Y2_RES1_O3, Tile_X0Y2_RES2_O0, Tile_X0Y2_RES2_O1, Tile_X0Y2_RES2_O2, Tile_X0Y2_RES2_O3, Tile_X7Y2_OPA_I0, Tile_X7Y2_OPA_I1, Tile_X7Y2_OPA_I2, Tile_X7Y2_OPA_I3, Tile_X7Y2_OPB_I0, Tile_X7Y2_OPB_I1, Tile_X7Y2_OPB_I2, Tile_X7Y2_OPB_I3, Tile_X7Y2_RES0_O0, Tile_X7Y2_RES0_O1, Tile_X7Y2_RES0_O2, Tile_X7Y2_RES0_O3, Tile_X7Y2_RES1_O0, Tile_X7Y2_RES1_O1, Tile_X7Y2_RES1_O2, Tile_X7Y2_RES1_O3, Tile_X7Y2_RES2_O0, Tile_X7Y2_RES2_O1, Tile_X7Y2_RES2_O2, Tile_X7Y2_RES2_O3, Tile_X0Y3_OPA_I0, Tile_X0Y3_OPA_I1, Tile_X0Y3_OPA_I2, Tile_X0Y3_OPA_I3, Tile_X0Y3_OPB_I0, Tile_X0Y3_OPB_I1, Tile_X0Y3_OPB_I2, Tile_X0Y3_OPB_I3, Tile_X0Y3_RES0_O0, Tile_X0Y3_RES0_O1, Tile_X0Y3_RES0_O2, Tile_X0Y3_RES0_O3, Tile_X0Y3_RES1_O0, Tile_X0Y3_RES1_O1, Tile_X0Y3_RES1_O2, Tile_X0Y3_RES1_O3, Tile_X0Y3_RES2_O0, Tile_X0Y3_RES2_O1, Tile_X0Y3_RES2_O2, Tile_X0Y3_RES2_O3, Tile_X7Y3_OPA_I0, Tile_X7Y3_OPA_I1, Tile_X7Y3_OPA_I2, Tile_X7Y3_OPA_I3, Tile_X7Y3_OPB_I0, Tile_X7Y3_OPB_I1, Tile_X7Y3_OPB_I2, Tile_X7Y3_OPB_I3, Tile_X7Y3_RES0_O0, Tile_X7Y3_RES0_O1, Tile_X7Y3_RES0_O2, Tile_X7Y3_RES0_O3, Tile_X7Y3_RES1_O0, Tile_X7Y3_RES1_O1, Tile_X7Y3_RES1_O2, Tile_X7Y3_RES1_O3, Tile_X7Y3_RES2_O0, Tile_X7Y3_RES2_O1, Tile_X7Y3_RES2_O2, Tile_X7Y3_RES2_O3, Tile_X0Y4_OPA_I0, Tile_X0Y4_OPA_I1, Tile_X0Y4_OPA_I2, Tile_X0Y4_OPA_I3, Tile_X0Y4_OPB_I0, Tile_X0Y4_OPB_I1, Tile_X0Y4_OPB_I2, Tile_X0Y4_OPB_I3, Tile_X0Y4_RES0_O0, Tile_X0Y4_RES0_O1, Tile_X0Y4_RES0_O2, Tile_X0Y4_RES0_O3, Tile_X0Y4_RES1_O0, Tile_X0Y4_RES1_O1, Tile_X0Y4_RES1_O2, Tile_X0Y4_RES1_O3, Tile_X0Y4_RES2_O0, Tile_X0Y4_RES2_O1, Tile_X0Y4_RES2_O2, Tile_X0Y4_RES2_O3, Tile_X7Y4_OPA_I0, Tile_X7Y4_OPA_I1, Tile_X7Y4_OPA_I2, Tile_X7Y4_OPA_I3, Tile_X7Y4_OPB_I0, Tile_X7Y4_OPB_I1, Tile_X7Y4_OPB_I2, Tile_X7Y4_OPB_I3, Tile_X7Y4_RES0_O0, Tile_X7Y4_RES0_O1, Tile_X7Y4_RES0_O2, Tile_X7Y4_RES0_O3, Tile_X7Y4_RES1_O0, Tile_X7Y4_RES1_O1, Tile_X7Y4_RES1_O2, Tile_X7Y4_RES1_O3, Tile_X7Y4_RES2_O0, Tile_X7Y4_RES2_O1, Tile_X7Y4_RES2_O2, Tile_X7Y4_RES2_O3, Tile_X0Y5_OPA_I0, Tile_X0Y5_OPA_I1, Tile_X0Y5_OPA_I2, Tile_X0Y5_OPA_I3, Tile_X0Y5_OPB_I0, Tile_X0Y5_OPB_I1, Tile_X0Y5_OPB_I2, Tile_X0Y5_OPB_I3, Tile_X0Y5_RES0_O0, Tile_X0Y5_RES0_O1, Tile_X0Y5_RES0_O2, Tile_X0Y5_RES0_O3, Tile_X0Y5_RES1_O0, Tile_X0Y5_RES1_O1, Tile_X0Y5_RES1_O2, Tile_X0Y5_RES1_O3, Tile_X0Y5_RES2_O0, Tile_X0Y5_RES2_O1, Tile_X0Y5_RES2_O2, Tile_X0Y5_RES2_O3, Tile_X7Y5_OPA_I0, Tile_X7Y5_OPA_I1, Tile_X7Y5_OPA_I2, Tile_X7Y5_OPA_I3, Tile_X7Y5_OPB_I0, Tile_X7Y5_OPB_I1, Tile_X7Y5_OPB_I2, Tile_X7Y5_OPB_I3, Tile_X7Y5_RES0_O0, Tile_X7Y5_RES0_O1, Tile_X7Y5_RES0_O2, Tile_X7Y5_RES0_O3, Tile_X7Y5_RES1_O0, Tile_X7Y5_RES1_O1, Tile_X7Y5_RES1_O2, Tile_X7Y5_RES1_O3, Tile_X7Y5_RES2_O0, Tile_X7Y5_RES2_O1, Tile_X7Y5_RES2_O2, Tile_X7Y5_RES2_O3, Tile_X0Y6_OPA_I0, Tile_X0Y6_OPA_I1, Tile_X0Y6_OPA_I2, Tile_X0Y6_OPA_I3, Tile_X0Y6_OPB_I0, Tile_X0Y6_OPB_I1, Tile_X0Y6_OPB_I2, Tile_X0Y6_OPB_I3, Tile_X0Y6_RES0_O0, Tile_X0Y6_RES0_O1, Tile_X0Y6_RES0_O2, Tile_X0Y6_RES0_O3, Tile_X0Y6_RES1_O0, Tile_X0Y6_RES1_O1, Tile_X0Y6_RES1_O2, Tile_X0Y6_RES1_O3, Tile_X0Y6_RES2_O0, Tile_X0Y6_RES2_O1, Tile_X0Y6_RES2_O2, Tile_X0Y6_RES2_O3, Tile_X7Y6_OPA_I0, Tile_X7Y6_OPA_I1, Tile_X7Y6_OPA_I2, Tile_X7Y6_OPA_I3, Tile_X7Y6_OPB_I0, Tile_X7Y6_OPB_I1, Tile_X7Y6_OPB_I2, Tile_X7Y6_OPB_I3, Tile_X7Y6_RES0_O0, Tile_X7Y6_RES0_O1, Tile_X7Y6_RES0_O2, Tile_X7Y6_RES0_O3, Tile_X7Y6_RES1_O0, Tile_X7Y6_RES1_O1, Tile_X7Y6_RES1_O2, Tile_X7Y6_RES1_O3, Tile_X7Y6_RES2_O0, Tile_X7Y6_RES2_O1, Tile_X7Y6_RES2_O2, Tile_X7Y6_RES2_O3, Tile_X0Y7_OPA_I0, Tile_X0Y7_OPA_I1, Tile_X0Y7_OPA_I2, Tile_X0Y7_OPA_I3, Tile_X0Y7_OPB_I0, Tile_X0Y7_OPB_I1, Tile_X0Y7_OPB_I2, Tile_X0Y7_OPB_I3, Tile_X0Y7_RES0_O0, Tile_X0Y7_RES0_O1, Tile_X0Y7_RES0_O2, Tile_X0Y7_RES0_O3, Tile_X0Y7_RES1_O0, Tile_X0Y7_RES1_O1, Tile_X0Y7_RES1_O2, Tile_X0Y7_RES1_O3, Tile_X0Y7_RES2_O0, Tile_X0Y7_RES2_O1, Tile_X0Y7_RES2_O2, Tile_X0Y7_RES2_O3, Tile_X7Y7_OPA_I0, Tile_X7Y7_OPA_I1, Tile_X7Y7_OPA_I2, Tile_X7Y7_OPA_I3, Tile_X7Y7_OPB_I0, Tile_X7Y7_OPB_I1, Tile_X7Y7_OPB_I2, Tile_X7Y7_OPB_I3, Tile_X7Y7_RES0_O0, Tile_X7Y7_RES0_O1, Tile_X7Y7_RES0_O2, Tile_X7Y7_RES0_O3, Tile_X7Y7_RES1_O0, Tile_X7Y7_RES1_O1, Tile_X7Y7_RES1_O2, Tile_X7Y7_RES1_O3, Tile_X7Y7_RES2_O0, Tile_X7Y7_RES2_O1, Tile_X7Y7_RES2_O2, Tile_X7Y7_RES2_O3, Tile_X0Y8_OPA_I0, Tile_X0Y8_OPA_I1, Tile_X0Y8_OPA_I2, Tile_X0Y8_OPA_I3, Tile_X0Y8_OPB_I0, Tile_X0Y8_OPB_I1, Tile_X0Y8_OPB_I2, Tile_X0Y8_OPB_I3, Tile_X0Y8_RES0_O0, Tile_X0Y8_RES0_O1, Tile_X0Y8_RES0_O2, Tile_X0Y8_RES0_O3, Tile_X0Y8_RES1_O0, Tile_X0Y8_RES1_O1, Tile_X0Y8_RES1_O2, Tile_X0Y8_RES1_O3, Tile_X0Y8_RES2_O0, Tile_X0Y8_RES2_O1, Tile_X0Y8_RES2_O2, Tile_X0Y8_RES2_O3, Tile_X7Y8_OPA_I0, Tile_X7Y8_OPA_I1, Tile_X7Y8_OPA_I2, Tile_X7Y8_OPA_I3, Tile_X7Y8_OPB_I0, Tile_X7Y8_OPB_I1, Tile_X7Y8_OPB_I2, Tile_X7Y8_OPB_I3, Tile_X7Y8_RES0_O0, Tile_X7Y8_RES0_O1, Tile_X7Y8_RES0_O2, Tile_X7Y8_RES0_O3, Tile_X7Y8_RES1_O0, Tile_X7Y8_RES1_O1, Tile_X7Y8_RES1_O2, Tile_X7Y8_RES1_O3, Tile_X7Y8_RES2_O0, Tile_X7Y8_RES2_O1, Tile_X7Y8_RES2_O2, Tile_X7Y8_RES2_O3, Tile_X0Y9_OPA_I0, Tile_X0Y9_OPA_I1, Tile_X0Y9_OPA_I2, Tile_X0Y9_OPA_I3, Tile_X0Y9_OPB_I0, Tile_X0Y9_OPB_I1, Tile_X0Y9_OPB_I2, Tile_X0Y9_OPB_I3, Tile_X0Y9_RES0_O0, Tile_X0Y9_RES0_O1, Tile_X0Y9_RES0_O2, Tile_X0Y9_RES0_O3, Tile_X0Y9_RES1_O0, Tile_X0Y9_RES1_O1, Tile_X0Y9_RES1_O2, Tile_X0Y9_RES1_O3, Tile_X0Y9_RES2_O0, Tile_X0Y9_RES2_O1, Tile_X0Y9_RES2_O2, Tile_X0Y9_RES2_O3, Tile_X7Y9_OPA_I0, Tile_X7Y9_OPA_I1, Tile_X7Y9_OPA_I2, Tile_X7Y9_OPA_I3, Tile_X7Y9_OPB_I0, Tile_X7Y9_OPB_I1, Tile_X7Y9_OPB_I2, Tile_X7Y9_OPB_I3, Tile_X7Y9_RES0_O0, Tile_X7Y9_RES0_O1, Tile_X7Y9_RES0_O2, Tile_X7Y9_RES0_O3, Tile_X7Y9_RES1_O0, Tile_X7Y9_RES1_O1, Tile_X7Y9_RES1_O2, Tile_X7Y9_RES1_O3, Tile_X7Y9_RES2_O0, Tile_X7Y9_RES2_O1, Tile_X7Y9_RES2_O2, Tile_X7Y9_RES2_O3, Tile_X0Y10_OPA_I0, Tile_X0Y10_OPA_I1, Tile_X0Y10_OPA_I2, Tile_X0Y10_OPA_I3, Tile_X0Y10_OPB_I0, Tile_X0Y10_OPB_I1, Tile_X0Y10_OPB_I2, Tile_X0Y10_OPB_I3, Tile_X0Y10_RES0_O0, Tile_X0Y10_RES0_O1, Tile_X0Y10_RES0_O2, Tile_X0Y10_RES0_O3, Tile_X0Y10_RES1_O0, Tile_X0Y10_RES1_O1, Tile_X0Y10_RES1_O2, Tile_X0Y10_RES1_O3, Tile_X0Y10_RES2_O0, Tile_X0Y10_RES2_O1, Tile_X0Y10_RES2_O2, Tile_X0Y10_RES2_O3, Tile_X7Y10_OPA_I0, Tile_X7Y10_OPA_I1, Tile_X7Y10_OPA_I2, Tile_X7Y10_OPA_I3, Tile_X7Y10_OPB_I0, Tile_X7Y10_OPB_I1, Tile_X7Y10_OPB_I2, Tile_X7Y10_OPB_I3, Tile_X7Y10_RES0_O0, Tile_X7Y10_RES0_O1, Tile_X7Y10_RES0_O2, Tile_X7Y10_RES0_O3, Tile_X7Y10_RES1_O0, Tile_X7Y10_RES1_O1, Tile_X7Y10_RES1_O2, Tile_X7Y10_RES1_O3, Tile_X7Y10_RES2_O0, Tile_X7Y10_RES2_O1, Tile_X7Y10_RES2_O2, Tile_X7Y10_RES2_O3, FrameData, FrameStrobe);
	parameter MaxFramesPerCol = 20;
	parameter FrameBitsPerRow = 32;
	parameter NoConfigBits = 0;
	input Tile_X0Y1_OPA_I0;  //EXTERNAL
	input Tile_X0Y1_OPA_I1;  //EXTERNAL
	input Tile_X0Y1_OPA_I2;  //EXTERNAL
	input Tile_X0Y1_OPA_I3;  //EXTERNAL
	input UserCLK;  //EXTERNAL //SHARED_PORT //## the EXTERNAL keyword will send this signal all the way to top and the --SHARED Allows multiple BELs usg the same port (e.g. for exportg a clock to the top)
	input Tile_X0Y1_OPB_I0;  //EXTERNAL
	input Tile_X0Y1_OPB_I1;  //EXTERNAL
	input Tile_X0Y1_OPB_I2;  //EXTERNAL
	input Tile_X0Y1_OPB_I3;  //EXTERNAL
	output Tile_X0Y1_RES0_O0;  //EXTERNAL
	output Tile_X0Y1_RES0_O1;  //EXTERNAL
	output Tile_X0Y1_RES0_O2;  //EXTERNAL
	output Tile_X0Y1_RES0_O3;  //EXTERNAL
	output Tile_X0Y1_RES1_O0;  //EXTERNAL
	output Tile_X0Y1_RES1_O1;  //EXTERNAL
	output Tile_X0Y1_RES1_O2;  //EXTERNAL
	output Tile_X0Y1_RES1_O3;  //EXTERNAL
	output Tile_X0Y1_RES2_O0;  //EXTERNAL
	output Tile_X0Y1_RES2_O1;  //EXTERNAL
	output Tile_X0Y1_RES2_O2;  //EXTERNAL
	output Tile_X0Y1_RES2_O3;  //EXTERNAL
	input Tile_X7Y1_OPA_I0;  //EXTERNAL
	input Tile_X7Y1_OPA_I1;  //EXTERNAL
	input Tile_X7Y1_OPA_I2;  //EXTERNAL
	input Tile_X7Y1_OPA_I3;  //EXTERNAL
	input Tile_X7Y1_OPB_I0;  //EXTERNAL
	input Tile_X7Y1_OPB_I1;  //EXTERNAL
	input Tile_X7Y1_OPB_I2;  //EXTERNAL
	input Tile_X7Y1_OPB_I3;  //EXTERNAL
	output Tile_X7Y1_RES0_O0;  //EXTERNAL
	output Tile_X7Y1_RES0_O1;  //EXTERNAL
	output Tile_X7Y1_RES0_O2;  //EXTERNAL
	output Tile_X7Y1_RES0_O3;  //EXTERNAL
	output Tile_X7Y1_RES1_O0;  //EXTERNAL
	output Tile_X7Y1_RES1_O1;  //EXTERNAL
	output Tile_X7Y1_RES1_O2;  //EXTERNAL
	output Tile_X7Y1_RES1_O3;  //EXTERNAL
	output Tile_X7Y1_RES2_O0;  //EXTERNAL
	output Tile_X7Y1_RES2_O1;  //EXTERNAL
	output Tile_X7Y1_RES2_O2;  //EXTERNAL
	output Tile_X7Y1_RES2_O3;  //EXTERNAL
	input Tile_X0Y2_OPA_I0;  //EXTERNAL
	input Tile_X0Y2_OPA_I1;  //EXTERNAL
	input Tile_X0Y2_OPA_I2;  //EXTERNAL
	input Tile_X0Y2_OPA_I3;  //EXTERNAL
	input Tile_X0Y2_OPB_I0;  //EXTERNAL
	input Tile_X0Y2_OPB_I1;  //EXTERNAL
	input Tile_X0Y2_OPB_I2;  //EXTERNAL
	input Tile_X0Y2_OPB_I3;  //EXTERNAL
	output Tile_X0Y2_RES0_O0;  //EXTERNAL
	output Tile_X0Y2_RES0_O1;  //EXTERNAL
	output Tile_X0Y2_RES0_O2;  //EXTERNAL
	output Tile_X0Y2_RES0_O3;  //EXTERNAL
	output Tile_X0Y2_RES1_O0;  //EXTERNAL
	output Tile_X0Y2_RES1_O1;  //EXTERNAL
	output Tile_X0Y2_RES1_O2;  //EXTERNAL
	output Tile_X0Y2_RES1_O3;  //EXTERNAL
	output Tile_X0Y2_RES2_O0;  //EXTERNAL
	output Tile_X0Y2_RES2_O1;  //EXTERNAL
	output Tile_X0Y2_RES2_O2;  //EXTERNAL
	output Tile_X0Y2_RES2_O3;  //EXTERNAL
	input Tile_X7Y2_OPA_I0;  //EXTERNAL
	input Tile_X7Y2_OPA_I1;  //EXTERNAL
	input Tile_X7Y2_OPA_I2;  //EXTERNAL
	input Tile_X7Y2_OPA_I3;  //EXTERNAL
	input Tile_X7Y2_OPB_I0;  //EXTERNAL
	input Tile_X7Y2_OPB_I1;  //EXTERNAL
	input Tile_X7Y2_OPB_I2;  //EXTERNAL
	input Tile_X7Y2_OPB_I3;  //EXTERNAL
	output Tile_X7Y2_RES0_O0;  //EXTERNAL
	output Tile_X7Y2_RES0_O1;  //EXTERNAL
	output Tile_X7Y2_RES0_O2;  //EXTERNAL
	output Tile_X7Y2_RES0_O3;  //EXTERNAL
	output Tile_X7Y2_RES1_O0;  //EXTERNAL
	output Tile_X7Y2_RES1_O1;  //EXTERNAL
	output Tile_X7Y2_RES1_O2;  //EXTERNAL
	output Tile_X7Y2_RES1_O3;  //EXTERNAL
	output Tile_X7Y2_RES2_O0;  //EXTERNAL
	output Tile_X7Y2_RES2_O1;  //EXTERNAL
	output Tile_X7Y2_RES2_O2;  //EXTERNAL
	output Tile_X7Y2_RES2_O3;  //EXTERNAL
	input Tile_X0Y3_OPA_I0;  //EXTERNAL
	input Tile_X0Y3_OPA_I1;  //EXTERNAL
	input Tile_X0Y3_OPA_I2;  //EXTERNAL
	input Tile_X0Y3_OPA_I3;  //EXTERNAL
	input Tile_X0Y3_OPB_I0;  //EXTERNAL
	input Tile_X0Y3_OPB_I1;  //EXTERNAL
	input Tile_X0Y3_OPB_I2;  //EXTERNAL
	input Tile_X0Y3_OPB_I3;  //EXTERNAL
	output Tile_X0Y3_RES0_O0;  //EXTERNAL
	output Tile_X0Y3_RES0_O1;  //EXTERNAL
	output Tile_X0Y3_RES0_O2;  //EXTERNAL
	output Tile_X0Y3_RES0_O3;  //EXTERNAL
	output Tile_X0Y3_RES1_O0;  //EXTERNAL
	output Tile_X0Y3_RES1_O1;  //EXTERNAL
	output Tile_X0Y3_RES1_O2;  //EXTERNAL
	output Tile_X0Y3_RES1_O3;  //EXTERNAL
	output Tile_X0Y3_RES2_O0;  //EXTERNAL
	output Tile_X0Y3_RES2_O1;  //EXTERNAL
	output Tile_X0Y3_RES2_O2;  //EXTERNAL
	output Tile_X0Y3_RES2_O3;  //EXTERNAL
	input Tile_X7Y3_OPA_I0;  //EXTERNAL
	input Tile_X7Y3_OPA_I1;  //EXTERNAL
	input Tile_X7Y3_OPA_I2;  //EXTERNAL
	input Tile_X7Y3_OPA_I3;  //EXTERNAL
	input Tile_X7Y3_OPB_I0;  //EXTERNAL
	input Tile_X7Y3_OPB_I1;  //EXTERNAL
	input Tile_X7Y3_OPB_I2;  //EXTERNAL
	input Tile_X7Y3_OPB_I3;  //EXTERNAL
	output Tile_X7Y3_RES0_O0;  //EXTERNAL
	output Tile_X7Y3_RES0_O1;  //EXTERNAL
	output Tile_X7Y3_RES0_O2;  //EXTERNAL
	output Tile_X7Y3_RES0_O3;  //EXTERNAL
	output Tile_X7Y3_RES1_O0;  //EXTERNAL
	output Tile_X7Y3_RES1_O1;  //EXTERNAL
	output Tile_X7Y3_RES1_O2;  //EXTERNAL
	output Tile_X7Y3_RES1_O3;  //EXTERNAL
	output Tile_X7Y3_RES2_O0;  //EXTERNAL
	output Tile_X7Y3_RES2_O1;  //EXTERNAL
	output Tile_X7Y3_RES2_O2;  //EXTERNAL
	output Tile_X7Y3_RES2_O3;  //EXTERNAL
	input Tile_X0Y4_OPA_I0;  //EXTERNAL
	input Tile_X0Y4_OPA_I1;  //EXTERNAL
	input Tile_X0Y4_OPA_I2;  //EXTERNAL
	input Tile_X0Y4_OPA_I3;  //EXTERNAL
	input Tile_X0Y4_OPB_I0;  //EXTERNAL
	input Tile_X0Y4_OPB_I1;  //EXTERNAL
	input Tile_X0Y4_OPB_I2;  //EXTERNAL
	input Tile_X0Y4_OPB_I3;  //EXTERNAL
	output Tile_X0Y4_RES0_O0;  //EXTERNAL
	output Tile_X0Y4_RES0_O1;  //EXTERNAL
	output Tile_X0Y4_RES0_O2;  //EXTERNAL
	output Tile_X0Y4_RES0_O3;  //EXTERNAL
	output Tile_X0Y4_RES1_O0;  //EXTERNAL
	output Tile_X0Y4_RES1_O1;  //EXTERNAL
	output Tile_X0Y4_RES1_O2;  //EXTERNAL
	output Tile_X0Y4_RES1_O3;  //EXTERNAL
	output Tile_X0Y4_RES2_O0;  //EXTERNAL
	output Tile_X0Y4_RES2_O1;  //EXTERNAL
	output Tile_X0Y4_RES2_O2;  //EXTERNAL
	output Tile_X0Y4_RES2_O3;  //EXTERNAL
	input Tile_X7Y4_OPA_I0;  //EXTERNAL
	input Tile_X7Y4_OPA_I1;  //EXTERNAL
	input Tile_X7Y4_OPA_I2;  //EXTERNAL
	input Tile_X7Y4_OPA_I3;  //EXTERNAL
	input Tile_X7Y4_OPB_I0;  //EXTERNAL
	input Tile_X7Y4_OPB_I1;  //EXTERNAL
	input Tile_X7Y4_OPB_I2;  //EXTERNAL
	input Tile_X7Y4_OPB_I3;  //EXTERNAL
	output Tile_X7Y4_RES0_O0;  //EXTERNAL
	output Tile_X7Y4_RES0_O1;  //EXTERNAL
	output Tile_X7Y4_RES0_O2;  //EXTERNAL
	output Tile_X7Y4_RES0_O3;  //EXTERNAL
	output Tile_X7Y4_RES1_O0;  //EXTERNAL
	output Tile_X7Y4_RES1_O1;  //EXTERNAL
	output Tile_X7Y4_RES1_O2;  //EXTERNAL
	output Tile_X7Y4_RES1_O3;  //EXTERNAL
	output Tile_X7Y4_RES2_O0;  //EXTERNAL
	output Tile_X7Y4_RES2_O1;  //EXTERNAL
	output Tile_X7Y4_RES2_O2;  //EXTERNAL
	output Tile_X7Y4_RES2_O3;  //EXTERNAL
	input Tile_X0Y5_OPA_I0;  //EXTERNAL
	input Tile_X0Y5_OPA_I1;  //EXTERNAL
	input Tile_X0Y5_OPA_I2;  //EXTERNAL
	input Tile_X0Y5_OPA_I3;  //EXTERNAL
	input Tile_X0Y5_OPB_I0;  //EXTERNAL
	input Tile_X0Y5_OPB_I1;  //EXTERNAL
	input Tile_X0Y5_OPB_I2;  //EXTERNAL
	input Tile_X0Y5_OPB_I3;  //EXTERNAL
	output Tile_X0Y5_RES0_O0;  //EXTERNAL
	output Tile_X0Y5_RES0_O1;  //EXTERNAL
	output Tile_X0Y5_RES0_O2;  //EXTERNAL
	output Tile_X0Y5_RES0_O3;  //EXTERNAL
	output Tile_X0Y5_RES1_O0;  //EXTERNAL
	output Tile_X0Y5_RES1_O1;  //EXTERNAL
	output Tile_X0Y5_RES1_O2;  //EXTERNAL
	output Tile_X0Y5_RES1_O3;  //EXTERNAL
	output Tile_X0Y5_RES2_O0;  //EXTERNAL
	output Tile_X0Y5_RES2_O1;  //EXTERNAL
	output Tile_X0Y5_RES2_O2;  //EXTERNAL
	output Tile_X0Y5_RES2_O3;  //EXTERNAL
	input Tile_X7Y5_OPA_I0;  //EXTERNAL
	input Tile_X7Y5_OPA_I1;  //EXTERNAL
	input Tile_X7Y5_OPA_I2;  //EXTERNAL
	input Tile_X7Y5_OPA_I3;  //EXTERNAL
	input Tile_X7Y5_OPB_I0;  //EXTERNAL
	input Tile_X7Y5_OPB_I1;  //EXTERNAL
	input Tile_X7Y5_OPB_I2;  //EXTERNAL
	input Tile_X7Y5_OPB_I3;  //EXTERNAL
	output Tile_X7Y5_RES0_O0;  //EXTERNAL
	output Tile_X7Y5_RES0_O1;  //EXTERNAL
	output Tile_X7Y5_RES0_O2;  //EXTERNAL
	output Tile_X7Y5_RES0_O3;  //EXTERNAL
	output Tile_X7Y5_RES1_O0;  //EXTERNAL
	output Tile_X7Y5_RES1_O1;  //EXTERNAL
	output Tile_X7Y5_RES1_O2;  //EXTERNAL
	output Tile_X7Y5_RES1_O3;  //EXTERNAL
	output Tile_X7Y5_RES2_O0;  //EXTERNAL
	output Tile_X7Y5_RES2_O1;  //EXTERNAL
	output Tile_X7Y5_RES2_O2;  //EXTERNAL
	output Tile_X7Y5_RES2_O3;  //EXTERNAL
	input Tile_X0Y6_OPA_I0;  //EXTERNAL
	input Tile_X0Y6_OPA_I1;  //EXTERNAL
	input Tile_X0Y6_OPA_I2;  //EXTERNAL
	input Tile_X0Y6_OPA_I3;  //EXTERNAL
	input Tile_X0Y6_OPB_I0;  //EXTERNAL
	input Tile_X0Y6_OPB_I1;  //EXTERNAL
	input Tile_X0Y6_OPB_I2;  //EXTERNAL
	input Tile_X0Y6_OPB_I3;  //EXTERNAL
	output Tile_X0Y6_RES0_O0;  //EXTERNAL
	output Tile_X0Y6_RES0_O1;  //EXTERNAL
	output Tile_X0Y6_RES0_O2;  //EXTERNAL
	output Tile_X0Y6_RES0_O3;  //EXTERNAL
	output Tile_X0Y6_RES1_O0;  //EXTERNAL
	output Tile_X0Y6_RES1_O1;  //EXTERNAL
	output Tile_X0Y6_RES1_O2;  //EXTERNAL
	output Tile_X0Y6_RES1_O3;  //EXTERNAL
	output Tile_X0Y6_RES2_O0;  //EXTERNAL
	output Tile_X0Y6_RES2_O1;  //EXTERNAL
	output Tile_X0Y6_RES2_O2;  //EXTERNAL
	output Tile_X0Y6_RES2_O3;  //EXTERNAL
	input Tile_X7Y6_OPA_I0;  //EXTERNAL
	input Tile_X7Y6_OPA_I1;  //EXTERNAL
	input Tile_X7Y6_OPA_I2;  //EXTERNAL
	input Tile_X7Y6_OPA_I3;  //EXTERNAL
	input Tile_X7Y6_OPB_I0;  //EXTERNAL
	input Tile_X7Y6_OPB_I1;  //EXTERNAL
	input Tile_X7Y6_OPB_I2;  //EXTERNAL
	input Tile_X7Y6_OPB_I3;  //EXTERNAL
	output Tile_X7Y6_RES0_O0;  //EXTERNAL
	output Tile_X7Y6_RES0_O1;  //EXTERNAL
	output Tile_X7Y6_RES0_O2;  //EXTERNAL
	output Tile_X7Y6_RES0_O3;  //EXTERNAL
	output Tile_X7Y6_RES1_O0;  //EXTERNAL
	output Tile_X7Y6_RES1_O1;  //EXTERNAL
	output Tile_X7Y6_RES1_O2;  //EXTERNAL
	output Tile_X7Y6_RES1_O3;  //EXTERNAL
	output Tile_X7Y6_RES2_O0;  //EXTERNAL
	output Tile_X7Y6_RES2_O1;  //EXTERNAL
	output Tile_X7Y6_RES2_O2;  //EXTERNAL
	output Tile_X7Y6_RES2_O3;  //EXTERNAL
	input Tile_X0Y7_OPA_I0;  //EXTERNAL
	input Tile_X0Y7_OPA_I1;  //EXTERNAL
	input Tile_X0Y7_OPA_I2;  //EXTERNAL
	input Tile_X0Y7_OPA_I3;  //EXTERNAL
	input Tile_X0Y7_OPB_I0;  //EXTERNAL
	input Tile_X0Y7_OPB_I1;  //EXTERNAL
	input Tile_X0Y7_OPB_I2;  //EXTERNAL
	input Tile_X0Y7_OPB_I3;  //EXTERNAL
	output Tile_X0Y7_RES0_O0;  //EXTERNAL
	output Tile_X0Y7_RES0_O1;  //EXTERNAL
	output Tile_X0Y7_RES0_O2;  //EXTERNAL
	output Tile_X0Y7_RES0_O3;  //EXTERNAL
	output Tile_X0Y7_RES1_O0;  //EXTERNAL
	output Tile_X0Y7_RES1_O1;  //EXTERNAL
	output Tile_X0Y7_RES1_O2;  //EXTERNAL
	output Tile_X0Y7_RES1_O3;  //EXTERNAL
	output Tile_X0Y7_RES2_O0;  //EXTERNAL
	output Tile_X0Y7_RES2_O1;  //EXTERNAL
	output Tile_X0Y7_RES2_O2;  //EXTERNAL
	output Tile_X0Y7_RES2_O3;  //EXTERNAL
	input Tile_X7Y7_OPA_I0;  //EXTERNAL
	input Tile_X7Y7_OPA_I1;  //EXTERNAL
	input Tile_X7Y7_OPA_I2;  //EXTERNAL
	input Tile_X7Y7_OPA_I3;  //EXTERNAL
	input Tile_X7Y7_OPB_I0;  //EXTERNAL
	input Tile_X7Y7_OPB_I1;  //EXTERNAL
	input Tile_X7Y7_OPB_I2;  //EXTERNAL
	input Tile_X7Y7_OPB_I3;  //EXTERNAL
	output Tile_X7Y7_RES0_O0;  //EXTERNAL
	output Tile_X7Y7_RES0_O1;  //EXTERNAL
	output Tile_X7Y7_RES0_O2;  //EXTERNAL
	output Tile_X7Y7_RES0_O3;  //EXTERNAL
	output Tile_X7Y7_RES1_O0;  //EXTERNAL
	output Tile_X7Y7_RES1_O1;  //EXTERNAL
	output Tile_X7Y7_RES1_O2;  //EXTERNAL
	output Tile_X7Y7_RES1_O3;  //EXTERNAL
	output Tile_X7Y7_RES2_O0;  //EXTERNAL
	output Tile_X7Y7_RES2_O1;  //EXTERNAL
	output Tile_X7Y7_RES2_O2;  //EXTERNAL
	output Tile_X7Y7_RES2_O3;  //EXTERNAL
	input Tile_X0Y8_OPA_I0;  //EXTERNAL
	input Tile_X0Y8_OPA_I1;  //EXTERNAL
	input Tile_X0Y8_OPA_I2;  //EXTERNAL
	input Tile_X0Y8_OPA_I3;  //EXTERNAL
	input Tile_X0Y8_OPB_I0;  //EXTERNAL
	input Tile_X0Y8_OPB_I1;  //EXTERNAL
	input Tile_X0Y8_OPB_I2;  //EXTERNAL
	input Tile_X0Y8_OPB_I3;  //EXTERNAL
	output Tile_X0Y8_RES0_O0;  //EXTERNAL
	output Tile_X0Y8_RES0_O1;  //EXTERNAL
	output Tile_X0Y8_RES0_O2;  //EXTERNAL
	output Tile_X0Y8_RES0_O3;  //EXTERNAL
	output Tile_X0Y8_RES1_O0;  //EXTERNAL
	output Tile_X0Y8_RES1_O1;  //EXTERNAL
	output Tile_X0Y8_RES1_O2;  //EXTERNAL
	output Tile_X0Y8_RES1_O3;  //EXTERNAL
	output Tile_X0Y8_RES2_O0;  //EXTERNAL
	output Tile_X0Y8_RES2_O1;  //EXTERNAL
	output Tile_X0Y8_RES2_O2;  //EXTERNAL
	output Tile_X0Y8_RES2_O3;  //EXTERNAL
	input Tile_X7Y8_OPA_I0;  //EXTERNAL
	input Tile_X7Y8_OPA_I1;  //EXTERNAL
	input Tile_X7Y8_OPA_I2;  //EXTERNAL
	input Tile_X7Y8_OPA_I3;  //EXTERNAL
	input Tile_X7Y8_OPB_I0;  //EXTERNAL
	input Tile_X7Y8_OPB_I1;  //EXTERNAL
	input Tile_X7Y8_OPB_I2;  //EXTERNAL
	input Tile_X7Y8_OPB_I3;  //EXTERNAL
	output Tile_X7Y8_RES0_O0;  //EXTERNAL
	output Tile_X7Y8_RES0_O1;  //EXTERNAL
	output Tile_X7Y8_RES0_O2;  //EXTERNAL
	output Tile_X7Y8_RES0_O3;  //EXTERNAL
	output Tile_X7Y8_RES1_O0;  //EXTERNAL
	output Tile_X7Y8_RES1_O1;  //EXTERNAL
	output Tile_X7Y8_RES1_O2;  //EXTERNAL
	output Tile_X7Y8_RES1_O3;  //EXTERNAL
	output Tile_X7Y8_RES2_O0;  //EXTERNAL
	output Tile_X7Y8_RES2_O1;  //EXTERNAL
	output Tile_X7Y8_RES2_O2;  //EXTERNAL
	output Tile_X7Y8_RES2_O3;  //EXTERNAL
	input Tile_X0Y9_OPA_I0;  //EXTERNAL
	input Tile_X0Y9_OPA_I1;  //EXTERNAL
	input Tile_X0Y9_OPA_I2;  //EXTERNAL
	input Tile_X0Y9_OPA_I3;  //EXTERNAL
	input Tile_X0Y9_OPB_I0;  //EXTERNAL
	input Tile_X0Y9_OPB_I1;  //EXTERNAL
	input Tile_X0Y9_OPB_I2;  //EXTERNAL
	input Tile_X0Y9_OPB_I3;  //EXTERNAL
	output Tile_X0Y9_RES0_O0;  //EXTERNAL
	output Tile_X0Y9_RES0_O1;  //EXTERNAL
	output Tile_X0Y9_RES0_O2;  //EXTERNAL
	output Tile_X0Y9_RES0_O3;  //EXTERNAL
	output Tile_X0Y9_RES1_O0;  //EXTERNAL
	output Tile_X0Y9_RES1_O1;  //EXTERNAL
	output Tile_X0Y9_RES1_O2;  //EXTERNAL
	output Tile_X0Y9_RES1_O3;  //EXTERNAL
	output Tile_X0Y9_RES2_O0;  //EXTERNAL
	output Tile_X0Y9_RES2_O1;  //EXTERNAL
	output Tile_X0Y9_RES2_O2;  //EXTERNAL
	output Tile_X0Y9_RES2_O3;  //EXTERNAL
	input Tile_X7Y9_OPA_I0;  //EXTERNAL
	input Tile_X7Y9_OPA_I1;  //EXTERNAL
	input Tile_X7Y9_OPA_I2;  //EXTERNAL
	input Tile_X7Y9_OPA_I3;  //EXTERNAL
	input Tile_X7Y9_OPB_I0;  //EXTERNAL
	input Tile_X7Y9_OPB_I1;  //EXTERNAL
	input Tile_X7Y9_OPB_I2;  //EXTERNAL
	input Tile_X7Y9_OPB_I3;  //EXTERNAL
	output Tile_X7Y9_RES0_O0;  //EXTERNAL
	output Tile_X7Y9_RES0_O1;  //EXTERNAL
	output Tile_X7Y9_RES0_O2;  //EXTERNAL
	output Tile_X7Y9_RES0_O3;  //EXTERNAL
	output Tile_X7Y9_RES1_O0;  //EXTERNAL
	output Tile_X7Y9_RES1_O1;  //EXTERNAL
	output Tile_X7Y9_RES1_O2;  //EXTERNAL
	output Tile_X7Y9_RES1_O3;  //EXTERNAL
	output Tile_X7Y9_RES2_O0;  //EXTERNAL
	output Tile_X7Y9_RES2_O1;  //EXTERNAL
	output Tile_X7Y9_RES2_O2;  //EXTERNAL
	output Tile_X7Y9_RES2_O3;  //EXTERNAL
	input Tile_X0Y10_OPA_I0;  //EXTERNAL
	input Tile_X0Y10_OPA_I1;  //EXTERNAL
	input Tile_X0Y10_OPA_I2;  //EXTERNAL
	input Tile_X0Y10_OPA_I3;  //EXTERNAL
	input Tile_X0Y10_OPB_I0;  //EXTERNAL
	input Tile_X0Y10_OPB_I1;  //EXTERNAL
	input Tile_X0Y10_OPB_I2;  //EXTERNAL
	input Tile_X0Y10_OPB_I3;  //EXTERNAL
	output Tile_X0Y10_RES0_O0;  //EXTERNAL
	output Tile_X0Y10_RES0_O1;  //EXTERNAL
	output Tile_X0Y10_RES0_O2;  //EXTERNAL
	output Tile_X0Y10_RES0_O3;  //EXTERNAL
	output Tile_X0Y10_RES1_O0;  //EXTERNAL
	output Tile_X0Y10_RES1_O1;  //EXTERNAL
	output Tile_X0Y10_RES1_O2;  //EXTERNAL
	output Tile_X0Y10_RES1_O3;  //EXTERNAL
	output Tile_X0Y10_RES2_O0;  //EXTERNAL
	output Tile_X0Y10_RES2_O1;  //EXTERNAL
	output Tile_X0Y10_RES2_O2;  //EXTERNAL
	output Tile_X0Y10_RES2_O3;  //EXTERNAL
	input Tile_X7Y10_OPA_I0;  //EXTERNAL
	input Tile_X7Y10_OPA_I1;  //EXTERNAL
	input Tile_X7Y10_OPA_I2;  //EXTERNAL
	input Tile_X7Y10_OPA_I3;  //EXTERNAL
	input Tile_X7Y10_OPB_I0;  //EXTERNAL
	input Tile_X7Y10_OPB_I1;  //EXTERNAL
	input Tile_X7Y10_OPB_I2;  //EXTERNAL
	input Tile_X7Y10_OPB_I3;  //EXTERNAL
	output Tile_X7Y10_RES0_O0;  //EXTERNAL
	output Tile_X7Y10_RES0_O1;  //EXTERNAL
	output Tile_X7Y10_RES0_O2;  //EXTERNAL
	output Tile_X7Y10_RES0_O3;  //EXTERNAL
	output Tile_X7Y10_RES1_O0;  //EXTERNAL
	output Tile_X7Y10_RES1_O1;  //EXTERNAL
	output Tile_X7Y10_RES1_O2;  //EXTERNAL
	output Tile_X7Y10_RES1_O3;  //EXTERNAL
	output Tile_X7Y10_RES2_O0;  //EXTERNAL
	output Tile_X7Y10_RES2_O1;  //EXTERNAL
	output Tile_X7Y10_RES2_O2;  //EXTERNAL
	output Tile_X7Y10_RES2_O3;  //EXTERNAL
	input [(FrameBitsPerRow*12)-1:0] FrameData;   // CONFIG_PORT this is a keyword needed to connect the tile to the bitstream frame register
	input [(MaxFramesPerCol*8)-1:0] FrameStrobe;   // CONFIG_PORT this is a keyword needed to connect the tile to the bitstream frame register 
	//global


//signal declarations
//configuration signal declarations

	wire [FrameBitsPerRow-1:0] Tile_Y0_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y1_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y2_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y3_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y4_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y5_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y6_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y7_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y8_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y9_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y10_FrameData;
	wire [FrameBitsPerRow-1:0] Tile_Y11_FrameData;
	wire [MaxFramesPerCol-1:0] Tile_X0_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X1_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X2_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X3_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X4_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X5_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X6_FrameStrobe;
	wire [MaxFramesPerCol-1:0] Tile_X7_FrameStrobe;
	wire [FrameBitsPerRow-1:0] Tile_X0Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y0_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y1_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y2_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y3_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y4_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y5_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y6_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y7_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y8_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y9_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y10_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X0Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X1Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X2Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X3Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X4Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X5Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X6Y11_FrameData_O;
	wire [FrameBitsPerRow-1:0] Tile_X7Y11_FrameData_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y0_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y1_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y2_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y3_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y4_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y5_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y6_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y7_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y8_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y9_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y10_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X0Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X1Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X2Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X3Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X4Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X5Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X6Y11_FrameStrobe_O;
	wire [MaxFramesPerCol-1:0] Tile_X7Y11_FrameStrobe_O;

//tile-to-tile signal declarations

	wire [3:0] Tile_X1Y0_S1BEG;
	wire [7:0] Tile_X1Y0_S2BEG;
	wire [7:0] Tile_X1Y0_S2BEGb;
	wire [15:0] Tile_X1Y0_S4BEG;
	wire [15:0] Tile_X1Y0_SS4BEG;
	wire [3:0] Tile_X2Y0_S1BEG;
	wire [7:0] Tile_X2Y0_S2BEG;
	wire [7:0] Tile_X2Y0_S2BEGb;
	wire [15:0] Tile_X2Y0_S4BEG;
	wire [15:0] Tile_X2Y0_SS4BEG;
	wire [3:0] Tile_X3Y0_S1BEG;
	wire [7:0] Tile_X3Y0_S2BEG;
	wire [7:0] Tile_X3Y0_S2BEGb;
	wire [15:0] Tile_X3Y0_S4BEG;
	wire [15:0] Tile_X3Y0_SS4BEG;
	wire [3:0] Tile_X4Y0_S1BEG;
	wire [7:0] Tile_X4Y0_S2BEG;
	wire [7:0] Tile_X4Y0_S2BEGb;
	wire [15:0] Tile_X4Y0_S4BEG;
	wire [15:0] Tile_X4Y0_SS4BEG;
	wire [3:0] Tile_X5Y0_S1BEG;
	wire [7:0] Tile_X5Y0_S2BEG;
	wire [7:0] Tile_X5Y0_S2BEGb;
	wire [15:0] Tile_X5Y0_S4BEG;
	wire [15:0] Tile_X5Y0_SS4BEG;
	wire [3:0] Tile_X6Y0_S1BEG;
	wire [7:0] Tile_X6Y0_S2BEG;
	wire [7:0] Tile_X6Y0_S2BEGb;
	wire [15:0] Tile_X6Y0_S4BEG;
	wire [15:0] Tile_X6Y0_SS4BEG;
	wire [3:0] Tile_X0Y1_E1BEG;
	wire [7:0] Tile_X0Y1_E2BEG;
	wire [7:0] Tile_X0Y1_E2BEGb;
	wire [15:0] Tile_X0Y1_EE4BEG;
	wire [11:0] Tile_X0Y1_E6BEG;
	wire [3:0] Tile_X1Y1_N1BEG;
	wire [7:0] Tile_X1Y1_N2BEG;
	wire [7:0] Tile_X1Y1_N2BEGb;
	wire [15:0] Tile_X1Y1_N4BEG;
	wire [15:0] Tile_X1Y1_NN4BEG;
	wire [3:0] Tile_X1Y1_E1BEG;
	wire [7:0] Tile_X1Y1_E2BEG;
	wire [7:0] Tile_X1Y1_E2BEGb;
	wire [15:0] Tile_X1Y1_EE4BEG;
	wire [11:0] Tile_X1Y1_E6BEG;
	wire [3:0] Tile_X1Y1_S1BEG;
	wire [7:0] Tile_X1Y1_S2BEG;
	wire [7:0] Tile_X1Y1_S2BEGb;
	wire [15:0] Tile_X1Y1_S4BEG;
	wire [15:0] Tile_X1Y1_SS4BEG;
	wire [17:0] Tile_X1Y1_top2bot;
	wire [3:0] Tile_X1Y1_W1BEG;
	wire [7:0] Tile_X1Y1_W2BEG;
	wire [7:0] Tile_X1Y1_W2BEGb;
	wire [15:0] Tile_X1Y1_WW4BEG;
	wire [11:0] Tile_X1Y1_W6BEG;
	wire [3:0] Tile_X2Y1_N1BEG;
	wire [7:0] Tile_X2Y1_N2BEG;
	wire [7:0] Tile_X2Y1_N2BEGb;
	wire [15:0] Tile_X2Y1_N4BEG;
	wire [15:0] Tile_X2Y1_NN4BEG;
	wire [0:0] Tile_X2Y1_Co;
	wire [3:0] Tile_X2Y1_E1BEG;
	wire [7:0] Tile_X2Y1_E2BEG;
	wire [7:0] Tile_X2Y1_E2BEGb;
	wire [15:0] Tile_X2Y1_EE4BEG;
	wire [11:0] Tile_X2Y1_E6BEG;
	wire [3:0] Tile_X2Y1_S1BEG;
	wire [7:0] Tile_X2Y1_S2BEG;
	wire [7:0] Tile_X2Y1_S2BEGb;
	wire [15:0] Tile_X2Y1_S4BEG;
	wire [15:0] Tile_X2Y1_SS4BEG;
	wire [3:0] Tile_X2Y1_W1BEG;
	wire [7:0] Tile_X2Y1_W2BEG;
	wire [7:0] Tile_X2Y1_W2BEGb;
	wire [15:0] Tile_X2Y1_WW4BEG;
	wire [11:0] Tile_X2Y1_W6BEG;
	wire [3:0] Tile_X3Y1_N1BEG;
	wire [7:0] Tile_X3Y1_N2BEG;
	wire [7:0] Tile_X3Y1_N2BEGb;
	wire [15:0] Tile_X3Y1_N4BEG;
	wire [15:0] Tile_X3Y1_NN4BEG;
	wire [0:0] Tile_X3Y1_Co;
	wire [3:0] Tile_X3Y1_E1BEG;
	wire [7:0] Tile_X3Y1_E2BEG;
	wire [7:0] Tile_X3Y1_E2BEGb;
	wire [15:0] Tile_X3Y1_EE4BEG;
	wire [11:0] Tile_X3Y1_E6BEG;
	wire [3:0] Tile_X3Y1_S1BEG;
	wire [7:0] Tile_X3Y1_S2BEG;
	wire [7:0] Tile_X3Y1_S2BEGb;
	wire [15:0] Tile_X3Y1_S4BEG;
	wire [15:0] Tile_X3Y1_SS4BEG;
	wire [3:0] Tile_X3Y1_W1BEG;
	wire [7:0] Tile_X3Y1_W2BEG;
	wire [7:0] Tile_X3Y1_W2BEGb;
	wire [15:0] Tile_X3Y1_WW4BEG;
	wire [11:0] Tile_X3Y1_W6BEG;
	wire [3:0] Tile_X4Y1_N1BEG;
	wire [7:0] Tile_X4Y1_N2BEG;
	wire [7:0] Tile_X4Y1_N2BEGb;
	wire [15:0] Tile_X4Y1_N4BEG;
	wire [15:0] Tile_X4Y1_NN4BEG;
	wire [0:0] Tile_X4Y1_Co;
	wire [3:0] Tile_X4Y1_E1BEG;
	wire [7:0] Tile_X4Y1_E2BEG;
	wire [7:0] Tile_X4Y1_E2BEGb;
	wire [15:0] Tile_X4Y1_EE4BEG;
	wire [11:0] Tile_X4Y1_E6BEG;
	wire [3:0] Tile_X4Y1_S1BEG;
	wire [7:0] Tile_X4Y1_S2BEG;
	wire [7:0] Tile_X4Y1_S2BEGb;
	wire [15:0] Tile_X4Y1_S4BEG;
	wire [15:0] Tile_X4Y1_SS4BEG;
	wire [3:0] Tile_X4Y1_W1BEG;
	wire [7:0] Tile_X4Y1_W2BEG;
	wire [7:0] Tile_X4Y1_W2BEGb;
	wire [15:0] Tile_X4Y1_WW4BEG;
	wire [11:0] Tile_X4Y1_W6BEG;
	wire [3:0] Tile_X5Y1_N1BEG;
	wire [7:0] Tile_X5Y1_N2BEG;
	wire [7:0] Tile_X5Y1_N2BEGb;
	wire [15:0] Tile_X5Y1_N4BEG;
	wire [15:0] Tile_X5Y1_NN4BEG;
	wire [3:0] Tile_X5Y1_E1BEG;
	wire [7:0] Tile_X5Y1_E2BEG;
	wire [7:0] Tile_X5Y1_E2BEGb;
	wire [15:0] Tile_X5Y1_EE4BEG;
	wire [11:0] Tile_X5Y1_E6BEG;
	wire [3:0] Tile_X5Y1_S1BEG;
	wire [7:0] Tile_X5Y1_S2BEG;
	wire [7:0] Tile_X5Y1_S2BEGb;
	wire [15:0] Tile_X5Y1_S4BEG;
	wire [15:0] Tile_X5Y1_SS4BEG;
	wire [17:0] Tile_X5Y1_top2bot;
	wire [3:0] Tile_X5Y1_W1BEG;
	wire [7:0] Tile_X5Y1_W2BEG;
	wire [7:0] Tile_X5Y1_W2BEGb;
	wire [15:0] Tile_X5Y1_WW4BEG;
	wire [11:0] Tile_X5Y1_W6BEG;
	wire [3:0] Tile_X6Y1_N1BEG;
	wire [7:0] Tile_X6Y1_N2BEG;
	wire [7:0] Tile_X6Y1_N2BEGb;
	wire [15:0] Tile_X6Y1_N4BEG;
	wire [15:0] Tile_X6Y1_NN4BEG;
	wire [0:0] Tile_X6Y1_Co;
	wire [3:0] Tile_X6Y1_E1BEG;
	wire [7:0] Tile_X6Y1_E2BEG;
	wire [7:0] Tile_X6Y1_E2BEGb;
	wire [15:0] Tile_X6Y1_EE4BEG;
	wire [11:0] Tile_X6Y1_E6BEG;
	wire [3:0] Tile_X6Y1_S1BEG;
	wire [7:0] Tile_X6Y1_S2BEG;
	wire [7:0] Tile_X6Y1_S2BEGb;
	wire [15:0] Tile_X6Y1_S4BEG;
	wire [15:0] Tile_X6Y1_SS4BEG;
	wire [3:0] Tile_X6Y1_W1BEG;
	wire [7:0] Tile_X6Y1_W2BEG;
	wire [7:0] Tile_X6Y1_W2BEGb;
	wire [15:0] Tile_X6Y1_WW4BEG;
	wire [11:0] Tile_X6Y1_W6BEG;
	wire [3:0] Tile_X7Y1_W1BEG;
	wire [7:0] Tile_X7Y1_W2BEG;
	wire [7:0] Tile_X7Y1_W2BEGb;
	wire [15:0] Tile_X7Y1_WW4BEG;
	wire [11:0] Tile_X7Y1_W6BEG;
	wire [3:0] Tile_X0Y2_E1BEG;
	wire [7:0] Tile_X0Y2_E2BEG;
	wire [7:0] Tile_X0Y2_E2BEGb;
	wire [15:0] Tile_X0Y2_EE4BEG;
	wire [11:0] Tile_X0Y2_E6BEG;
	wire [3:0] Tile_X1Y2_N1BEG;
	wire [7:0] Tile_X1Y2_N2BEG;
	wire [7:0] Tile_X1Y2_N2BEGb;
	wire [15:0] Tile_X1Y2_N4BEG;
	wire [15:0] Tile_X1Y2_NN4BEG;
	wire [9:0] Tile_X1Y2_bot2top;
	wire [3:0] Tile_X1Y2_E1BEG;
	wire [7:0] Tile_X1Y2_E2BEG;
	wire [7:0] Tile_X1Y2_E2BEGb;
	wire [15:0] Tile_X1Y2_EE4BEG;
	wire [11:0] Tile_X1Y2_E6BEG;
	wire [3:0] Tile_X1Y2_S1BEG;
	wire [7:0] Tile_X1Y2_S2BEG;
	wire [7:0] Tile_X1Y2_S2BEGb;
	wire [15:0] Tile_X1Y2_S4BEG;
	wire [15:0] Tile_X1Y2_SS4BEG;
	wire [3:0] Tile_X1Y2_W1BEG;
	wire [7:0] Tile_X1Y2_W2BEG;
	wire [7:0] Tile_X1Y2_W2BEGb;
	wire [15:0] Tile_X1Y2_WW4BEG;
	wire [11:0] Tile_X1Y2_W6BEG;
	wire [3:0] Tile_X2Y2_N1BEG;
	wire [7:0] Tile_X2Y2_N2BEG;
	wire [7:0] Tile_X2Y2_N2BEGb;
	wire [15:0] Tile_X2Y2_N4BEG;
	wire [15:0] Tile_X2Y2_NN4BEG;
	wire [0:0] Tile_X2Y2_Co;
	wire [3:0] Tile_X2Y2_E1BEG;
	wire [7:0] Tile_X2Y2_E2BEG;
	wire [7:0] Tile_X2Y2_E2BEGb;
	wire [15:0] Tile_X2Y2_EE4BEG;
	wire [11:0] Tile_X2Y2_E6BEG;
	wire [3:0] Tile_X2Y2_S1BEG;
	wire [7:0] Tile_X2Y2_S2BEG;
	wire [7:0] Tile_X2Y2_S2BEGb;
	wire [15:0] Tile_X2Y2_S4BEG;
	wire [15:0] Tile_X2Y2_SS4BEG;
	wire [3:0] Tile_X2Y2_W1BEG;
	wire [7:0] Tile_X2Y2_W2BEG;
	wire [7:0] Tile_X2Y2_W2BEGb;
	wire [15:0] Tile_X2Y2_WW4BEG;
	wire [11:0] Tile_X2Y2_W6BEG;
	wire [3:0] Tile_X3Y2_N1BEG;
	wire [7:0] Tile_X3Y2_N2BEG;
	wire [7:0] Tile_X3Y2_N2BEGb;
	wire [15:0] Tile_X3Y2_N4BEG;
	wire [15:0] Tile_X3Y2_NN4BEG;
	wire [0:0] Tile_X3Y2_Co;
	wire [3:0] Tile_X3Y2_E1BEG;
	wire [7:0] Tile_X3Y2_E2BEG;
	wire [7:0] Tile_X3Y2_E2BEGb;
	wire [15:0] Tile_X3Y2_EE4BEG;
	wire [11:0] Tile_X3Y2_E6BEG;
	wire [3:0] Tile_X3Y2_S1BEG;
	wire [7:0] Tile_X3Y2_S2BEG;
	wire [7:0] Tile_X3Y2_S2BEGb;
	wire [15:0] Tile_X3Y2_S4BEG;
	wire [15:0] Tile_X3Y2_SS4BEG;
	wire [3:0] Tile_X3Y2_W1BEG;
	wire [7:0] Tile_X3Y2_W2BEG;
	wire [7:0] Tile_X3Y2_W2BEGb;
	wire [15:0] Tile_X3Y2_WW4BEG;
	wire [11:0] Tile_X3Y2_W6BEG;
	wire [3:0] Tile_X4Y2_N1BEG;
	wire [7:0] Tile_X4Y2_N2BEG;
	wire [7:0] Tile_X4Y2_N2BEGb;
	wire [15:0] Tile_X4Y2_N4BEG;
	wire [15:0] Tile_X4Y2_NN4BEG;
	wire [0:0] Tile_X4Y2_Co;
	wire [3:0] Tile_X4Y2_E1BEG;
	wire [7:0] Tile_X4Y2_E2BEG;
	wire [7:0] Tile_X4Y2_E2BEGb;
	wire [15:0] Tile_X4Y2_EE4BEG;
	wire [11:0] Tile_X4Y2_E6BEG;
	wire [3:0] Tile_X4Y2_S1BEG;
	wire [7:0] Tile_X4Y2_S2BEG;
	wire [7:0] Tile_X4Y2_S2BEGb;
	wire [15:0] Tile_X4Y2_S4BEG;
	wire [15:0] Tile_X4Y2_SS4BEG;
	wire [3:0] Tile_X4Y2_W1BEG;
	wire [7:0] Tile_X4Y2_W2BEG;
	wire [7:0] Tile_X4Y2_W2BEGb;
	wire [15:0] Tile_X4Y2_WW4BEG;
	wire [11:0] Tile_X4Y2_W6BEG;
	wire [3:0] Tile_X5Y2_N1BEG;
	wire [7:0] Tile_X5Y2_N2BEG;
	wire [7:0] Tile_X5Y2_N2BEGb;
	wire [15:0] Tile_X5Y2_N4BEG;
	wire [15:0] Tile_X5Y2_NN4BEG;
	wire [9:0] Tile_X5Y2_bot2top;
	wire [3:0] Tile_X5Y2_E1BEG;
	wire [7:0] Tile_X5Y2_E2BEG;
	wire [7:0] Tile_X5Y2_E2BEGb;
	wire [15:0] Tile_X5Y2_EE4BEG;
	wire [11:0] Tile_X5Y2_E6BEG;
	wire [3:0] Tile_X5Y2_S1BEG;
	wire [7:0] Tile_X5Y2_S2BEG;
	wire [7:0] Tile_X5Y2_S2BEGb;
	wire [15:0] Tile_X5Y2_S4BEG;
	wire [15:0] Tile_X5Y2_SS4BEG;
	wire [3:0] Tile_X5Y2_W1BEG;
	wire [7:0] Tile_X5Y2_W2BEG;
	wire [7:0] Tile_X5Y2_W2BEGb;
	wire [15:0] Tile_X5Y2_WW4BEG;
	wire [11:0] Tile_X5Y2_W6BEG;
	wire [3:0] Tile_X6Y2_N1BEG;
	wire [7:0] Tile_X6Y2_N2BEG;
	wire [7:0] Tile_X6Y2_N2BEGb;
	wire [15:0] Tile_X6Y2_N4BEG;
	wire [15:0] Tile_X6Y2_NN4BEG;
	wire [0:0] Tile_X6Y2_Co;
	wire [3:0] Tile_X6Y2_E1BEG;
	wire [7:0] Tile_X6Y2_E2BEG;
	wire [7:0] Tile_X6Y2_E2BEGb;
	wire [15:0] Tile_X6Y2_EE4BEG;
	wire [11:0] Tile_X6Y2_E6BEG;
	wire [3:0] Tile_X6Y2_S1BEG;
	wire [7:0] Tile_X6Y2_S2BEG;
	wire [7:0] Tile_X6Y2_S2BEGb;
	wire [15:0] Tile_X6Y2_S4BEG;
	wire [15:0] Tile_X6Y2_SS4BEG;
	wire [3:0] Tile_X6Y2_W1BEG;
	wire [7:0] Tile_X6Y2_W2BEG;
	wire [7:0] Tile_X6Y2_W2BEGb;
	wire [15:0] Tile_X6Y2_WW4BEG;
	wire [11:0] Tile_X6Y2_W6BEG;
	wire [3:0] Tile_X7Y2_W1BEG;
	wire [7:0] Tile_X7Y2_W2BEG;
	wire [7:0] Tile_X7Y2_W2BEGb;
	wire [15:0] Tile_X7Y2_WW4BEG;
	wire [11:0] Tile_X7Y2_W6BEG;
	wire [3:0] Tile_X0Y3_E1BEG;
	wire [7:0] Tile_X0Y3_E2BEG;
	wire [7:0] Tile_X0Y3_E2BEGb;
	wire [15:0] Tile_X0Y3_EE4BEG;
	wire [11:0] Tile_X0Y3_E6BEG;
	wire [3:0] Tile_X1Y3_N1BEG;
	wire [7:0] Tile_X1Y3_N2BEG;
	wire [7:0] Tile_X1Y3_N2BEGb;
	wire [15:0] Tile_X1Y3_N4BEG;
	wire [15:0] Tile_X1Y3_NN4BEG;
	wire [3:0] Tile_X1Y3_E1BEG;
	wire [7:0] Tile_X1Y3_E2BEG;
	wire [7:0] Tile_X1Y3_E2BEGb;
	wire [15:0] Tile_X1Y3_EE4BEG;
	wire [11:0] Tile_X1Y3_E6BEG;
	wire [3:0] Tile_X1Y3_S1BEG;
	wire [7:0] Tile_X1Y3_S2BEG;
	wire [7:0] Tile_X1Y3_S2BEGb;
	wire [15:0] Tile_X1Y3_S4BEG;
	wire [15:0] Tile_X1Y3_SS4BEG;
	wire [17:0] Tile_X1Y3_top2bot;
	wire [3:0] Tile_X1Y3_W1BEG;
	wire [7:0] Tile_X1Y3_W2BEG;
	wire [7:0] Tile_X1Y3_W2BEGb;
	wire [15:0] Tile_X1Y3_WW4BEG;
	wire [11:0] Tile_X1Y3_W6BEG;
	wire [3:0] Tile_X2Y3_N1BEG;
	wire [7:0] Tile_X2Y3_N2BEG;
	wire [7:0] Tile_X2Y3_N2BEGb;
	wire [15:0] Tile_X2Y3_N4BEG;
	wire [15:0] Tile_X2Y3_NN4BEG;
	wire [0:0] Tile_X2Y3_Co;
	wire [3:0] Tile_X2Y3_E1BEG;
	wire [7:0] Tile_X2Y3_E2BEG;
	wire [7:0] Tile_X2Y3_E2BEGb;
	wire [15:0] Tile_X2Y3_EE4BEG;
	wire [11:0] Tile_X2Y3_E6BEG;
	wire [3:0] Tile_X2Y3_S1BEG;
	wire [7:0] Tile_X2Y3_S2BEG;
	wire [7:0] Tile_X2Y3_S2BEGb;
	wire [15:0] Tile_X2Y3_S4BEG;
	wire [15:0] Tile_X2Y3_SS4BEG;
	wire [3:0] Tile_X2Y3_W1BEG;
	wire [7:0] Tile_X2Y3_W2BEG;
	wire [7:0] Tile_X2Y3_W2BEGb;
	wire [15:0] Tile_X2Y3_WW4BEG;
	wire [11:0] Tile_X2Y3_W6BEG;
	wire [3:0] Tile_X3Y3_N1BEG;
	wire [7:0] Tile_X3Y3_N2BEG;
	wire [7:0] Tile_X3Y3_N2BEGb;
	wire [15:0] Tile_X3Y3_N4BEG;
	wire [15:0] Tile_X3Y3_NN4BEG;
	wire [0:0] Tile_X3Y3_Co;
	wire [3:0] Tile_X3Y3_E1BEG;
	wire [7:0] Tile_X3Y3_E2BEG;
	wire [7:0] Tile_X3Y3_E2BEGb;
	wire [15:0] Tile_X3Y3_EE4BEG;
	wire [11:0] Tile_X3Y3_E6BEG;
	wire [3:0] Tile_X3Y3_S1BEG;
	wire [7:0] Tile_X3Y3_S2BEG;
	wire [7:0] Tile_X3Y3_S2BEGb;
	wire [15:0] Tile_X3Y3_S4BEG;
	wire [15:0] Tile_X3Y3_SS4BEG;
	wire [3:0] Tile_X3Y3_W1BEG;
	wire [7:0] Tile_X3Y3_W2BEG;
	wire [7:0] Tile_X3Y3_W2BEGb;
	wire [15:0] Tile_X3Y3_WW4BEG;
	wire [11:0] Tile_X3Y3_W6BEG;
	wire [3:0] Tile_X4Y3_N1BEG;
	wire [7:0] Tile_X4Y3_N2BEG;
	wire [7:0] Tile_X4Y3_N2BEGb;
	wire [15:0] Tile_X4Y3_N4BEG;
	wire [15:0] Tile_X4Y3_NN4BEG;
	wire [0:0] Tile_X4Y3_Co;
	wire [3:0] Tile_X4Y3_E1BEG;
	wire [7:0] Tile_X4Y3_E2BEG;
	wire [7:0] Tile_X4Y3_E2BEGb;
	wire [15:0] Tile_X4Y3_EE4BEG;
	wire [11:0] Tile_X4Y3_E6BEG;
	wire [3:0] Tile_X4Y3_S1BEG;
	wire [7:0] Tile_X4Y3_S2BEG;
	wire [7:0] Tile_X4Y3_S2BEGb;
	wire [15:0] Tile_X4Y3_S4BEG;
	wire [15:0] Tile_X4Y3_SS4BEG;
	wire [3:0] Tile_X4Y3_W1BEG;
	wire [7:0] Tile_X4Y3_W2BEG;
	wire [7:0] Tile_X4Y3_W2BEGb;
	wire [15:0] Tile_X4Y3_WW4BEG;
	wire [11:0] Tile_X4Y3_W6BEG;
	wire [3:0] Tile_X5Y3_N1BEG;
	wire [7:0] Tile_X5Y3_N2BEG;
	wire [7:0] Tile_X5Y3_N2BEGb;
	wire [15:0] Tile_X5Y3_N4BEG;
	wire [15:0] Tile_X5Y3_NN4BEG;
	wire [3:0] Tile_X5Y3_E1BEG;
	wire [7:0] Tile_X5Y3_E2BEG;
	wire [7:0] Tile_X5Y3_E2BEGb;
	wire [15:0] Tile_X5Y3_EE4BEG;
	wire [11:0] Tile_X5Y3_E6BEG;
	wire [3:0] Tile_X5Y3_S1BEG;
	wire [7:0] Tile_X5Y3_S2BEG;
	wire [7:0] Tile_X5Y3_S2BEGb;
	wire [15:0] Tile_X5Y3_S4BEG;
	wire [15:0] Tile_X5Y3_SS4BEG;
	wire [17:0] Tile_X5Y3_top2bot;
	wire [3:0] Tile_X5Y3_W1BEG;
	wire [7:0] Tile_X5Y3_W2BEG;
	wire [7:0] Tile_X5Y3_W2BEGb;
	wire [15:0] Tile_X5Y3_WW4BEG;
	wire [11:0] Tile_X5Y3_W6BEG;
	wire [3:0] Tile_X6Y3_N1BEG;
	wire [7:0] Tile_X6Y3_N2BEG;
	wire [7:0] Tile_X6Y3_N2BEGb;
	wire [15:0] Tile_X6Y3_N4BEG;
	wire [15:0] Tile_X6Y3_NN4BEG;
	wire [0:0] Tile_X6Y3_Co;
	wire [3:0] Tile_X6Y3_E1BEG;
	wire [7:0] Tile_X6Y3_E2BEG;
	wire [7:0] Tile_X6Y3_E2BEGb;
	wire [15:0] Tile_X6Y3_EE4BEG;
	wire [11:0] Tile_X6Y3_E6BEG;
	wire [3:0] Tile_X6Y3_S1BEG;
	wire [7:0] Tile_X6Y3_S2BEG;
	wire [7:0] Tile_X6Y3_S2BEGb;
	wire [15:0] Tile_X6Y3_S4BEG;
	wire [15:0] Tile_X6Y3_SS4BEG;
	wire [3:0] Tile_X6Y3_W1BEG;
	wire [7:0] Tile_X6Y3_W2BEG;
	wire [7:0] Tile_X6Y3_W2BEGb;
	wire [15:0] Tile_X6Y3_WW4BEG;
	wire [11:0] Tile_X6Y3_W6BEG;
	wire [3:0] Tile_X7Y3_W1BEG;
	wire [7:0] Tile_X7Y3_W2BEG;
	wire [7:0] Tile_X7Y3_W2BEGb;
	wire [15:0] Tile_X7Y3_WW4BEG;
	wire [11:0] Tile_X7Y3_W6BEG;
	wire [3:0] Tile_X0Y4_E1BEG;
	wire [7:0] Tile_X0Y4_E2BEG;
	wire [7:0] Tile_X0Y4_E2BEGb;
	wire [15:0] Tile_X0Y4_EE4BEG;
	wire [11:0] Tile_X0Y4_E6BEG;
	wire [3:0] Tile_X1Y4_N1BEG;
	wire [7:0] Tile_X1Y4_N2BEG;
	wire [7:0] Tile_X1Y4_N2BEGb;
	wire [15:0] Tile_X1Y4_N4BEG;
	wire [15:0] Tile_X1Y4_NN4BEG;
	wire [9:0] Tile_X1Y4_bot2top;
	wire [3:0] Tile_X1Y4_E1BEG;
	wire [7:0] Tile_X1Y4_E2BEG;
	wire [7:0] Tile_X1Y4_E2BEGb;
	wire [15:0] Tile_X1Y4_EE4BEG;
	wire [11:0] Tile_X1Y4_E6BEG;
	wire [3:0] Tile_X1Y4_S1BEG;
	wire [7:0] Tile_X1Y4_S2BEG;
	wire [7:0] Tile_X1Y4_S2BEGb;
	wire [15:0] Tile_X1Y4_S4BEG;
	wire [15:0] Tile_X1Y4_SS4BEG;
	wire [3:0] Tile_X1Y4_W1BEG;
	wire [7:0] Tile_X1Y4_W2BEG;
	wire [7:0] Tile_X1Y4_W2BEGb;
	wire [15:0] Tile_X1Y4_WW4BEG;
	wire [11:0] Tile_X1Y4_W6BEG;
	wire [3:0] Tile_X2Y4_N1BEG;
	wire [7:0] Tile_X2Y4_N2BEG;
	wire [7:0] Tile_X2Y4_N2BEGb;
	wire [15:0] Tile_X2Y4_N4BEG;
	wire [15:0] Tile_X2Y4_NN4BEG;
	wire [0:0] Tile_X2Y4_Co;
	wire [3:0] Tile_X2Y4_E1BEG;
	wire [7:0] Tile_X2Y4_E2BEG;
	wire [7:0] Tile_X2Y4_E2BEGb;
	wire [15:0] Tile_X2Y4_EE4BEG;
	wire [11:0] Tile_X2Y4_E6BEG;
	wire [3:0] Tile_X2Y4_S1BEG;
	wire [7:0] Tile_X2Y4_S2BEG;
	wire [7:0] Tile_X2Y4_S2BEGb;
	wire [15:0] Tile_X2Y4_S4BEG;
	wire [15:0] Tile_X2Y4_SS4BEG;
	wire [3:0] Tile_X2Y4_W1BEG;
	wire [7:0] Tile_X2Y4_W2BEG;
	wire [7:0] Tile_X2Y4_W2BEGb;
	wire [15:0] Tile_X2Y4_WW4BEG;
	wire [11:0] Tile_X2Y4_W6BEG;
	wire [3:0] Tile_X3Y4_N1BEG;
	wire [7:0] Tile_X3Y4_N2BEG;
	wire [7:0] Tile_X3Y4_N2BEGb;
	wire [15:0] Tile_X3Y4_N4BEG;
	wire [15:0] Tile_X3Y4_NN4BEG;
	wire [0:0] Tile_X3Y4_Co;
	wire [3:0] Tile_X3Y4_E1BEG;
	wire [7:0] Tile_X3Y4_E2BEG;
	wire [7:0] Tile_X3Y4_E2BEGb;
	wire [15:0] Tile_X3Y4_EE4BEG;
	wire [11:0] Tile_X3Y4_E6BEG;
	wire [3:0] Tile_X3Y4_S1BEG;
	wire [7:0] Tile_X3Y4_S2BEG;
	wire [7:0] Tile_X3Y4_S2BEGb;
	wire [15:0] Tile_X3Y4_S4BEG;
	wire [15:0] Tile_X3Y4_SS4BEG;
	wire [3:0] Tile_X3Y4_W1BEG;
	wire [7:0] Tile_X3Y4_W2BEG;
	wire [7:0] Tile_X3Y4_W2BEGb;
	wire [15:0] Tile_X3Y4_WW4BEG;
	wire [11:0] Tile_X3Y4_W6BEG;
	wire [3:0] Tile_X4Y4_N1BEG;
	wire [7:0] Tile_X4Y4_N2BEG;
	wire [7:0] Tile_X4Y4_N2BEGb;
	wire [15:0] Tile_X4Y4_N4BEG;
	wire [15:0] Tile_X4Y4_NN4BEG;
	wire [0:0] Tile_X4Y4_Co;
	wire [3:0] Tile_X4Y4_E1BEG;
	wire [7:0] Tile_X4Y4_E2BEG;
	wire [7:0] Tile_X4Y4_E2BEGb;
	wire [15:0] Tile_X4Y4_EE4BEG;
	wire [11:0] Tile_X4Y4_E6BEG;
	wire [3:0] Tile_X4Y4_S1BEG;
	wire [7:0] Tile_X4Y4_S2BEG;
	wire [7:0] Tile_X4Y4_S2BEGb;
	wire [15:0] Tile_X4Y4_S4BEG;
	wire [15:0] Tile_X4Y4_SS4BEG;
	wire [3:0] Tile_X4Y4_W1BEG;
	wire [7:0] Tile_X4Y4_W2BEG;
	wire [7:0] Tile_X4Y4_W2BEGb;
	wire [15:0] Tile_X4Y4_WW4BEG;
	wire [11:0] Tile_X4Y4_W6BEG;
	wire [3:0] Tile_X5Y4_N1BEG;
	wire [7:0] Tile_X5Y4_N2BEG;
	wire [7:0] Tile_X5Y4_N2BEGb;
	wire [15:0] Tile_X5Y4_N4BEG;
	wire [15:0] Tile_X5Y4_NN4BEG;
	wire [9:0] Tile_X5Y4_bot2top;
	wire [3:0] Tile_X5Y4_E1BEG;
	wire [7:0] Tile_X5Y4_E2BEG;
	wire [7:0] Tile_X5Y4_E2BEGb;
	wire [15:0] Tile_X5Y4_EE4BEG;
	wire [11:0] Tile_X5Y4_E6BEG;
	wire [3:0] Tile_X5Y4_S1BEG;
	wire [7:0] Tile_X5Y4_S2BEG;
	wire [7:0] Tile_X5Y4_S2BEGb;
	wire [15:0] Tile_X5Y4_S4BEG;
	wire [15:0] Tile_X5Y4_SS4BEG;
	wire [3:0] Tile_X5Y4_W1BEG;
	wire [7:0] Tile_X5Y4_W2BEG;
	wire [7:0] Tile_X5Y4_W2BEGb;
	wire [15:0] Tile_X5Y4_WW4BEG;
	wire [11:0] Tile_X5Y4_W6BEG;
	wire [3:0] Tile_X6Y4_N1BEG;
	wire [7:0] Tile_X6Y4_N2BEG;
	wire [7:0] Tile_X6Y4_N2BEGb;
	wire [15:0] Tile_X6Y4_N4BEG;
	wire [15:0] Tile_X6Y4_NN4BEG;
	wire [0:0] Tile_X6Y4_Co;
	wire [3:0] Tile_X6Y4_E1BEG;
	wire [7:0] Tile_X6Y4_E2BEG;
	wire [7:0] Tile_X6Y4_E2BEGb;
	wire [15:0] Tile_X6Y4_EE4BEG;
	wire [11:0] Tile_X6Y4_E6BEG;
	wire [3:0] Tile_X6Y4_S1BEG;
	wire [7:0] Tile_X6Y4_S2BEG;
	wire [7:0] Tile_X6Y4_S2BEGb;
	wire [15:0] Tile_X6Y4_S4BEG;
	wire [15:0] Tile_X6Y4_SS4BEG;
	wire [3:0] Tile_X6Y4_W1BEG;
	wire [7:0] Tile_X6Y4_W2BEG;
	wire [7:0] Tile_X6Y4_W2BEGb;
	wire [15:0] Tile_X6Y4_WW4BEG;
	wire [11:0] Tile_X6Y4_W6BEG;
	wire [3:0] Tile_X7Y4_W1BEG;
	wire [7:0] Tile_X7Y4_W2BEG;
	wire [7:0] Tile_X7Y4_W2BEGb;
	wire [15:0] Tile_X7Y4_WW4BEG;
	wire [11:0] Tile_X7Y4_W6BEG;
	wire [3:0] Tile_X0Y5_E1BEG;
	wire [7:0] Tile_X0Y5_E2BEG;
	wire [7:0] Tile_X0Y5_E2BEGb;
	wire [15:0] Tile_X0Y5_EE4BEG;
	wire [11:0] Tile_X0Y5_E6BEG;
	wire [3:0] Tile_X1Y5_N1BEG;
	wire [7:0] Tile_X1Y5_N2BEG;
	wire [7:0] Tile_X1Y5_N2BEGb;
	wire [15:0] Tile_X1Y5_N4BEG;
	wire [15:0] Tile_X1Y5_NN4BEG;
	wire [3:0] Tile_X1Y5_E1BEG;
	wire [7:0] Tile_X1Y5_E2BEG;
	wire [7:0] Tile_X1Y5_E2BEGb;
	wire [15:0] Tile_X1Y5_EE4BEG;
	wire [11:0] Tile_X1Y5_E6BEG;
	wire [3:0] Tile_X1Y5_S1BEG;
	wire [7:0] Tile_X1Y5_S2BEG;
	wire [7:0] Tile_X1Y5_S2BEGb;
	wire [15:0] Tile_X1Y5_S4BEG;
	wire [15:0] Tile_X1Y5_SS4BEG;
	wire [17:0] Tile_X1Y5_top2bot;
	wire [3:0] Tile_X1Y5_W1BEG;
	wire [7:0] Tile_X1Y5_W2BEG;
	wire [7:0] Tile_X1Y5_W2BEGb;
	wire [15:0] Tile_X1Y5_WW4BEG;
	wire [11:0] Tile_X1Y5_W6BEG;
	wire [3:0] Tile_X2Y5_N1BEG;
	wire [7:0] Tile_X2Y5_N2BEG;
	wire [7:0] Tile_X2Y5_N2BEGb;
	wire [15:0] Tile_X2Y5_N4BEG;
	wire [15:0] Tile_X2Y5_NN4BEG;
	wire [0:0] Tile_X2Y5_Co;
	wire [3:0] Tile_X2Y5_E1BEG;
	wire [7:0] Tile_X2Y5_E2BEG;
	wire [7:0] Tile_X2Y5_E2BEGb;
	wire [15:0] Tile_X2Y5_EE4BEG;
	wire [11:0] Tile_X2Y5_E6BEG;
	wire [3:0] Tile_X2Y5_S1BEG;
	wire [7:0] Tile_X2Y5_S2BEG;
	wire [7:0] Tile_X2Y5_S2BEGb;
	wire [15:0] Tile_X2Y5_S4BEG;
	wire [15:0] Tile_X2Y5_SS4BEG;
	wire [3:0] Tile_X2Y5_W1BEG;
	wire [7:0] Tile_X2Y5_W2BEG;
	wire [7:0] Tile_X2Y5_W2BEGb;
	wire [15:0] Tile_X2Y5_WW4BEG;
	wire [11:0] Tile_X2Y5_W6BEG;
	wire [3:0] Tile_X3Y5_N1BEG;
	wire [7:0] Tile_X3Y5_N2BEG;
	wire [7:0] Tile_X3Y5_N2BEGb;
	wire [15:0] Tile_X3Y5_N4BEG;
	wire [15:0] Tile_X3Y5_NN4BEG;
	wire [0:0] Tile_X3Y5_Co;
	wire [3:0] Tile_X3Y5_E1BEG;
	wire [7:0] Tile_X3Y5_E2BEG;
	wire [7:0] Tile_X3Y5_E2BEGb;
	wire [15:0] Tile_X3Y5_EE4BEG;
	wire [11:0] Tile_X3Y5_E6BEG;
	wire [3:0] Tile_X3Y5_S1BEG;
	wire [7:0] Tile_X3Y5_S2BEG;
	wire [7:0] Tile_X3Y5_S2BEGb;
	wire [15:0] Tile_X3Y5_S4BEG;
	wire [15:0] Tile_X3Y5_SS4BEG;
	wire [3:0] Tile_X3Y5_W1BEG;
	wire [7:0] Tile_X3Y5_W2BEG;
	wire [7:0] Tile_X3Y5_W2BEGb;
	wire [15:0] Tile_X3Y5_WW4BEG;
	wire [11:0] Tile_X3Y5_W6BEG;
	wire [3:0] Tile_X4Y5_N1BEG;
	wire [7:0] Tile_X4Y5_N2BEG;
	wire [7:0] Tile_X4Y5_N2BEGb;
	wire [15:0] Tile_X4Y5_N4BEG;
	wire [15:0] Tile_X4Y5_NN4BEG;
	wire [0:0] Tile_X4Y5_Co;
	wire [3:0] Tile_X4Y5_E1BEG;
	wire [7:0] Tile_X4Y5_E2BEG;
	wire [7:0] Tile_X4Y5_E2BEGb;
	wire [15:0] Tile_X4Y5_EE4BEG;
	wire [11:0] Tile_X4Y5_E6BEG;
	wire [3:0] Tile_X4Y5_S1BEG;
	wire [7:0] Tile_X4Y5_S2BEG;
	wire [7:0] Tile_X4Y5_S2BEGb;
	wire [15:0] Tile_X4Y5_S4BEG;
	wire [15:0] Tile_X4Y5_SS4BEG;
	wire [3:0] Tile_X4Y5_W1BEG;
	wire [7:0] Tile_X4Y5_W2BEG;
	wire [7:0] Tile_X4Y5_W2BEGb;
	wire [15:0] Tile_X4Y5_WW4BEG;
	wire [11:0] Tile_X4Y5_W6BEG;
	wire [3:0] Tile_X5Y5_N1BEG;
	wire [7:0] Tile_X5Y5_N2BEG;
	wire [7:0] Tile_X5Y5_N2BEGb;
	wire [15:0] Tile_X5Y5_N4BEG;
	wire [15:0] Tile_X5Y5_NN4BEG;
	wire [3:0] Tile_X5Y5_E1BEG;
	wire [7:0] Tile_X5Y5_E2BEG;
	wire [7:0] Tile_X5Y5_E2BEGb;
	wire [15:0] Tile_X5Y5_EE4BEG;
	wire [11:0] Tile_X5Y5_E6BEG;
	wire [3:0] Tile_X5Y5_S1BEG;
	wire [7:0] Tile_X5Y5_S2BEG;
	wire [7:0] Tile_X5Y5_S2BEGb;
	wire [15:0] Tile_X5Y5_S4BEG;
	wire [15:0] Tile_X5Y5_SS4BEG;
	wire [17:0] Tile_X5Y5_top2bot;
	wire [3:0] Tile_X5Y5_W1BEG;
	wire [7:0] Tile_X5Y5_W2BEG;
	wire [7:0] Tile_X5Y5_W2BEGb;
	wire [15:0] Tile_X5Y5_WW4BEG;
	wire [11:0] Tile_X5Y5_W6BEG;
	wire [3:0] Tile_X6Y5_N1BEG;
	wire [7:0] Tile_X6Y5_N2BEG;
	wire [7:0] Tile_X6Y5_N2BEGb;
	wire [15:0] Tile_X6Y5_N4BEG;
	wire [15:0] Tile_X6Y5_NN4BEG;
	wire [0:0] Tile_X6Y5_Co;
	wire [3:0] Tile_X6Y5_E1BEG;
	wire [7:0] Tile_X6Y5_E2BEG;
	wire [7:0] Tile_X6Y5_E2BEGb;
	wire [15:0] Tile_X6Y5_EE4BEG;
	wire [11:0] Tile_X6Y5_E6BEG;
	wire [3:0] Tile_X6Y5_S1BEG;
	wire [7:0] Tile_X6Y5_S2BEG;
	wire [7:0] Tile_X6Y5_S2BEGb;
	wire [15:0] Tile_X6Y5_S4BEG;
	wire [15:0] Tile_X6Y5_SS4BEG;
	wire [3:0] Tile_X6Y5_W1BEG;
	wire [7:0] Tile_X6Y5_W2BEG;
	wire [7:0] Tile_X6Y5_W2BEGb;
	wire [15:0] Tile_X6Y5_WW4BEG;
	wire [11:0] Tile_X6Y5_W6BEG;
	wire [3:0] Tile_X7Y5_W1BEG;
	wire [7:0] Tile_X7Y5_W2BEG;
	wire [7:0] Tile_X7Y5_W2BEGb;
	wire [15:0] Tile_X7Y5_WW4BEG;
	wire [11:0] Tile_X7Y5_W6BEG;
	wire [3:0] Tile_X0Y6_E1BEG;
	wire [7:0] Tile_X0Y6_E2BEG;
	wire [7:0] Tile_X0Y6_E2BEGb;
	wire [15:0] Tile_X0Y6_EE4BEG;
	wire [11:0] Tile_X0Y6_E6BEG;
	wire [3:0] Tile_X1Y6_N1BEG;
	wire [7:0] Tile_X1Y6_N2BEG;
	wire [7:0] Tile_X1Y6_N2BEGb;
	wire [15:0] Tile_X1Y6_N4BEG;
	wire [15:0] Tile_X1Y6_NN4BEG;
	wire [9:0] Tile_X1Y6_bot2top;
	wire [3:0] Tile_X1Y6_E1BEG;
	wire [7:0] Tile_X1Y6_E2BEG;
	wire [7:0] Tile_X1Y6_E2BEGb;
	wire [15:0] Tile_X1Y6_EE4BEG;
	wire [11:0] Tile_X1Y6_E6BEG;
	wire [3:0] Tile_X1Y6_S1BEG;
	wire [7:0] Tile_X1Y6_S2BEG;
	wire [7:0] Tile_X1Y6_S2BEGb;
	wire [15:0] Tile_X1Y6_S4BEG;
	wire [15:0] Tile_X1Y6_SS4BEG;
	wire [3:0] Tile_X1Y6_W1BEG;
	wire [7:0] Tile_X1Y6_W2BEG;
	wire [7:0] Tile_X1Y6_W2BEGb;
	wire [15:0] Tile_X1Y6_WW4BEG;
	wire [11:0] Tile_X1Y6_W6BEG;
	wire [3:0] Tile_X2Y6_N1BEG;
	wire [7:0] Tile_X2Y6_N2BEG;
	wire [7:0] Tile_X2Y6_N2BEGb;
	wire [15:0] Tile_X2Y6_N4BEG;
	wire [15:0] Tile_X2Y6_NN4BEG;
	wire [0:0] Tile_X2Y6_Co;
	wire [3:0] Tile_X2Y6_E1BEG;
	wire [7:0] Tile_X2Y6_E2BEG;
	wire [7:0] Tile_X2Y6_E2BEGb;
	wire [15:0] Tile_X2Y6_EE4BEG;
	wire [11:0] Tile_X2Y6_E6BEG;
	wire [3:0] Tile_X2Y6_S1BEG;
	wire [7:0] Tile_X2Y6_S2BEG;
	wire [7:0] Tile_X2Y6_S2BEGb;
	wire [15:0] Tile_X2Y6_S4BEG;
	wire [15:0] Tile_X2Y6_SS4BEG;
	wire [3:0] Tile_X2Y6_W1BEG;
	wire [7:0] Tile_X2Y6_W2BEG;
	wire [7:0] Tile_X2Y6_W2BEGb;
	wire [15:0] Tile_X2Y6_WW4BEG;
	wire [11:0] Tile_X2Y6_W6BEG;
	wire [3:0] Tile_X3Y6_N1BEG;
	wire [7:0] Tile_X3Y6_N2BEG;
	wire [7:0] Tile_X3Y6_N2BEGb;
	wire [15:0] Tile_X3Y6_N4BEG;
	wire [15:0] Tile_X3Y6_NN4BEG;
	wire [0:0] Tile_X3Y6_Co;
	wire [3:0] Tile_X3Y6_E1BEG;
	wire [7:0] Tile_X3Y6_E2BEG;
	wire [7:0] Tile_X3Y6_E2BEGb;
	wire [15:0] Tile_X3Y6_EE4BEG;
	wire [11:0] Tile_X3Y6_E6BEG;
	wire [3:0] Tile_X3Y6_S1BEG;
	wire [7:0] Tile_X3Y6_S2BEG;
	wire [7:0] Tile_X3Y6_S2BEGb;
	wire [15:0] Tile_X3Y6_S4BEG;
	wire [15:0] Tile_X3Y6_SS4BEG;
	wire [3:0] Tile_X3Y6_W1BEG;
	wire [7:0] Tile_X3Y6_W2BEG;
	wire [7:0] Tile_X3Y6_W2BEGb;
	wire [15:0] Tile_X3Y6_WW4BEG;
	wire [11:0] Tile_X3Y6_W6BEG;
	wire [3:0] Tile_X4Y6_N1BEG;
	wire [7:0] Tile_X4Y6_N2BEG;
	wire [7:0] Tile_X4Y6_N2BEGb;
	wire [15:0] Tile_X4Y6_N4BEG;
	wire [15:0] Tile_X4Y6_NN4BEG;
	wire [0:0] Tile_X4Y6_Co;
	wire [3:0] Tile_X4Y6_E1BEG;
	wire [7:0] Tile_X4Y6_E2BEG;
	wire [7:0] Tile_X4Y6_E2BEGb;
	wire [15:0] Tile_X4Y6_EE4BEG;
	wire [11:0] Tile_X4Y6_E6BEG;
	wire [3:0] Tile_X4Y6_S1BEG;
	wire [7:0] Tile_X4Y6_S2BEG;
	wire [7:0] Tile_X4Y6_S2BEGb;
	wire [15:0] Tile_X4Y6_S4BEG;
	wire [15:0] Tile_X4Y6_SS4BEG;
	wire [3:0] Tile_X4Y6_W1BEG;
	wire [7:0] Tile_X4Y6_W2BEG;
	wire [7:0] Tile_X4Y6_W2BEGb;
	wire [15:0] Tile_X4Y6_WW4BEG;
	wire [11:0] Tile_X4Y6_W6BEG;
	wire [3:0] Tile_X5Y6_N1BEG;
	wire [7:0] Tile_X5Y6_N2BEG;
	wire [7:0] Tile_X5Y6_N2BEGb;
	wire [15:0] Tile_X5Y6_N4BEG;
	wire [15:0] Tile_X5Y6_NN4BEG;
	wire [9:0] Tile_X5Y6_bot2top;
	wire [3:0] Tile_X5Y6_E1BEG;
	wire [7:0] Tile_X5Y6_E2BEG;
	wire [7:0] Tile_X5Y6_E2BEGb;
	wire [15:0] Tile_X5Y6_EE4BEG;
	wire [11:0] Tile_X5Y6_E6BEG;
	wire [3:0] Tile_X5Y6_S1BEG;
	wire [7:0] Tile_X5Y6_S2BEG;
	wire [7:0] Tile_X5Y6_S2BEGb;
	wire [15:0] Tile_X5Y6_S4BEG;
	wire [15:0] Tile_X5Y6_SS4BEG;
	wire [3:0] Tile_X5Y6_W1BEG;
	wire [7:0] Tile_X5Y6_W2BEG;
	wire [7:0] Tile_X5Y6_W2BEGb;
	wire [15:0] Tile_X5Y6_WW4BEG;
	wire [11:0] Tile_X5Y6_W6BEG;
	wire [3:0] Tile_X6Y6_N1BEG;
	wire [7:0] Tile_X6Y6_N2BEG;
	wire [7:0] Tile_X6Y6_N2BEGb;
	wire [15:0] Tile_X6Y6_N4BEG;
	wire [15:0] Tile_X6Y6_NN4BEG;
	wire [0:0] Tile_X6Y6_Co;
	wire [3:0] Tile_X6Y6_E1BEG;
	wire [7:0] Tile_X6Y6_E2BEG;
	wire [7:0] Tile_X6Y6_E2BEGb;
	wire [15:0] Tile_X6Y6_EE4BEG;
	wire [11:0] Tile_X6Y6_E6BEG;
	wire [3:0] Tile_X6Y6_S1BEG;
	wire [7:0] Tile_X6Y6_S2BEG;
	wire [7:0] Tile_X6Y6_S2BEGb;
	wire [15:0] Tile_X6Y6_S4BEG;
	wire [15:0] Tile_X6Y6_SS4BEG;
	wire [3:0] Tile_X6Y6_W1BEG;
	wire [7:0] Tile_X6Y6_W2BEG;
	wire [7:0] Tile_X6Y6_W2BEGb;
	wire [15:0] Tile_X6Y6_WW4BEG;
	wire [11:0] Tile_X6Y6_W6BEG;
	wire [3:0] Tile_X7Y6_W1BEG;
	wire [7:0] Tile_X7Y6_W2BEG;
	wire [7:0] Tile_X7Y6_W2BEGb;
	wire [15:0] Tile_X7Y6_WW4BEG;
	wire [11:0] Tile_X7Y6_W6BEG;
	wire [3:0] Tile_X0Y7_E1BEG;
	wire [7:0] Tile_X0Y7_E2BEG;
	wire [7:0] Tile_X0Y7_E2BEGb;
	wire [15:0] Tile_X0Y7_EE4BEG;
	wire [11:0] Tile_X0Y7_E6BEG;
	wire [3:0] Tile_X1Y7_N1BEG;
	wire [7:0] Tile_X1Y7_N2BEG;
	wire [7:0] Tile_X1Y7_N2BEGb;
	wire [15:0] Tile_X1Y7_N4BEG;
	wire [15:0] Tile_X1Y7_NN4BEG;
	wire [3:0] Tile_X1Y7_E1BEG;
	wire [7:0] Tile_X1Y7_E2BEG;
	wire [7:0] Tile_X1Y7_E2BEGb;
	wire [15:0] Tile_X1Y7_EE4BEG;
	wire [11:0] Tile_X1Y7_E6BEG;
	wire [3:0] Tile_X1Y7_S1BEG;
	wire [7:0] Tile_X1Y7_S2BEG;
	wire [7:0] Tile_X1Y7_S2BEGb;
	wire [15:0] Tile_X1Y7_S4BEG;
	wire [15:0] Tile_X1Y7_SS4BEG;
	wire [17:0] Tile_X1Y7_top2bot;
	wire [3:0] Tile_X1Y7_W1BEG;
	wire [7:0] Tile_X1Y7_W2BEG;
	wire [7:0] Tile_X1Y7_W2BEGb;
	wire [15:0] Tile_X1Y7_WW4BEG;
	wire [11:0] Tile_X1Y7_W6BEG;
	wire [3:0] Tile_X2Y7_N1BEG;
	wire [7:0] Tile_X2Y7_N2BEG;
	wire [7:0] Tile_X2Y7_N2BEGb;
	wire [15:0] Tile_X2Y7_N4BEG;
	wire [15:0] Tile_X2Y7_NN4BEG;
	wire [0:0] Tile_X2Y7_Co;
	wire [3:0] Tile_X2Y7_E1BEG;
	wire [7:0] Tile_X2Y7_E2BEG;
	wire [7:0] Tile_X2Y7_E2BEGb;
	wire [15:0] Tile_X2Y7_EE4BEG;
	wire [11:0] Tile_X2Y7_E6BEG;
	wire [3:0] Tile_X2Y7_S1BEG;
	wire [7:0] Tile_X2Y7_S2BEG;
	wire [7:0] Tile_X2Y7_S2BEGb;
	wire [15:0] Tile_X2Y7_S4BEG;
	wire [15:0] Tile_X2Y7_SS4BEG;
	wire [3:0] Tile_X2Y7_W1BEG;
	wire [7:0] Tile_X2Y7_W2BEG;
	wire [7:0] Tile_X2Y7_W2BEGb;
	wire [15:0] Tile_X2Y7_WW4BEG;
	wire [11:0] Tile_X2Y7_W6BEG;
	wire [3:0] Tile_X3Y7_N1BEG;
	wire [7:0] Tile_X3Y7_N2BEG;
	wire [7:0] Tile_X3Y7_N2BEGb;
	wire [15:0] Tile_X3Y7_N4BEG;
	wire [15:0] Tile_X3Y7_NN4BEG;
	wire [0:0] Tile_X3Y7_Co;
	wire [3:0] Tile_X3Y7_E1BEG;
	wire [7:0] Tile_X3Y7_E2BEG;
	wire [7:0] Tile_X3Y7_E2BEGb;
	wire [15:0] Tile_X3Y7_EE4BEG;
	wire [11:0] Tile_X3Y7_E6BEG;
	wire [3:0] Tile_X3Y7_S1BEG;
	wire [7:0] Tile_X3Y7_S2BEG;
	wire [7:0] Tile_X3Y7_S2BEGb;
	wire [15:0] Tile_X3Y7_S4BEG;
	wire [15:0] Tile_X3Y7_SS4BEG;
	wire [3:0] Tile_X3Y7_W1BEG;
	wire [7:0] Tile_X3Y7_W2BEG;
	wire [7:0] Tile_X3Y7_W2BEGb;
	wire [15:0] Tile_X3Y7_WW4BEG;
	wire [11:0] Tile_X3Y7_W6BEG;
	wire [3:0] Tile_X4Y7_N1BEG;
	wire [7:0] Tile_X4Y7_N2BEG;
	wire [7:0] Tile_X4Y7_N2BEGb;
	wire [15:0] Tile_X4Y7_N4BEG;
	wire [15:0] Tile_X4Y7_NN4BEG;
	wire [0:0] Tile_X4Y7_Co;
	wire [3:0] Tile_X4Y7_E1BEG;
	wire [7:0] Tile_X4Y7_E2BEG;
	wire [7:0] Tile_X4Y7_E2BEGb;
	wire [15:0] Tile_X4Y7_EE4BEG;
	wire [11:0] Tile_X4Y7_E6BEG;
	wire [3:0] Tile_X4Y7_S1BEG;
	wire [7:0] Tile_X4Y7_S2BEG;
	wire [7:0] Tile_X4Y7_S2BEGb;
	wire [15:0] Tile_X4Y7_S4BEG;
	wire [15:0] Tile_X4Y7_SS4BEG;
	wire [3:0] Tile_X4Y7_W1BEG;
	wire [7:0] Tile_X4Y7_W2BEG;
	wire [7:0] Tile_X4Y7_W2BEGb;
	wire [15:0] Tile_X4Y7_WW4BEG;
	wire [11:0] Tile_X4Y7_W6BEG;
	wire [3:0] Tile_X5Y7_N1BEG;
	wire [7:0] Tile_X5Y7_N2BEG;
	wire [7:0] Tile_X5Y7_N2BEGb;
	wire [15:0] Tile_X5Y7_N4BEG;
	wire [15:0] Tile_X5Y7_NN4BEG;
	wire [3:0] Tile_X5Y7_E1BEG;
	wire [7:0] Tile_X5Y7_E2BEG;
	wire [7:0] Tile_X5Y7_E2BEGb;
	wire [15:0] Tile_X5Y7_EE4BEG;
	wire [11:0] Tile_X5Y7_E6BEG;
	wire [3:0] Tile_X5Y7_S1BEG;
	wire [7:0] Tile_X5Y7_S2BEG;
	wire [7:0] Tile_X5Y7_S2BEGb;
	wire [15:0] Tile_X5Y7_S4BEG;
	wire [15:0] Tile_X5Y7_SS4BEG;
	wire [17:0] Tile_X5Y7_top2bot;
	wire [3:0] Tile_X5Y7_W1BEG;
	wire [7:0] Tile_X5Y7_W2BEG;
	wire [7:0] Tile_X5Y7_W2BEGb;
	wire [15:0] Tile_X5Y7_WW4BEG;
	wire [11:0] Tile_X5Y7_W6BEG;
	wire [3:0] Tile_X6Y7_N1BEG;
	wire [7:0] Tile_X6Y7_N2BEG;
	wire [7:0] Tile_X6Y7_N2BEGb;
	wire [15:0] Tile_X6Y7_N4BEG;
	wire [15:0] Tile_X6Y7_NN4BEG;
	wire [0:0] Tile_X6Y7_Co;
	wire [3:0] Tile_X6Y7_E1BEG;
	wire [7:0] Tile_X6Y7_E2BEG;
	wire [7:0] Tile_X6Y7_E2BEGb;
	wire [15:0] Tile_X6Y7_EE4BEG;
	wire [11:0] Tile_X6Y7_E6BEG;
	wire [3:0] Tile_X6Y7_S1BEG;
	wire [7:0] Tile_X6Y7_S2BEG;
	wire [7:0] Tile_X6Y7_S2BEGb;
	wire [15:0] Tile_X6Y7_S4BEG;
	wire [15:0] Tile_X6Y7_SS4BEG;
	wire [3:0] Tile_X6Y7_W1BEG;
	wire [7:0] Tile_X6Y7_W2BEG;
	wire [7:0] Tile_X6Y7_W2BEGb;
	wire [15:0] Tile_X6Y7_WW4BEG;
	wire [11:0] Tile_X6Y7_W6BEG;
	wire [3:0] Tile_X7Y7_W1BEG;
	wire [7:0] Tile_X7Y7_W2BEG;
	wire [7:0] Tile_X7Y7_W2BEGb;
	wire [15:0] Tile_X7Y7_WW4BEG;
	wire [11:0] Tile_X7Y7_W6BEG;
	wire [3:0] Tile_X0Y8_E1BEG;
	wire [7:0] Tile_X0Y8_E2BEG;
	wire [7:0] Tile_X0Y8_E2BEGb;
	wire [15:0] Tile_X0Y8_EE4BEG;
	wire [11:0] Tile_X0Y8_E6BEG;
	wire [3:0] Tile_X1Y8_N1BEG;
	wire [7:0] Tile_X1Y8_N2BEG;
	wire [7:0] Tile_X1Y8_N2BEGb;
	wire [15:0] Tile_X1Y8_N4BEG;
	wire [15:0] Tile_X1Y8_NN4BEG;
	wire [9:0] Tile_X1Y8_bot2top;
	wire [3:0] Tile_X1Y8_E1BEG;
	wire [7:0] Tile_X1Y8_E2BEG;
	wire [7:0] Tile_X1Y8_E2BEGb;
	wire [15:0] Tile_X1Y8_EE4BEG;
	wire [11:0] Tile_X1Y8_E6BEG;
	wire [3:0] Tile_X1Y8_S1BEG;
	wire [7:0] Tile_X1Y8_S2BEG;
	wire [7:0] Tile_X1Y8_S2BEGb;
	wire [15:0] Tile_X1Y8_S4BEG;
	wire [15:0] Tile_X1Y8_SS4BEG;
	wire [3:0] Tile_X1Y8_W1BEG;
	wire [7:0] Tile_X1Y8_W2BEG;
	wire [7:0] Tile_X1Y8_W2BEGb;
	wire [15:0] Tile_X1Y8_WW4BEG;
	wire [11:0] Tile_X1Y8_W6BEG;
	wire [3:0] Tile_X2Y8_N1BEG;
	wire [7:0] Tile_X2Y8_N2BEG;
	wire [7:0] Tile_X2Y8_N2BEGb;
	wire [15:0] Tile_X2Y8_N4BEG;
	wire [15:0] Tile_X2Y8_NN4BEG;
	wire [0:0] Tile_X2Y8_Co;
	wire [3:0] Tile_X2Y8_E1BEG;
	wire [7:0] Tile_X2Y8_E2BEG;
	wire [7:0] Tile_X2Y8_E2BEGb;
	wire [15:0] Tile_X2Y8_EE4BEG;
	wire [11:0] Tile_X2Y8_E6BEG;
	wire [3:0] Tile_X2Y8_S1BEG;
	wire [7:0] Tile_X2Y8_S2BEG;
	wire [7:0] Tile_X2Y8_S2BEGb;
	wire [15:0] Tile_X2Y8_S4BEG;
	wire [15:0] Tile_X2Y8_SS4BEG;
	wire [3:0] Tile_X2Y8_W1BEG;
	wire [7:0] Tile_X2Y8_W2BEG;
	wire [7:0] Tile_X2Y8_W2BEGb;
	wire [15:0] Tile_X2Y8_WW4BEG;
	wire [11:0] Tile_X2Y8_W6BEG;
	wire [3:0] Tile_X3Y8_N1BEG;
	wire [7:0] Tile_X3Y8_N2BEG;
	wire [7:0] Tile_X3Y8_N2BEGb;
	wire [15:0] Tile_X3Y8_N4BEG;
	wire [15:0] Tile_X3Y8_NN4BEG;
	wire [0:0] Tile_X3Y8_Co;
	wire [3:0] Tile_X3Y8_E1BEG;
	wire [7:0] Tile_X3Y8_E2BEG;
	wire [7:0] Tile_X3Y8_E2BEGb;
	wire [15:0] Tile_X3Y8_EE4BEG;
	wire [11:0] Tile_X3Y8_E6BEG;
	wire [3:0] Tile_X3Y8_S1BEG;
	wire [7:0] Tile_X3Y8_S2BEG;
	wire [7:0] Tile_X3Y8_S2BEGb;
	wire [15:0] Tile_X3Y8_S4BEG;
	wire [15:0] Tile_X3Y8_SS4BEG;
	wire [3:0] Tile_X3Y8_W1BEG;
	wire [7:0] Tile_X3Y8_W2BEG;
	wire [7:0] Tile_X3Y8_W2BEGb;
	wire [15:0] Tile_X3Y8_WW4BEG;
	wire [11:0] Tile_X3Y8_W6BEG;
	wire [3:0] Tile_X4Y8_N1BEG;
	wire [7:0] Tile_X4Y8_N2BEG;
	wire [7:0] Tile_X4Y8_N2BEGb;
	wire [15:0] Tile_X4Y8_N4BEG;
	wire [15:0] Tile_X4Y8_NN4BEG;
	wire [0:0] Tile_X4Y8_Co;
	wire [3:0] Tile_X4Y8_E1BEG;
	wire [7:0] Tile_X4Y8_E2BEG;
	wire [7:0] Tile_X4Y8_E2BEGb;
	wire [15:0] Tile_X4Y8_EE4BEG;
	wire [11:0] Tile_X4Y8_E6BEG;
	wire [3:0] Tile_X4Y8_S1BEG;
	wire [7:0] Tile_X4Y8_S2BEG;
	wire [7:0] Tile_X4Y8_S2BEGb;
	wire [15:0] Tile_X4Y8_S4BEG;
	wire [15:0] Tile_X4Y8_SS4BEG;
	wire [3:0] Tile_X4Y8_W1BEG;
	wire [7:0] Tile_X4Y8_W2BEG;
	wire [7:0] Tile_X4Y8_W2BEGb;
	wire [15:0] Tile_X4Y8_WW4BEG;
	wire [11:0] Tile_X4Y8_W6BEG;
	wire [3:0] Tile_X5Y8_N1BEG;
	wire [7:0] Tile_X5Y8_N2BEG;
	wire [7:0] Tile_X5Y8_N2BEGb;
	wire [15:0] Tile_X5Y8_N4BEG;
	wire [15:0] Tile_X5Y8_NN4BEG;
	wire [9:0] Tile_X5Y8_bot2top;
	wire [3:0] Tile_X5Y8_E1BEG;
	wire [7:0] Tile_X5Y8_E2BEG;
	wire [7:0] Tile_X5Y8_E2BEGb;
	wire [15:0] Tile_X5Y8_EE4BEG;
	wire [11:0] Tile_X5Y8_E6BEG;
	wire [3:0] Tile_X5Y8_S1BEG;
	wire [7:0] Tile_X5Y8_S2BEG;
	wire [7:0] Tile_X5Y8_S2BEGb;
	wire [15:0] Tile_X5Y8_S4BEG;
	wire [15:0] Tile_X5Y8_SS4BEG;
	wire [3:0] Tile_X5Y8_W1BEG;
	wire [7:0] Tile_X5Y8_W2BEG;
	wire [7:0] Tile_X5Y8_W2BEGb;
	wire [15:0] Tile_X5Y8_WW4BEG;
	wire [11:0] Tile_X5Y8_W6BEG;
	wire [3:0] Tile_X6Y8_N1BEG;
	wire [7:0] Tile_X6Y8_N2BEG;
	wire [7:0] Tile_X6Y8_N2BEGb;
	wire [15:0] Tile_X6Y8_N4BEG;
	wire [15:0] Tile_X6Y8_NN4BEG;
	wire [0:0] Tile_X6Y8_Co;
	wire [3:0] Tile_X6Y8_E1BEG;
	wire [7:0] Tile_X6Y8_E2BEG;
	wire [7:0] Tile_X6Y8_E2BEGb;
	wire [15:0] Tile_X6Y8_EE4BEG;
	wire [11:0] Tile_X6Y8_E6BEG;
	wire [3:0] Tile_X6Y8_S1BEG;
	wire [7:0] Tile_X6Y8_S2BEG;
	wire [7:0] Tile_X6Y8_S2BEGb;
	wire [15:0] Tile_X6Y8_S4BEG;
	wire [15:0] Tile_X6Y8_SS4BEG;
	wire [3:0] Tile_X6Y8_W1BEG;
	wire [7:0] Tile_X6Y8_W2BEG;
	wire [7:0] Tile_X6Y8_W2BEGb;
	wire [15:0] Tile_X6Y8_WW4BEG;
	wire [11:0] Tile_X6Y8_W6BEG;
	wire [3:0] Tile_X7Y8_W1BEG;
	wire [7:0] Tile_X7Y8_W2BEG;
	wire [7:0] Tile_X7Y8_W2BEGb;
	wire [15:0] Tile_X7Y8_WW4BEG;
	wire [11:0] Tile_X7Y8_W6BEG;
	wire [3:0] Tile_X0Y9_E1BEG;
	wire [7:0] Tile_X0Y9_E2BEG;
	wire [7:0] Tile_X0Y9_E2BEGb;
	wire [15:0] Tile_X0Y9_EE4BEG;
	wire [11:0] Tile_X0Y9_E6BEG;
	wire [3:0] Tile_X1Y9_N1BEG;
	wire [7:0] Tile_X1Y9_N2BEG;
	wire [7:0] Tile_X1Y9_N2BEGb;
	wire [15:0] Tile_X1Y9_N4BEG;
	wire [15:0] Tile_X1Y9_NN4BEG;
	wire [3:0] Tile_X1Y9_E1BEG;
	wire [7:0] Tile_X1Y9_E2BEG;
	wire [7:0] Tile_X1Y9_E2BEGb;
	wire [15:0] Tile_X1Y9_EE4BEG;
	wire [11:0] Tile_X1Y9_E6BEG;
	wire [3:0] Tile_X1Y9_S1BEG;
	wire [7:0] Tile_X1Y9_S2BEG;
	wire [7:0] Tile_X1Y9_S2BEGb;
	wire [15:0] Tile_X1Y9_S4BEG;
	wire [15:0] Tile_X1Y9_SS4BEG;
	wire [17:0] Tile_X1Y9_top2bot;
	wire [3:0] Tile_X1Y9_W1BEG;
	wire [7:0] Tile_X1Y9_W2BEG;
	wire [7:0] Tile_X1Y9_W2BEGb;
	wire [15:0] Tile_X1Y9_WW4BEG;
	wire [11:0] Tile_X1Y9_W6BEG;
	wire [3:0] Tile_X2Y9_N1BEG;
	wire [7:0] Tile_X2Y9_N2BEG;
	wire [7:0] Tile_X2Y9_N2BEGb;
	wire [15:0] Tile_X2Y9_N4BEG;
	wire [15:0] Tile_X2Y9_NN4BEG;
	wire [0:0] Tile_X2Y9_Co;
	wire [3:0] Tile_X2Y9_E1BEG;
	wire [7:0] Tile_X2Y9_E2BEG;
	wire [7:0] Tile_X2Y9_E2BEGb;
	wire [15:0] Tile_X2Y9_EE4BEG;
	wire [11:0] Tile_X2Y9_E6BEG;
	wire [3:0] Tile_X2Y9_S1BEG;
	wire [7:0] Tile_X2Y9_S2BEG;
	wire [7:0] Tile_X2Y9_S2BEGb;
	wire [15:0] Tile_X2Y9_S4BEG;
	wire [15:0] Tile_X2Y9_SS4BEG;
	wire [3:0] Tile_X2Y9_W1BEG;
	wire [7:0] Tile_X2Y9_W2BEG;
	wire [7:0] Tile_X2Y9_W2BEGb;
	wire [15:0] Tile_X2Y9_WW4BEG;
	wire [11:0] Tile_X2Y9_W6BEG;
	wire [3:0] Tile_X3Y9_N1BEG;
	wire [7:0] Tile_X3Y9_N2BEG;
	wire [7:0] Tile_X3Y9_N2BEGb;
	wire [15:0] Tile_X3Y9_N4BEG;
	wire [15:0] Tile_X3Y9_NN4BEG;
	wire [0:0] Tile_X3Y9_Co;
	wire [3:0] Tile_X3Y9_E1BEG;
	wire [7:0] Tile_X3Y9_E2BEG;
	wire [7:0] Tile_X3Y9_E2BEGb;
	wire [15:0] Tile_X3Y9_EE4BEG;
	wire [11:0] Tile_X3Y9_E6BEG;
	wire [3:0] Tile_X3Y9_S1BEG;
	wire [7:0] Tile_X3Y9_S2BEG;
	wire [7:0] Tile_X3Y9_S2BEGb;
	wire [15:0] Tile_X3Y9_S4BEG;
	wire [15:0] Tile_X3Y9_SS4BEG;
	wire [3:0] Tile_X3Y9_W1BEG;
	wire [7:0] Tile_X3Y9_W2BEG;
	wire [7:0] Tile_X3Y9_W2BEGb;
	wire [15:0] Tile_X3Y9_WW4BEG;
	wire [11:0] Tile_X3Y9_W6BEG;
	wire [3:0] Tile_X4Y9_N1BEG;
	wire [7:0] Tile_X4Y9_N2BEG;
	wire [7:0] Tile_X4Y9_N2BEGb;
	wire [15:0] Tile_X4Y9_N4BEG;
	wire [15:0] Tile_X4Y9_NN4BEG;
	wire [0:0] Tile_X4Y9_Co;
	wire [3:0] Tile_X4Y9_E1BEG;
	wire [7:0] Tile_X4Y9_E2BEG;
	wire [7:0] Tile_X4Y9_E2BEGb;
	wire [15:0] Tile_X4Y9_EE4BEG;
	wire [11:0] Tile_X4Y9_E6BEG;
	wire [3:0] Tile_X4Y9_S1BEG;
	wire [7:0] Tile_X4Y9_S2BEG;
	wire [7:0] Tile_X4Y9_S2BEGb;
	wire [15:0] Tile_X4Y9_S4BEG;
	wire [15:0] Tile_X4Y9_SS4BEG;
	wire [3:0] Tile_X4Y9_W1BEG;
	wire [7:0] Tile_X4Y9_W2BEG;
	wire [7:0] Tile_X4Y9_W2BEGb;
	wire [15:0] Tile_X4Y9_WW4BEG;
	wire [11:0] Tile_X4Y9_W6BEG;
	wire [3:0] Tile_X5Y9_N1BEG;
	wire [7:0] Tile_X5Y9_N2BEG;
	wire [7:0] Tile_X5Y9_N2BEGb;
	wire [15:0] Tile_X5Y9_N4BEG;
	wire [15:0] Tile_X5Y9_NN4BEG;
	wire [3:0] Tile_X5Y9_E1BEG;
	wire [7:0] Tile_X5Y9_E2BEG;
	wire [7:0] Tile_X5Y9_E2BEGb;
	wire [15:0] Tile_X5Y9_EE4BEG;
	wire [11:0] Tile_X5Y9_E6BEG;
	wire [3:0] Tile_X5Y9_S1BEG;
	wire [7:0] Tile_X5Y9_S2BEG;
	wire [7:0] Tile_X5Y9_S2BEGb;
	wire [15:0] Tile_X5Y9_S4BEG;
	wire [15:0] Tile_X5Y9_SS4BEG;
	wire [17:0] Tile_X5Y9_top2bot;
	wire [3:0] Tile_X5Y9_W1BEG;
	wire [7:0] Tile_X5Y9_W2BEG;
	wire [7:0] Tile_X5Y9_W2BEGb;
	wire [15:0] Tile_X5Y9_WW4BEG;
	wire [11:0] Tile_X5Y9_W6BEG;
	wire [3:0] Tile_X6Y9_N1BEG;
	wire [7:0] Tile_X6Y9_N2BEG;
	wire [7:0] Tile_X6Y9_N2BEGb;
	wire [15:0] Tile_X6Y9_N4BEG;
	wire [15:0] Tile_X6Y9_NN4BEG;
	wire [0:0] Tile_X6Y9_Co;
	wire [3:0] Tile_X6Y9_E1BEG;
	wire [7:0] Tile_X6Y9_E2BEG;
	wire [7:0] Tile_X6Y9_E2BEGb;
	wire [15:0] Tile_X6Y9_EE4BEG;
	wire [11:0] Tile_X6Y9_E6BEG;
	wire [3:0] Tile_X6Y9_S1BEG;
	wire [7:0] Tile_X6Y9_S2BEG;
	wire [7:0] Tile_X6Y9_S2BEGb;
	wire [15:0] Tile_X6Y9_S4BEG;
	wire [15:0] Tile_X6Y9_SS4BEG;
	wire [3:0] Tile_X6Y9_W1BEG;
	wire [7:0] Tile_X6Y9_W2BEG;
	wire [7:0] Tile_X6Y9_W2BEGb;
	wire [15:0] Tile_X6Y9_WW4BEG;
	wire [11:0] Tile_X6Y9_W6BEG;
	wire [3:0] Tile_X7Y9_W1BEG;
	wire [7:0] Tile_X7Y9_W2BEG;
	wire [7:0] Tile_X7Y9_W2BEGb;
	wire [15:0] Tile_X7Y9_WW4BEG;
	wire [11:0] Tile_X7Y9_W6BEG;
	wire [3:0] Tile_X0Y10_E1BEG;
	wire [7:0] Tile_X0Y10_E2BEG;
	wire [7:0] Tile_X0Y10_E2BEGb;
	wire [15:0] Tile_X0Y10_EE4BEG;
	wire [11:0] Tile_X0Y10_E6BEG;
	wire [3:0] Tile_X1Y10_N1BEG;
	wire [7:0] Tile_X1Y10_N2BEG;
	wire [7:0] Tile_X1Y10_N2BEGb;
	wire [15:0] Tile_X1Y10_N4BEG;
	wire [15:0] Tile_X1Y10_NN4BEG;
	wire [9:0] Tile_X1Y10_bot2top;
	wire [3:0] Tile_X1Y10_E1BEG;
	wire [7:0] Tile_X1Y10_E2BEG;
	wire [7:0] Tile_X1Y10_E2BEGb;
	wire [15:0] Tile_X1Y10_EE4BEG;
	wire [11:0] Tile_X1Y10_E6BEG;
	wire [3:0] Tile_X1Y10_S1BEG;
	wire [7:0] Tile_X1Y10_S2BEG;
	wire [7:0] Tile_X1Y10_S2BEGb;
	wire [15:0] Tile_X1Y10_S4BEG;
	wire [15:0] Tile_X1Y10_SS4BEG;
	wire [3:0] Tile_X1Y10_W1BEG;
	wire [7:0] Tile_X1Y10_W2BEG;
	wire [7:0] Tile_X1Y10_W2BEGb;
	wire [15:0] Tile_X1Y10_WW4BEG;
	wire [11:0] Tile_X1Y10_W6BEG;
	wire [3:0] Tile_X2Y10_N1BEG;
	wire [7:0] Tile_X2Y10_N2BEG;
	wire [7:0] Tile_X2Y10_N2BEGb;
	wire [15:0] Tile_X2Y10_N4BEG;
	wire [15:0] Tile_X2Y10_NN4BEG;
	wire [0:0] Tile_X2Y10_Co;
	wire [3:0] Tile_X2Y10_E1BEG;
	wire [7:0] Tile_X2Y10_E2BEG;
	wire [7:0] Tile_X2Y10_E2BEGb;
	wire [15:0] Tile_X2Y10_EE4BEG;
	wire [11:0] Tile_X2Y10_E6BEG;
	wire [3:0] Tile_X2Y10_S1BEG;
	wire [7:0] Tile_X2Y10_S2BEG;
	wire [7:0] Tile_X2Y10_S2BEGb;
	wire [15:0] Tile_X2Y10_S4BEG;
	wire [15:0] Tile_X2Y10_SS4BEG;
	wire [3:0] Tile_X2Y10_W1BEG;
	wire [7:0] Tile_X2Y10_W2BEG;
	wire [7:0] Tile_X2Y10_W2BEGb;
	wire [15:0] Tile_X2Y10_WW4BEG;
	wire [11:0] Tile_X2Y10_W6BEG;
	wire [3:0] Tile_X3Y10_N1BEG;
	wire [7:0] Tile_X3Y10_N2BEG;
	wire [7:0] Tile_X3Y10_N2BEGb;
	wire [15:0] Tile_X3Y10_N4BEG;
	wire [15:0] Tile_X3Y10_NN4BEG;
	wire [0:0] Tile_X3Y10_Co;
	wire [3:0] Tile_X3Y10_E1BEG;
	wire [7:0] Tile_X3Y10_E2BEG;
	wire [7:0] Tile_X3Y10_E2BEGb;
	wire [15:0] Tile_X3Y10_EE4BEG;
	wire [11:0] Tile_X3Y10_E6BEG;
	wire [3:0] Tile_X3Y10_S1BEG;
	wire [7:0] Tile_X3Y10_S2BEG;
	wire [7:0] Tile_X3Y10_S2BEGb;
	wire [15:0] Tile_X3Y10_S4BEG;
	wire [15:0] Tile_X3Y10_SS4BEG;
	wire [3:0] Tile_X3Y10_W1BEG;
	wire [7:0] Tile_X3Y10_W2BEG;
	wire [7:0] Tile_X3Y10_W2BEGb;
	wire [15:0] Tile_X3Y10_WW4BEG;
	wire [11:0] Tile_X3Y10_W6BEG;
	wire [3:0] Tile_X4Y10_N1BEG;
	wire [7:0] Tile_X4Y10_N2BEG;
	wire [7:0] Tile_X4Y10_N2BEGb;
	wire [15:0] Tile_X4Y10_N4BEG;
	wire [15:0] Tile_X4Y10_NN4BEG;
	wire [0:0] Tile_X4Y10_Co;
	wire [3:0] Tile_X4Y10_E1BEG;
	wire [7:0] Tile_X4Y10_E2BEG;
	wire [7:0] Tile_X4Y10_E2BEGb;
	wire [15:0] Tile_X4Y10_EE4BEG;
	wire [11:0] Tile_X4Y10_E6BEG;
	wire [3:0] Tile_X4Y10_S1BEG;
	wire [7:0] Tile_X4Y10_S2BEG;
	wire [7:0] Tile_X4Y10_S2BEGb;
	wire [15:0] Tile_X4Y10_S4BEG;
	wire [15:0] Tile_X4Y10_SS4BEG;
	wire [3:0] Tile_X4Y10_W1BEG;
	wire [7:0] Tile_X4Y10_W2BEG;
	wire [7:0] Tile_X4Y10_W2BEGb;
	wire [15:0] Tile_X4Y10_WW4BEG;
	wire [11:0] Tile_X4Y10_W6BEG;
	wire [3:0] Tile_X5Y10_N1BEG;
	wire [7:0] Tile_X5Y10_N2BEG;
	wire [7:0] Tile_X5Y10_N2BEGb;
	wire [15:0] Tile_X5Y10_N4BEG;
	wire [15:0] Tile_X5Y10_NN4BEG;
	wire [9:0] Tile_X5Y10_bot2top;
	wire [3:0] Tile_X5Y10_E1BEG;
	wire [7:0] Tile_X5Y10_E2BEG;
	wire [7:0] Tile_X5Y10_E2BEGb;
	wire [15:0] Tile_X5Y10_EE4BEG;
	wire [11:0] Tile_X5Y10_E6BEG;
	wire [3:0] Tile_X5Y10_S1BEG;
	wire [7:0] Tile_X5Y10_S2BEG;
	wire [7:0] Tile_X5Y10_S2BEGb;
	wire [15:0] Tile_X5Y10_S4BEG;
	wire [15:0] Tile_X5Y10_SS4BEG;
	wire [3:0] Tile_X5Y10_W1BEG;
	wire [7:0] Tile_X5Y10_W2BEG;
	wire [7:0] Tile_X5Y10_W2BEGb;
	wire [15:0] Tile_X5Y10_WW4BEG;
	wire [11:0] Tile_X5Y10_W6BEG;
	wire [3:0] Tile_X6Y10_N1BEG;
	wire [7:0] Tile_X6Y10_N2BEG;
	wire [7:0] Tile_X6Y10_N2BEGb;
	wire [15:0] Tile_X6Y10_N4BEG;
	wire [15:0] Tile_X6Y10_NN4BEG;
	wire [0:0] Tile_X6Y10_Co;
	wire [3:0] Tile_X6Y10_E1BEG;
	wire [7:0] Tile_X6Y10_E2BEG;
	wire [7:0] Tile_X6Y10_E2BEGb;
	wire [15:0] Tile_X6Y10_EE4BEG;
	wire [11:0] Tile_X6Y10_E6BEG;
	wire [3:0] Tile_X6Y10_S1BEG;
	wire [7:0] Tile_X6Y10_S2BEG;
	wire [7:0] Tile_X6Y10_S2BEGb;
	wire [15:0] Tile_X6Y10_S4BEG;
	wire [15:0] Tile_X6Y10_SS4BEG;
	wire [3:0] Tile_X6Y10_W1BEG;
	wire [7:0] Tile_X6Y10_W2BEG;
	wire [7:0] Tile_X6Y10_W2BEGb;
	wire [15:0] Tile_X6Y10_WW4BEG;
	wire [11:0] Tile_X6Y10_W6BEG;
	wire [3:0] Tile_X7Y10_W1BEG;
	wire [7:0] Tile_X7Y10_W2BEG;
	wire [7:0] Tile_X7Y10_W2BEGb;
	wire [15:0] Tile_X7Y10_WW4BEG;
	wire [11:0] Tile_X7Y10_W6BEG;
	wire [3:0] Tile_X1Y11_N1BEG;
	wire [7:0] Tile_X1Y11_N2BEG;
	wire [7:0] Tile_X1Y11_N2BEGb;
	wire [15:0] Tile_X1Y11_N4BEG;
	wire [15:0] Tile_X1Y11_NN4BEG;
	wire [3:0] Tile_X2Y11_N1BEG;
	wire [7:0] Tile_X2Y11_N2BEG;
	wire [7:0] Tile_X2Y11_N2BEGb;
	wire [15:0] Tile_X2Y11_N4BEG;
	wire [15:0] Tile_X2Y11_NN4BEG;
	wire [0:0] Tile_X2Y11_Co;
	wire [3:0] Tile_X3Y11_N1BEG;
	wire [7:0] Tile_X3Y11_N2BEG;
	wire [7:0] Tile_X3Y11_N2BEGb;
	wire [15:0] Tile_X3Y11_N4BEG;
	wire [15:0] Tile_X3Y11_NN4BEG;
	wire [0:0] Tile_X3Y11_Co;
	wire [3:0] Tile_X4Y11_N1BEG;
	wire [7:0] Tile_X4Y11_N2BEG;
	wire [7:0] Tile_X4Y11_N2BEGb;
	wire [15:0] Tile_X4Y11_N4BEG;
	wire [15:0] Tile_X4Y11_NN4BEG;
	wire [0:0] Tile_X4Y11_Co;
	wire [3:0] Tile_X5Y11_N1BEG;
	wire [7:0] Tile_X5Y11_N2BEG;
	wire [7:0] Tile_X5Y11_N2BEGb;
	wire [15:0] Tile_X5Y11_N4BEG;
	wire [15:0] Tile_X5Y11_NN4BEG;
	wire [3:0] Tile_X6Y11_N1BEG;
	wire [7:0] Tile_X6Y11_N2BEG;
	wire [7:0] Tile_X6Y11_N2BEGb;
	wire [15:0] Tile_X6Y11_N4BEG;
	wire [15:0] Tile_X6Y11_NN4BEG;
	wire [0:0] Tile_X6Y11_Co;

	assign Tile_Y0_FrameData = FrameData[(FrameBitsPerRow*(0+1))-1:FrameBitsPerRow*0];
	assign Tile_Y1_FrameData = FrameData[(FrameBitsPerRow*(1+1))-1:FrameBitsPerRow*1];
	assign Tile_Y2_FrameData = FrameData[(FrameBitsPerRow*(2+1))-1:FrameBitsPerRow*2];
	assign Tile_Y3_FrameData = FrameData[(FrameBitsPerRow*(3+1))-1:FrameBitsPerRow*3];
	assign Tile_Y4_FrameData = FrameData[(FrameBitsPerRow*(4+1))-1:FrameBitsPerRow*4];
	assign Tile_Y5_FrameData = FrameData[(FrameBitsPerRow*(5+1))-1:FrameBitsPerRow*5];
	assign Tile_Y6_FrameData = FrameData[(FrameBitsPerRow*(6+1))-1:FrameBitsPerRow*6];
	assign Tile_Y7_FrameData = FrameData[(FrameBitsPerRow*(7+1))-1:FrameBitsPerRow*7];
	assign Tile_Y8_FrameData = FrameData[(FrameBitsPerRow*(8+1))-1:FrameBitsPerRow*8];
	assign Tile_Y9_FrameData = FrameData[(FrameBitsPerRow*(9+1))-1:FrameBitsPerRow*9];
	assign Tile_Y10_FrameData = FrameData[(FrameBitsPerRow*(10+1))-1:FrameBitsPerRow*10];
	assign Tile_Y11_FrameData = FrameData[(FrameBitsPerRow*(11+1))-1:FrameBitsPerRow*11];
	assign Tile_X0_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(0+1))-1:MaxFramesPerCol*0];
	assign Tile_X1_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(1+1))-1:MaxFramesPerCol*1];
	assign Tile_X2_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(2+1))-1:MaxFramesPerCol*2];
	assign Tile_X3_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(3+1))-1:MaxFramesPerCol*3];
	assign Tile_X4_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(4+1))-1:MaxFramesPerCol*4];
	assign Tile_X5_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(5+1))-1:MaxFramesPerCol*5];
	assign Tile_X6_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(6+1))-1:MaxFramesPerCol*6];
	assign Tile_X7_FrameStrobe = FrameStrobe[(MaxFramesPerCol*(7+1))-1:MaxFramesPerCol*7];

//tile instantiations

	N_term_DSP Tile_X1Y0_N_term_DSP (
	.N1END(Tile_X1Y1_N1BEG[3:0]),
	.N2MID(Tile_X1Y1_N2BEG[7:0]),
	.N2END(Tile_X1Y1_N2BEGb[7:0]),
	.N4END(Tile_X1Y1_N4BEG[15:0]),
	.NN4END(Tile_X1Y1_NN4BEG[15:0]),
	.S1BEG(Tile_X1Y0_S1BEG[3:0]),
	.S2BEG(Tile_X1Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X1Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X1Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X1Y0_SS4BEG[15:0]),
	.FrameData(Tile_Y0_FrameData), 
	.FrameData_O(Tile_X1Y0_FrameData_O), 
	.FrameStrobe(Tile_X1Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X1Y0_FrameStrobe_O)
	);

	N_term_single Tile_X2Y0_N_term_single (
	.N1END(Tile_X2Y1_N1BEG[3:0]),
	.N2MID(Tile_X2Y1_N2BEG[7:0]),
	.N2END(Tile_X2Y1_N2BEGb[7:0]),
	.N4END(Tile_X2Y1_N4BEG[15:0]),
	.NN4END(Tile_X2Y1_NN4BEG[15:0]),
	.Ci(Tile_X2Y1_Co[0:0]),
	.S1BEG(Tile_X2Y0_S1BEG[3:0]),
	.S2BEG(Tile_X2Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y0_SS4BEG[15:0]),
	.FrameData(Tile_X1Y0_FrameData_O), 
	.FrameData_O(Tile_X2Y0_FrameData_O), 
	.FrameStrobe(Tile_X2Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y0_FrameStrobe_O)
	);

	N_term_single Tile_X3Y0_N_term_single (
	.N1END(Tile_X3Y1_N1BEG[3:0]),
	.N2MID(Tile_X3Y1_N2BEG[7:0]),
	.N2END(Tile_X3Y1_N2BEGb[7:0]),
	.N4END(Tile_X3Y1_N4BEG[15:0]),
	.NN4END(Tile_X3Y1_NN4BEG[15:0]),
	.Ci(Tile_X3Y1_Co[0:0]),
	.S1BEG(Tile_X3Y0_S1BEG[3:0]),
	.S2BEG(Tile_X3Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y0_SS4BEG[15:0]),
	.FrameData(Tile_X2Y0_FrameData_O), 
	.FrameData_O(Tile_X3Y0_FrameData_O), 
	.FrameStrobe(Tile_X3Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y0_FrameStrobe_O)
	);

	N_term_single Tile_X4Y0_N_term_single (
	.N1END(Tile_X4Y1_N1BEG[3:0]),
	.N2MID(Tile_X4Y1_N2BEG[7:0]),
	.N2END(Tile_X4Y1_N2BEGb[7:0]),
	.N4END(Tile_X4Y1_N4BEG[15:0]),
	.NN4END(Tile_X4Y1_NN4BEG[15:0]),
	.Ci(Tile_X4Y1_Co[0:0]),
	.S1BEG(Tile_X4Y0_S1BEG[3:0]),
	.S2BEG(Tile_X4Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y0_SS4BEG[15:0]),
	.FrameData(Tile_X3Y0_FrameData_O), 
	.FrameData_O(Tile_X4Y0_FrameData_O), 
	.FrameStrobe(Tile_X4Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y0_FrameStrobe_O)
	);

	N_term_DSP Tile_X5Y0_N_term_DSP (
	.N1END(Tile_X5Y1_N1BEG[3:0]),
	.N2MID(Tile_X5Y1_N2BEG[7:0]),
	.N2END(Tile_X5Y1_N2BEGb[7:0]),
	.N4END(Tile_X5Y1_N4BEG[15:0]),
	.NN4END(Tile_X5Y1_NN4BEG[15:0]),
	.S1BEG(Tile_X5Y0_S1BEG[3:0]),
	.S2BEG(Tile_X5Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X5Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X5Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X5Y0_SS4BEG[15:0]),
	.FrameData(Tile_X4Y0_FrameData_O), 
	.FrameData_O(Tile_X5Y0_FrameData_O), 
	.FrameStrobe(Tile_X5Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X5Y0_FrameStrobe_O)
	);

	N_term_single Tile_X6Y0_N_term_single (
	.N1END(Tile_X6Y1_N1BEG[3:0]),
	.N2MID(Tile_X6Y1_N2BEG[7:0]),
	.N2END(Tile_X6Y1_N2BEGb[7:0]),
	.N4END(Tile_X6Y1_N4BEG[15:0]),
	.NN4END(Tile_X6Y1_NN4BEG[15:0]),
	.Ci(Tile_X6Y1_Co[0:0]),
	.S1BEG(Tile_X6Y0_S1BEG[3:0]),
	.S2BEG(Tile_X6Y0_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y0_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y0_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y0_SS4BEG[15:0]),
	.FrameData(Tile_X5Y0_FrameData_O), 
	.FrameData_O(Tile_X6Y0_FrameData_O), 
	.FrameStrobe(Tile_X6Y1_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y0_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y1_W_CPU_IO (
	.W1END(Tile_X1Y1_W1BEG[3:0]),
	.W2MID(Tile_X1Y1_W2BEG[7:0]),
	.W2END(Tile_X1Y1_W2BEGb[7:0]),
	.WW4END(Tile_X1Y1_WW4BEG[15:0]),
	.W6END(Tile_X1Y1_W6BEG[11:0]),
	.E1BEG(Tile_X0Y1_E1BEG[3:0]),
	.E2BEG(Tile_X0Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y1_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y1_OPA_I0),
	.OPA_I1(Tile_X0Y1_OPA_I1),
	.OPA_I2(Tile_X0Y1_OPA_I2),
	.OPA_I3(Tile_X0Y1_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y1_OPB_I0),
	.OPB_I1(Tile_X0Y1_OPB_I1),
	.OPB_I2(Tile_X0Y1_OPB_I2),
	.OPB_I3(Tile_X0Y1_OPB_I3),
	.RES0_O0(Tile_X0Y1_RES0_O0),
	.RES0_O1(Tile_X0Y1_RES0_O1),
	.RES0_O2(Tile_X0Y1_RES0_O2),
	.RES0_O3(Tile_X0Y1_RES0_O3),
	.RES1_O0(Tile_X0Y1_RES1_O0),
	.RES1_O1(Tile_X0Y1_RES1_O1),
	.RES1_O2(Tile_X0Y1_RES1_O2),
	.RES1_O3(Tile_X0Y1_RES1_O3),
	.RES2_O0(Tile_X0Y1_RES2_O0),
	.RES2_O1(Tile_X0Y1_RES2_O1),
	.RES2_O2(Tile_X0Y1_RES2_O2),
	.RES2_O3(Tile_X0Y1_RES2_O3),
	.FrameData(Tile_Y1_FrameData), 
	.FrameData_O(Tile_X0Y1_FrameData_O), 
	.FrameStrobe(Tile_X0Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y1_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y1_LUT4AB (
	.N1END(Tile_X2Y2_N1BEG[3:0]),
	.N2MID(Tile_X2Y2_N2BEG[7:0]),
	.N2END(Tile_X2Y2_N2BEGb[7:0]),
	.N4END(Tile_X2Y2_N4BEG[15:0]),
	.NN4END(Tile_X2Y2_NN4BEG[15:0]),
	.Ci(Tile_X2Y2_Co[0:0]),
	.E1END(Tile_X1Y1_E1BEG[3:0]),
	.E2MID(Tile_X1Y1_E2BEG[7:0]),
	.E2END(Tile_X1Y1_E2BEGb[7:0]),
	.EE4END(Tile_X1Y1_EE4BEG[15:0]),
	.E6END(Tile_X1Y1_E6BEG[11:0]),
	.S1END(Tile_X2Y0_S1BEG[3:0]),
	.S2MID(Tile_X2Y0_S2BEG[7:0]),
	.S2END(Tile_X2Y0_S2BEGb[7:0]),
	.S4END(Tile_X2Y0_S4BEG[15:0]),
	.SS4END(Tile_X2Y0_SS4BEG[15:0]),
	.W1END(Tile_X3Y1_W1BEG[3:0]),
	.W2MID(Tile_X3Y1_W2BEG[7:0]),
	.W2END(Tile_X3Y1_W2BEGb[7:0]),
	.WW4END(Tile_X3Y1_WW4BEG[15:0]),
	.W6END(Tile_X3Y1_W6BEG[11:0]),
	.N1BEG(Tile_X2Y1_N1BEG[3:0]),
	.N2BEG(Tile_X2Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y1_NN4BEG[15:0]),
	.Co(Tile_X2Y1_Co[0:0]),
	.E1BEG(Tile_X2Y1_E1BEG[3:0]),
	.E2BEG(Tile_X2Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y1_E6BEG[11:0]),
	.S1BEG(Tile_X2Y1_S1BEG[3:0]),
	.S2BEG(Tile_X2Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y1_W1BEG[3:0]),
	.W2BEG(Tile_X2Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y1_FrameData_O), 
	.FrameData_O(Tile_X2Y1_FrameData_O), 
	.FrameStrobe(Tile_X2Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y1_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y1_LUT4AB (
	.N1END(Tile_X3Y2_N1BEG[3:0]),
	.N2MID(Tile_X3Y2_N2BEG[7:0]),
	.N2END(Tile_X3Y2_N2BEGb[7:0]),
	.N4END(Tile_X3Y2_N4BEG[15:0]),
	.NN4END(Tile_X3Y2_NN4BEG[15:0]),
	.Ci(Tile_X3Y2_Co[0:0]),
	.E1END(Tile_X2Y1_E1BEG[3:0]),
	.E2MID(Tile_X2Y1_E2BEG[7:0]),
	.E2END(Tile_X2Y1_E2BEGb[7:0]),
	.EE4END(Tile_X2Y1_EE4BEG[15:0]),
	.E6END(Tile_X2Y1_E6BEG[11:0]),
	.S1END(Tile_X3Y0_S1BEG[3:0]),
	.S2MID(Tile_X3Y0_S2BEG[7:0]),
	.S2END(Tile_X3Y0_S2BEGb[7:0]),
	.S4END(Tile_X3Y0_S4BEG[15:0]),
	.SS4END(Tile_X3Y0_SS4BEG[15:0]),
	.W1END(Tile_X4Y1_W1BEG[3:0]),
	.W2MID(Tile_X4Y1_W2BEG[7:0]),
	.W2END(Tile_X4Y1_W2BEGb[7:0]),
	.WW4END(Tile_X4Y1_WW4BEG[15:0]),
	.W6END(Tile_X4Y1_W6BEG[11:0]),
	.N1BEG(Tile_X3Y1_N1BEG[3:0]),
	.N2BEG(Tile_X3Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y1_NN4BEG[15:0]),
	.Co(Tile_X3Y1_Co[0:0]),
	.E1BEG(Tile_X3Y1_E1BEG[3:0]),
	.E2BEG(Tile_X3Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y1_E6BEG[11:0]),
	.S1BEG(Tile_X3Y1_S1BEG[3:0]),
	.S2BEG(Tile_X3Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y1_W1BEG[3:0]),
	.W2BEG(Tile_X3Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y1_FrameData_O), 
	.FrameData_O(Tile_X3Y1_FrameData_O), 
	.FrameStrobe(Tile_X3Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y1_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y1_LUT4AB (
	.N1END(Tile_X4Y2_N1BEG[3:0]),
	.N2MID(Tile_X4Y2_N2BEG[7:0]),
	.N2END(Tile_X4Y2_N2BEGb[7:0]),
	.N4END(Tile_X4Y2_N4BEG[15:0]),
	.NN4END(Tile_X4Y2_NN4BEG[15:0]),
	.Ci(Tile_X4Y2_Co[0:0]),
	.E1END(Tile_X3Y1_E1BEG[3:0]),
	.E2MID(Tile_X3Y1_E2BEG[7:0]),
	.E2END(Tile_X3Y1_E2BEGb[7:0]),
	.EE4END(Tile_X3Y1_EE4BEG[15:0]),
	.E6END(Tile_X3Y1_E6BEG[11:0]),
	.S1END(Tile_X4Y0_S1BEG[3:0]),
	.S2MID(Tile_X4Y0_S2BEG[7:0]),
	.S2END(Tile_X4Y0_S2BEGb[7:0]),
	.S4END(Tile_X4Y0_S4BEG[15:0]),
	.SS4END(Tile_X4Y0_SS4BEG[15:0]),
	.W1END(Tile_X5Y1_W1BEG[3:0]),
	.W2MID(Tile_X5Y1_W2BEG[7:0]),
	.W2END(Tile_X5Y1_W2BEGb[7:0]),
	.WW4END(Tile_X5Y1_WW4BEG[15:0]),
	.W6END(Tile_X5Y1_W6BEG[11:0]),
	.N1BEG(Tile_X4Y1_N1BEG[3:0]),
	.N2BEG(Tile_X4Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y1_NN4BEG[15:0]),
	.Co(Tile_X4Y1_Co[0:0]),
	.E1BEG(Tile_X4Y1_E1BEG[3:0]),
	.E2BEG(Tile_X4Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y1_E6BEG[11:0]),
	.S1BEG(Tile_X4Y1_S1BEG[3:0]),
	.S2BEG(Tile_X4Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y1_W1BEG[3:0]),
	.W2BEG(Tile_X4Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y1_FrameData_O), 
	.FrameData_O(Tile_X4Y1_FrameData_O), 
	.FrameStrobe(Tile_X4Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y1_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y1_LUT4AB (
	.N1END(Tile_X6Y2_N1BEG[3:0]),
	.N2MID(Tile_X6Y2_N2BEG[7:0]),
	.N2END(Tile_X6Y2_N2BEGb[7:0]),
	.N4END(Tile_X6Y2_N4BEG[15:0]),
	.NN4END(Tile_X6Y2_NN4BEG[15:0]),
	.Ci(Tile_X6Y2_Co[0:0]),
	.E1END(Tile_X5Y1_E1BEG[3:0]),
	.E2MID(Tile_X5Y1_E2BEG[7:0]),
	.E2END(Tile_X5Y1_E2BEGb[7:0]),
	.EE4END(Tile_X5Y1_EE4BEG[15:0]),
	.E6END(Tile_X5Y1_E6BEG[11:0]),
	.S1END(Tile_X6Y0_S1BEG[3:0]),
	.S2MID(Tile_X6Y0_S2BEG[7:0]),
	.S2END(Tile_X6Y0_S2BEGb[7:0]),
	.S4END(Tile_X6Y0_S4BEG[15:0]),
	.SS4END(Tile_X6Y0_SS4BEG[15:0]),
	.W1END(Tile_X7Y1_W1BEG[3:0]),
	.W2MID(Tile_X7Y1_W2BEG[7:0]),
	.W2END(Tile_X7Y1_W2BEGb[7:0]),
	.WW4END(Tile_X7Y1_WW4BEG[15:0]),
	.W6END(Tile_X7Y1_W6BEG[11:0]),
	.N1BEG(Tile_X6Y1_N1BEG[3:0]),
	.N2BEG(Tile_X6Y1_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y1_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y1_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y1_NN4BEG[15:0]),
	.Co(Tile_X6Y1_Co[0:0]),
	.E1BEG(Tile_X6Y1_E1BEG[3:0]),
	.E2BEG(Tile_X6Y1_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y1_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y1_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y1_E6BEG[11:0]),
	.S1BEG(Tile_X6Y1_S1BEG[3:0]),
	.S2BEG(Tile_X6Y1_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y1_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y1_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y1_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y1_W1BEG[3:0]),
	.W2BEG(Tile_X6Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y1_FrameData_O), 
	.FrameData_O(Tile_X6Y1_FrameData_O), 
	.FrameStrobe(Tile_X6Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y1_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y1_E_CPU_IO (
	.E1END(Tile_X6Y1_E1BEG[3:0]),
	.E2MID(Tile_X6Y1_E2BEG[7:0]),
	.E2END(Tile_X6Y1_E2BEGb[7:0]),
	.EE4END(Tile_X6Y1_EE4BEG[15:0]),
	.E6END(Tile_X6Y1_E6BEG[11:0]),
	.W1BEG(Tile_X7Y1_W1BEG[3:0]),
	.W2BEG(Tile_X7Y1_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y1_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y1_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y1_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y1_OPA_I0),
	.OPA_I1(Tile_X7Y1_OPA_I1),
	.OPA_I2(Tile_X7Y1_OPA_I2),
	.OPA_I3(Tile_X7Y1_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y1_OPB_I0),
	.OPB_I1(Tile_X7Y1_OPB_I1),
	.OPB_I2(Tile_X7Y1_OPB_I2),
	.OPB_I3(Tile_X7Y1_OPB_I3),
	.RES0_O0(Tile_X7Y1_RES0_O0),
	.RES0_O1(Tile_X7Y1_RES0_O1),
	.RES0_O2(Tile_X7Y1_RES0_O2),
	.RES0_O3(Tile_X7Y1_RES0_O3),
	.RES1_O0(Tile_X7Y1_RES1_O0),
	.RES1_O1(Tile_X7Y1_RES1_O1),
	.RES1_O2(Tile_X7Y1_RES1_O2),
	.RES1_O3(Tile_X7Y1_RES1_O3),
	.RES2_O0(Tile_X7Y1_RES2_O0),
	.RES2_O1(Tile_X7Y1_RES2_O1),
	.RES2_O2(Tile_X7Y1_RES2_O2),
	.RES2_O3(Tile_X7Y1_RES2_O3),
	.FrameData(Tile_X6Y1_FrameData_O), 
	.FrameData_O(Tile_X7Y1_FrameData_O), 
	.FrameStrobe(Tile_X7Y2_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y1_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y2_W_CPU_IO (
	.W1END(Tile_X1Y2_W1BEG[3:0]),
	.W2MID(Tile_X1Y2_W2BEG[7:0]),
	.W2END(Tile_X1Y2_W2BEGb[7:0]),
	.WW4END(Tile_X1Y2_WW4BEG[15:0]),
	.W6END(Tile_X1Y2_W6BEG[11:0]),
	.E1BEG(Tile_X0Y2_E1BEG[3:0]),
	.E2BEG(Tile_X0Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y2_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y2_OPA_I0),
	.OPA_I1(Tile_X0Y2_OPA_I1),
	.OPA_I2(Tile_X0Y2_OPA_I2),
	.OPA_I3(Tile_X0Y2_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y2_OPB_I0),
	.OPB_I1(Tile_X0Y2_OPB_I1),
	.OPB_I2(Tile_X0Y2_OPB_I2),
	.OPB_I3(Tile_X0Y2_OPB_I3),
	.RES0_O0(Tile_X0Y2_RES0_O0),
	.RES0_O1(Tile_X0Y2_RES0_O1),
	.RES0_O2(Tile_X0Y2_RES0_O2),
	.RES0_O3(Tile_X0Y2_RES0_O3),
	.RES1_O0(Tile_X0Y2_RES1_O0),
	.RES1_O1(Tile_X0Y2_RES1_O1),
	.RES1_O2(Tile_X0Y2_RES1_O2),
	.RES1_O3(Tile_X0Y2_RES1_O3),
	.RES2_O0(Tile_X0Y2_RES2_O0),
	.RES2_O1(Tile_X0Y2_RES2_O1),
	.RES2_O2(Tile_X0Y2_RES2_O2),
	.RES2_O3(Tile_X0Y2_RES2_O3),
	.FrameData(Tile_Y2_FrameData), 
	.FrameData_O(Tile_X0Y2_FrameData_O), 
	.FrameStrobe(Tile_X0Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y2_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y2_LUT4AB (
	.N1END(Tile_X2Y3_N1BEG[3:0]),
	.N2MID(Tile_X2Y3_N2BEG[7:0]),
	.N2END(Tile_X2Y3_N2BEGb[7:0]),
	.N4END(Tile_X2Y3_N4BEG[15:0]),
	.NN4END(Tile_X2Y3_NN4BEG[15:0]),
	.Ci(Tile_X2Y3_Co[0:0]),
	.E1END(Tile_X1Y2_E1BEG[3:0]),
	.E2MID(Tile_X1Y2_E2BEG[7:0]),
	.E2END(Tile_X1Y2_E2BEGb[7:0]),
	.EE4END(Tile_X1Y2_EE4BEG[15:0]),
	.E6END(Tile_X1Y2_E6BEG[11:0]),
	.S1END(Tile_X2Y1_S1BEG[3:0]),
	.S2MID(Tile_X2Y1_S2BEG[7:0]),
	.S2END(Tile_X2Y1_S2BEGb[7:0]),
	.S4END(Tile_X2Y1_S4BEG[15:0]),
	.SS4END(Tile_X2Y1_SS4BEG[15:0]),
	.W1END(Tile_X3Y2_W1BEG[3:0]),
	.W2MID(Tile_X3Y2_W2BEG[7:0]),
	.W2END(Tile_X3Y2_W2BEGb[7:0]),
	.WW4END(Tile_X3Y2_WW4BEG[15:0]),
	.W6END(Tile_X3Y2_W6BEG[11:0]),
	.N1BEG(Tile_X2Y2_N1BEG[3:0]),
	.N2BEG(Tile_X2Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y2_NN4BEG[15:0]),
	.Co(Tile_X2Y2_Co[0:0]),
	.E1BEG(Tile_X2Y2_E1BEG[3:0]),
	.E2BEG(Tile_X2Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y2_E6BEG[11:0]),
	.S1BEG(Tile_X2Y2_S1BEG[3:0]),
	.S2BEG(Tile_X2Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y2_W1BEG[3:0]),
	.W2BEG(Tile_X2Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y2_FrameData_O), 
	.FrameData_O(Tile_X2Y2_FrameData_O), 
	.FrameStrobe(Tile_X2Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y2_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y2_LUT4AB (
	.N1END(Tile_X3Y3_N1BEG[3:0]),
	.N2MID(Tile_X3Y3_N2BEG[7:0]),
	.N2END(Tile_X3Y3_N2BEGb[7:0]),
	.N4END(Tile_X3Y3_N4BEG[15:0]),
	.NN4END(Tile_X3Y3_NN4BEG[15:0]),
	.Ci(Tile_X3Y3_Co[0:0]),
	.E1END(Tile_X2Y2_E1BEG[3:0]),
	.E2MID(Tile_X2Y2_E2BEG[7:0]),
	.E2END(Tile_X2Y2_E2BEGb[7:0]),
	.EE4END(Tile_X2Y2_EE4BEG[15:0]),
	.E6END(Tile_X2Y2_E6BEG[11:0]),
	.S1END(Tile_X3Y1_S1BEG[3:0]),
	.S2MID(Tile_X3Y1_S2BEG[7:0]),
	.S2END(Tile_X3Y1_S2BEGb[7:0]),
	.S4END(Tile_X3Y1_S4BEG[15:0]),
	.SS4END(Tile_X3Y1_SS4BEG[15:0]),
	.W1END(Tile_X4Y2_W1BEG[3:0]),
	.W2MID(Tile_X4Y2_W2BEG[7:0]),
	.W2END(Tile_X4Y2_W2BEGb[7:0]),
	.WW4END(Tile_X4Y2_WW4BEG[15:0]),
	.W6END(Tile_X4Y2_W6BEG[11:0]),
	.N1BEG(Tile_X3Y2_N1BEG[3:0]),
	.N2BEG(Tile_X3Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y2_NN4BEG[15:0]),
	.Co(Tile_X3Y2_Co[0:0]),
	.E1BEG(Tile_X3Y2_E1BEG[3:0]),
	.E2BEG(Tile_X3Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y2_E6BEG[11:0]),
	.S1BEG(Tile_X3Y2_S1BEG[3:0]),
	.S2BEG(Tile_X3Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y2_W1BEG[3:0]),
	.W2BEG(Tile_X3Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y2_FrameData_O), 
	.FrameData_O(Tile_X3Y2_FrameData_O), 
	.FrameStrobe(Tile_X3Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y2_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y2_LUT4AB (
	.N1END(Tile_X4Y3_N1BEG[3:0]),
	.N2MID(Tile_X4Y3_N2BEG[7:0]),
	.N2END(Tile_X4Y3_N2BEGb[7:0]),
	.N4END(Tile_X4Y3_N4BEG[15:0]),
	.NN4END(Tile_X4Y3_NN4BEG[15:0]),
	.Ci(Tile_X4Y3_Co[0:0]),
	.E1END(Tile_X3Y2_E1BEG[3:0]),
	.E2MID(Tile_X3Y2_E2BEG[7:0]),
	.E2END(Tile_X3Y2_E2BEGb[7:0]),
	.EE4END(Tile_X3Y2_EE4BEG[15:0]),
	.E6END(Tile_X3Y2_E6BEG[11:0]),
	.S1END(Tile_X4Y1_S1BEG[3:0]),
	.S2MID(Tile_X4Y1_S2BEG[7:0]),
	.S2END(Tile_X4Y1_S2BEGb[7:0]),
	.S4END(Tile_X4Y1_S4BEG[15:0]),
	.SS4END(Tile_X4Y1_SS4BEG[15:0]),
	.W1END(Tile_X5Y2_W1BEG[3:0]),
	.W2MID(Tile_X5Y2_W2BEG[7:0]),
	.W2END(Tile_X5Y2_W2BEGb[7:0]),
	.WW4END(Tile_X5Y2_WW4BEG[15:0]),
	.W6END(Tile_X5Y2_W6BEG[11:0]),
	.N1BEG(Tile_X4Y2_N1BEG[3:0]),
	.N2BEG(Tile_X4Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y2_NN4BEG[15:0]),
	.Co(Tile_X4Y2_Co[0:0]),
	.E1BEG(Tile_X4Y2_E1BEG[3:0]),
	.E2BEG(Tile_X4Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y2_E6BEG[11:0]),
	.S1BEG(Tile_X4Y2_S1BEG[3:0]),
	.S2BEG(Tile_X4Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y2_W1BEG[3:0]),
	.W2BEG(Tile_X4Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y2_FrameData_O), 
	.FrameData_O(Tile_X4Y2_FrameData_O), 
	.FrameStrobe(Tile_X4Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y2_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y2_LUT4AB (
	.N1END(Tile_X6Y3_N1BEG[3:0]),
	.N2MID(Tile_X6Y3_N2BEG[7:0]),
	.N2END(Tile_X6Y3_N2BEGb[7:0]),
	.N4END(Tile_X6Y3_N4BEG[15:0]),
	.NN4END(Tile_X6Y3_NN4BEG[15:0]),
	.Ci(Tile_X6Y3_Co[0:0]),
	.E1END(Tile_X5Y2_E1BEG[3:0]),
	.E2MID(Tile_X5Y2_E2BEG[7:0]),
	.E2END(Tile_X5Y2_E2BEGb[7:0]),
	.EE4END(Tile_X5Y2_EE4BEG[15:0]),
	.E6END(Tile_X5Y2_E6BEG[11:0]),
	.S1END(Tile_X6Y1_S1BEG[3:0]),
	.S2MID(Tile_X6Y1_S2BEG[7:0]),
	.S2END(Tile_X6Y1_S2BEGb[7:0]),
	.S4END(Tile_X6Y1_S4BEG[15:0]),
	.SS4END(Tile_X6Y1_SS4BEG[15:0]),
	.W1END(Tile_X7Y2_W1BEG[3:0]),
	.W2MID(Tile_X7Y2_W2BEG[7:0]),
	.W2END(Tile_X7Y2_W2BEGb[7:0]),
	.WW4END(Tile_X7Y2_WW4BEG[15:0]),
	.W6END(Tile_X7Y2_W6BEG[11:0]),
	.N1BEG(Tile_X6Y2_N1BEG[3:0]),
	.N2BEG(Tile_X6Y2_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y2_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y2_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y2_NN4BEG[15:0]),
	.Co(Tile_X6Y2_Co[0:0]),
	.E1BEG(Tile_X6Y2_E1BEG[3:0]),
	.E2BEG(Tile_X6Y2_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y2_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y2_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y2_E6BEG[11:0]),
	.S1BEG(Tile_X6Y2_S1BEG[3:0]),
	.S2BEG(Tile_X6Y2_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y2_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y2_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y2_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y2_W1BEG[3:0]),
	.W2BEG(Tile_X6Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y2_FrameData_O), 
	.FrameData_O(Tile_X6Y2_FrameData_O), 
	.FrameStrobe(Tile_X6Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y2_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y2_E_CPU_IO (
	.E1END(Tile_X6Y2_E1BEG[3:0]),
	.E2MID(Tile_X6Y2_E2BEG[7:0]),
	.E2END(Tile_X6Y2_E2BEGb[7:0]),
	.EE4END(Tile_X6Y2_EE4BEG[15:0]),
	.E6END(Tile_X6Y2_E6BEG[11:0]),
	.W1BEG(Tile_X7Y2_W1BEG[3:0]),
	.W2BEG(Tile_X7Y2_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y2_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y2_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y2_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y2_OPA_I0),
	.OPA_I1(Tile_X7Y2_OPA_I1),
	.OPA_I2(Tile_X7Y2_OPA_I2),
	.OPA_I3(Tile_X7Y2_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y2_OPB_I0),
	.OPB_I1(Tile_X7Y2_OPB_I1),
	.OPB_I2(Tile_X7Y2_OPB_I2),
	.OPB_I3(Tile_X7Y2_OPB_I3),
	.RES0_O0(Tile_X7Y2_RES0_O0),
	.RES0_O1(Tile_X7Y2_RES0_O1),
	.RES0_O2(Tile_X7Y2_RES0_O2),
	.RES0_O3(Tile_X7Y2_RES0_O3),
	.RES1_O0(Tile_X7Y2_RES1_O0),
	.RES1_O1(Tile_X7Y2_RES1_O1),
	.RES1_O2(Tile_X7Y2_RES1_O2),
	.RES1_O3(Tile_X7Y2_RES1_O3),
	.RES2_O0(Tile_X7Y2_RES2_O0),
	.RES2_O1(Tile_X7Y2_RES2_O1),
	.RES2_O2(Tile_X7Y2_RES2_O2),
	.RES2_O3(Tile_X7Y2_RES2_O3),
	.FrameData(Tile_X6Y2_FrameData_O), 
	.FrameData_O(Tile_X7Y2_FrameData_O), 
	.FrameStrobe(Tile_X7Y3_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y2_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y3_W_CPU_IO (
	.W1END(Tile_X1Y3_W1BEG[3:0]),
	.W2MID(Tile_X1Y3_W2BEG[7:0]),
	.W2END(Tile_X1Y3_W2BEGb[7:0]),
	.WW4END(Tile_X1Y3_WW4BEG[15:0]),
	.W6END(Tile_X1Y3_W6BEG[11:0]),
	.E1BEG(Tile_X0Y3_E1BEG[3:0]),
	.E2BEG(Tile_X0Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y3_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y3_OPA_I0),
	.OPA_I1(Tile_X0Y3_OPA_I1),
	.OPA_I2(Tile_X0Y3_OPA_I2),
	.OPA_I3(Tile_X0Y3_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y3_OPB_I0),
	.OPB_I1(Tile_X0Y3_OPB_I1),
	.OPB_I2(Tile_X0Y3_OPB_I2),
	.OPB_I3(Tile_X0Y3_OPB_I3),
	.RES0_O0(Tile_X0Y3_RES0_O0),
	.RES0_O1(Tile_X0Y3_RES0_O1),
	.RES0_O2(Tile_X0Y3_RES0_O2),
	.RES0_O3(Tile_X0Y3_RES0_O3),
	.RES1_O0(Tile_X0Y3_RES1_O0),
	.RES1_O1(Tile_X0Y3_RES1_O1),
	.RES1_O2(Tile_X0Y3_RES1_O2),
	.RES1_O3(Tile_X0Y3_RES1_O3),
	.RES2_O0(Tile_X0Y3_RES2_O0),
	.RES2_O1(Tile_X0Y3_RES2_O1),
	.RES2_O2(Tile_X0Y3_RES2_O2),
	.RES2_O3(Tile_X0Y3_RES2_O3),
	.FrameData(Tile_Y3_FrameData), 
	.FrameData_O(Tile_X0Y3_FrameData_O), 
	.FrameStrobe(Tile_X0Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y3_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y3_LUT4AB (
	.N1END(Tile_X2Y4_N1BEG[3:0]),
	.N2MID(Tile_X2Y4_N2BEG[7:0]),
	.N2END(Tile_X2Y4_N2BEGb[7:0]),
	.N4END(Tile_X2Y4_N4BEG[15:0]),
	.NN4END(Tile_X2Y4_NN4BEG[15:0]),
	.Ci(Tile_X2Y4_Co[0:0]),
	.E1END(Tile_X1Y3_E1BEG[3:0]),
	.E2MID(Tile_X1Y3_E2BEG[7:0]),
	.E2END(Tile_X1Y3_E2BEGb[7:0]),
	.EE4END(Tile_X1Y3_EE4BEG[15:0]),
	.E6END(Tile_X1Y3_E6BEG[11:0]),
	.S1END(Tile_X2Y2_S1BEG[3:0]),
	.S2MID(Tile_X2Y2_S2BEG[7:0]),
	.S2END(Tile_X2Y2_S2BEGb[7:0]),
	.S4END(Tile_X2Y2_S4BEG[15:0]),
	.SS4END(Tile_X2Y2_SS4BEG[15:0]),
	.W1END(Tile_X3Y3_W1BEG[3:0]),
	.W2MID(Tile_X3Y3_W2BEG[7:0]),
	.W2END(Tile_X3Y3_W2BEGb[7:0]),
	.WW4END(Tile_X3Y3_WW4BEG[15:0]),
	.W6END(Tile_X3Y3_W6BEG[11:0]),
	.N1BEG(Tile_X2Y3_N1BEG[3:0]),
	.N2BEG(Tile_X2Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y3_NN4BEG[15:0]),
	.Co(Tile_X2Y3_Co[0:0]),
	.E1BEG(Tile_X2Y3_E1BEG[3:0]),
	.E2BEG(Tile_X2Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y3_E6BEG[11:0]),
	.S1BEG(Tile_X2Y3_S1BEG[3:0]),
	.S2BEG(Tile_X2Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y3_W1BEG[3:0]),
	.W2BEG(Tile_X2Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y3_FrameData_O), 
	.FrameData_O(Tile_X2Y3_FrameData_O), 
	.FrameStrobe(Tile_X2Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y3_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y3_LUT4AB (
	.N1END(Tile_X3Y4_N1BEG[3:0]),
	.N2MID(Tile_X3Y4_N2BEG[7:0]),
	.N2END(Tile_X3Y4_N2BEGb[7:0]),
	.N4END(Tile_X3Y4_N4BEG[15:0]),
	.NN4END(Tile_X3Y4_NN4BEG[15:0]),
	.Ci(Tile_X3Y4_Co[0:0]),
	.E1END(Tile_X2Y3_E1BEG[3:0]),
	.E2MID(Tile_X2Y3_E2BEG[7:0]),
	.E2END(Tile_X2Y3_E2BEGb[7:0]),
	.EE4END(Tile_X2Y3_EE4BEG[15:0]),
	.E6END(Tile_X2Y3_E6BEG[11:0]),
	.S1END(Tile_X3Y2_S1BEG[3:0]),
	.S2MID(Tile_X3Y2_S2BEG[7:0]),
	.S2END(Tile_X3Y2_S2BEGb[7:0]),
	.S4END(Tile_X3Y2_S4BEG[15:0]),
	.SS4END(Tile_X3Y2_SS4BEG[15:0]),
	.W1END(Tile_X4Y3_W1BEG[3:0]),
	.W2MID(Tile_X4Y3_W2BEG[7:0]),
	.W2END(Tile_X4Y3_W2BEGb[7:0]),
	.WW4END(Tile_X4Y3_WW4BEG[15:0]),
	.W6END(Tile_X4Y3_W6BEG[11:0]),
	.N1BEG(Tile_X3Y3_N1BEG[3:0]),
	.N2BEG(Tile_X3Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y3_NN4BEG[15:0]),
	.Co(Tile_X3Y3_Co[0:0]),
	.E1BEG(Tile_X3Y3_E1BEG[3:0]),
	.E2BEG(Tile_X3Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y3_E6BEG[11:0]),
	.S1BEG(Tile_X3Y3_S1BEG[3:0]),
	.S2BEG(Tile_X3Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y3_W1BEG[3:0]),
	.W2BEG(Tile_X3Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y3_FrameData_O), 
	.FrameData_O(Tile_X3Y3_FrameData_O), 
	.FrameStrobe(Tile_X3Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y3_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y3_LUT4AB (
	.N1END(Tile_X4Y4_N1BEG[3:0]),
	.N2MID(Tile_X4Y4_N2BEG[7:0]),
	.N2END(Tile_X4Y4_N2BEGb[7:0]),
	.N4END(Tile_X4Y4_N4BEG[15:0]),
	.NN4END(Tile_X4Y4_NN4BEG[15:0]),
	.Ci(Tile_X4Y4_Co[0:0]),
	.E1END(Tile_X3Y3_E1BEG[3:0]),
	.E2MID(Tile_X3Y3_E2BEG[7:0]),
	.E2END(Tile_X3Y3_E2BEGb[7:0]),
	.EE4END(Tile_X3Y3_EE4BEG[15:0]),
	.E6END(Tile_X3Y3_E6BEG[11:0]),
	.S1END(Tile_X4Y2_S1BEG[3:0]),
	.S2MID(Tile_X4Y2_S2BEG[7:0]),
	.S2END(Tile_X4Y2_S2BEGb[7:0]),
	.S4END(Tile_X4Y2_S4BEG[15:0]),
	.SS4END(Tile_X4Y2_SS4BEG[15:0]),
	.W1END(Tile_X5Y3_W1BEG[3:0]),
	.W2MID(Tile_X5Y3_W2BEG[7:0]),
	.W2END(Tile_X5Y3_W2BEGb[7:0]),
	.WW4END(Tile_X5Y3_WW4BEG[15:0]),
	.W6END(Tile_X5Y3_W6BEG[11:0]),
	.N1BEG(Tile_X4Y3_N1BEG[3:0]),
	.N2BEG(Tile_X4Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y3_NN4BEG[15:0]),
	.Co(Tile_X4Y3_Co[0:0]),
	.E1BEG(Tile_X4Y3_E1BEG[3:0]),
	.E2BEG(Tile_X4Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y3_E6BEG[11:0]),
	.S1BEG(Tile_X4Y3_S1BEG[3:0]),
	.S2BEG(Tile_X4Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y3_W1BEG[3:0]),
	.W2BEG(Tile_X4Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y3_FrameData_O), 
	.FrameData_O(Tile_X4Y3_FrameData_O), 
	.FrameStrobe(Tile_X4Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y3_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y3_LUT4AB (
	.N1END(Tile_X6Y4_N1BEG[3:0]),
	.N2MID(Tile_X6Y4_N2BEG[7:0]),
	.N2END(Tile_X6Y4_N2BEGb[7:0]),
	.N4END(Tile_X6Y4_N4BEG[15:0]),
	.NN4END(Tile_X6Y4_NN4BEG[15:0]),
	.Ci(Tile_X6Y4_Co[0:0]),
	.E1END(Tile_X5Y3_E1BEG[3:0]),
	.E2MID(Tile_X5Y3_E2BEG[7:0]),
	.E2END(Tile_X5Y3_E2BEGb[7:0]),
	.EE4END(Tile_X5Y3_EE4BEG[15:0]),
	.E6END(Tile_X5Y3_E6BEG[11:0]),
	.S1END(Tile_X6Y2_S1BEG[3:0]),
	.S2MID(Tile_X6Y2_S2BEG[7:0]),
	.S2END(Tile_X6Y2_S2BEGb[7:0]),
	.S4END(Tile_X6Y2_S4BEG[15:0]),
	.SS4END(Tile_X6Y2_SS4BEG[15:0]),
	.W1END(Tile_X7Y3_W1BEG[3:0]),
	.W2MID(Tile_X7Y3_W2BEG[7:0]),
	.W2END(Tile_X7Y3_W2BEGb[7:0]),
	.WW4END(Tile_X7Y3_WW4BEG[15:0]),
	.W6END(Tile_X7Y3_W6BEG[11:0]),
	.N1BEG(Tile_X6Y3_N1BEG[3:0]),
	.N2BEG(Tile_X6Y3_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y3_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y3_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y3_NN4BEG[15:0]),
	.Co(Tile_X6Y3_Co[0:0]),
	.E1BEG(Tile_X6Y3_E1BEG[3:0]),
	.E2BEG(Tile_X6Y3_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y3_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y3_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y3_E6BEG[11:0]),
	.S1BEG(Tile_X6Y3_S1BEG[3:0]),
	.S2BEG(Tile_X6Y3_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y3_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y3_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y3_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y3_W1BEG[3:0]),
	.W2BEG(Tile_X6Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y3_FrameData_O), 
	.FrameData_O(Tile_X6Y3_FrameData_O), 
	.FrameStrobe(Tile_X6Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y3_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y3_E_CPU_IO (
	.E1END(Tile_X6Y3_E1BEG[3:0]),
	.E2MID(Tile_X6Y3_E2BEG[7:0]),
	.E2END(Tile_X6Y3_E2BEGb[7:0]),
	.EE4END(Tile_X6Y3_EE4BEG[15:0]),
	.E6END(Tile_X6Y3_E6BEG[11:0]),
	.W1BEG(Tile_X7Y3_W1BEG[3:0]),
	.W2BEG(Tile_X7Y3_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y3_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y3_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y3_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y3_OPA_I0),
	.OPA_I1(Tile_X7Y3_OPA_I1),
	.OPA_I2(Tile_X7Y3_OPA_I2),
	.OPA_I3(Tile_X7Y3_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y3_OPB_I0),
	.OPB_I1(Tile_X7Y3_OPB_I1),
	.OPB_I2(Tile_X7Y3_OPB_I2),
	.OPB_I3(Tile_X7Y3_OPB_I3),
	.RES0_O0(Tile_X7Y3_RES0_O0),
	.RES0_O1(Tile_X7Y3_RES0_O1),
	.RES0_O2(Tile_X7Y3_RES0_O2),
	.RES0_O3(Tile_X7Y3_RES0_O3),
	.RES1_O0(Tile_X7Y3_RES1_O0),
	.RES1_O1(Tile_X7Y3_RES1_O1),
	.RES1_O2(Tile_X7Y3_RES1_O2),
	.RES1_O3(Tile_X7Y3_RES1_O3),
	.RES2_O0(Tile_X7Y3_RES2_O0),
	.RES2_O1(Tile_X7Y3_RES2_O1),
	.RES2_O2(Tile_X7Y3_RES2_O2),
	.RES2_O3(Tile_X7Y3_RES2_O3),
	.FrameData(Tile_X6Y3_FrameData_O), 
	.FrameData_O(Tile_X7Y3_FrameData_O), 
	.FrameStrobe(Tile_X7Y4_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y3_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y4_W_CPU_IO (
	.W1END(Tile_X1Y4_W1BEG[3:0]),
	.W2MID(Tile_X1Y4_W2BEG[7:0]),
	.W2END(Tile_X1Y4_W2BEGb[7:0]),
	.WW4END(Tile_X1Y4_WW4BEG[15:0]),
	.W6END(Tile_X1Y4_W6BEG[11:0]),
	.E1BEG(Tile_X0Y4_E1BEG[3:0]),
	.E2BEG(Tile_X0Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y4_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y4_OPA_I0),
	.OPA_I1(Tile_X0Y4_OPA_I1),
	.OPA_I2(Tile_X0Y4_OPA_I2),
	.OPA_I3(Tile_X0Y4_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y4_OPB_I0),
	.OPB_I1(Tile_X0Y4_OPB_I1),
	.OPB_I2(Tile_X0Y4_OPB_I2),
	.OPB_I3(Tile_X0Y4_OPB_I3),
	.RES0_O0(Tile_X0Y4_RES0_O0),
	.RES0_O1(Tile_X0Y4_RES0_O1),
	.RES0_O2(Tile_X0Y4_RES0_O2),
	.RES0_O3(Tile_X0Y4_RES0_O3),
	.RES1_O0(Tile_X0Y4_RES1_O0),
	.RES1_O1(Tile_X0Y4_RES1_O1),
	.RES1_O2(Tile_X0Y4_RES1_O2),
	.RES1_O3(Tile_X0Y4_RES1_O3),
	.RES2_O0(Tile_X0Y4_RES2_O0),
	.RES2_O1(Tile_X0Y4_RES2_O1),
	.RES2_O2(Tile_X0Y4_RES2_O2),
	.RES2_O3(Tile_X0Y4_RES2_O3),
	.FrameData(Tile_Y4_FrameData), 
	.FrameData_O(Tile_X0Y4_FrameData_O), 
	.FrameStrobe(Tile_X0Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y4_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y4_LUT4AB (
	.N1END(Tile_X2Y5_N1BEG[3:0]),
	.N2MID(Tile_X2Y5_N2BEG[7:0]),
	.N2END(Tile_X2Y5_N2BEGb[7:0]),
	.N4END(Tile_X2Y5_N4BEG[15:0]),
	.NN4END(Tile_X2Y5_NN4BEG[15:0]),
	.Ci(Tile_X2Y5_Co[0:0]),
	.E1END(Tile_X1Y4_E1BEG[3:0]),
	.E2MID(Tile_X1Y4_E2BEG[7:0]),
	.E2END(Tile_X1Y4_E2BEGb[7:0]),
	.EE4END(Tile_X1Y4_EE4BEG[15:0]),
	.E6END(Tile_X1Y4_E6BEG[11:0]),
	.S1END(Tile_X2Y3_S1BEG[3:0]),
	.S2MID(Tile_X2Y3_S2BEG[7:0]),
	.S2END(Tile_X2Y3_S2BEGb[7:0]),
	.S4END(Tile_X2Y3_S4BEG[15:0]),
	.SS4END(Tile_X2Y3_SS4BEG[15:0]),
	.W1END(Tile_X3Y4_W1BEG[3:0]),
	.W2MID(Tile_X3Y4_W2BEG[7:0]),
	.W2END(Tile_X3Y4_W2BEGb[7:0]),
	.WW4END(Tile_X3Y4_WW4BEG[15:0]),
	.W6END(Tile_X3Y4_W6BEG[11:0]),
	.N1BEG(Tile_X2Y4_N1BEG[3:0]),
	.N2BEG(Tile_X2Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y4_NN4BEG[15:0]),
	.Co(Tile_X2Y4_Co[0:0]),
	.E1BEG(Tile_X2Y4_E1BEG[3:0]),
	.E2BEG(Tile_X2Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y4_E6BEG[11:0]),
	.S1BEG(Tile_X2Y4_S1BEG[3:0]),
	.S2BEG(Tile_X2Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y4_W1BEG[3:0]),
	.W2BEG(Tile_X2Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y4_FrameData_O), 
	.FrameData_O(Tile_X2Y4_FrameData_O), 
	.FrameStrobe(Tile_X2Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y4_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y4_LUT4AB (
	.N1END(Tile_X3Y5_N1BEG[3:0]),
	.N2MID(Tile_X3Y5_N2BEG[7:0]),
	.N2END(Tile_X3Y5_N2BEGb[7:0]),
	.N4END(Tile_X3Y5_N4BEG[15:0]),
	.NN4END(Tile_X3Y5_NN4BEG[15:0]),
	.Ci(Tile_X3Y5_Co[0:0]),
	.E1END(Tile_X2Y4_E1BEG[3:0]),
	.E2MID(Tile_X2Y4_E2BEG[7:0]),
	.E2END(Tile_X2Y4_E2BEGb[7:0]),
	.EE4END(Tile_X2Y4_EE4BEG[15:0]),
	.E6END(Tile_X2Y4_E6BEG[11:0]),
	.S1END(Tile_X3Y3_S1BEG[3:0]),
	.S2MID(Tile_X3Y3_S2BEG[7:0]),
	.S2END(Tile_X3Y3_S2BEGb[7:0]),
	.S4END(Tile_X3Y3_S4BEG[15:0]),
	.SS4END(Tile_X3Y3_SS4BEG[15:0]),
	.W1END(Tile_X4Y4_W1BEG[3:0]),
	.W2MID(Tile_X4Y4_W2BEG[7:0]),
	.W2END(Tile_X4Y4_W2BEGb[7:0]),
	.WW4END(Tile_X4Y4_WW4BEG[15:0]),
	.W6END(Tile_X4Y4_W6BEG[11:0]),
	.N1BEG(Tile_X3Y4_N1BEG[3:0]),
	.N2BEG(Tile_X3Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y4_NN4BEG[15:0]),
	.Co(Tile_X3Y4_Co[0:0]),
	.E1BEG(Tile_X3Y4_E1BEG[3:0]),
	.E2BEG(Tile_X3Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y4_E6BEG[11:0]),
	.S1BEG(Tile_X3Y4_S1BEG[3:0]),
	.S2BEG(Tile_X3Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y4_W1BEG[3:0]),
	.W2BEG(Tile_X3Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y4_FrameData_O), 
	.FrameData_O(Tile_X3Y4_FrameData_O), 
	.FrameStrobe(Tile_X3Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y4_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y4_LUT4AB (
	.N1END(Tile_X4Y5_N1BEG[3:0]),
	.N2MID(Tile_X4Y5_N2BEG[7:0]),
	.N2END(Tile_X4Y5_N2BEGb[7:0]),
	.N4END(Tile_X4Y5_N4BEG[15:0]),
	.NN4END(Tile_X4Y5_NN4BEG[15:0]),
	.Ci(Tile_X4Y5_Co[0:0]),
	.E1END(Tile_X3Y4_E1BEG[3:0]),
	.E2MID(Tile_X3Y4_E2BEG[7:0]),
	.E2END(Tile_X3Y4_E2BEGb[7:0]),
	.EE4END(Tile_X3Y4_EE4BEG[15:0]),
	.E6END(Tile_X3Y4_E6BEG[11:0]),
	.S1END(Tile_X4Y3_S1BEG[3:0]),
	.S2MID(Tile_X4Y3_S2BEG[7:0]),
	.S2END(Tile_X4Y3_S2BEGb[7:0]),
	.S4END(Tile_X4Y3_S4BEG[15:0]),
	.SS4END(Tile_X4Y3_SS4BEG[15:0]),
	.W1END(Tile_X5Y4_W1BEG[3:0]),
	.W2MID(Tile_X5Y4_W2BEG[7:0]),
	.W2END(Tile_X5Y4_W2BEGb[7:0]),
	.WW4END(Tile_X5Y4_WW4BEG[15:0]),
	.W6END(Tile_X5Y4_W6BEG[11:0]),
	.N1BEG(Tile_X4Y4_N1BEG[3:0]),
	.N2BEG(Tile_X4Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y4_NN4BEG[15:0]),
	.Co(Tile_X4Y4_Co[0:0]),
	.E1BEG(Tile_X4Y4_E1BEG[3:0]),
	.E2BEG(Tile_X4Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y4_E6BEG[11:0]),
	.S1BEG(Tile_X4Y4_S1BEG[3:0]),
	.S2BEG(Tile_X4Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y4_W1BEG[3:0]),
	.W2BEG(Tile_X4Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y4_FrameData_O), 
	.FrameData_O(Tile_X4Y4_FrameData_O), 
	.FrameStrobe(Tile_X4Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y4_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y4_LUT4AB (
	.N1END(Tile_X6Y5_N1BEG[3:0]),
	.N2MID(Tile_X6Y5_N2BEG[7:0]),
	.N2END(Tile_X6Y5_N2BEGb[7:0]),
	.N4END(Tile_X6Y5_N4BEG[15:0]),
	.NN4END(Tile_X6Y5_NN4BEG[15:0]),
	.Ci(Tile_X6Y5_Co[0:0]),
	.E1END(Tile_X5Y4_E1BEG[3:0]),
	.E2MID(Tile_X5Y4_E2BEG[7:0]),
	.E2END(Tile_X5Y4_E2BEGb[7:0]),
	.EE4END(Tile_X5Y4_EE4BEG[15:0]),
	.E6END(Tile_X5Y4_E6BEG[11:0]),
	.S1END(Tile_X6Y3_S1BEG[3:0]),
	.S2MID(Tile_X6Y3_S2BEG[7:0]),
	.S2END(Tile_X6Y3_S2BEGb[7:0]),
	.S4END(Tile_X6Y3_S4BEG[15:0]),
	.SS4END(Tile_X6Y3_SS4BEG[15:0]),
	.W1END(Tile_X7Y4_W1BEG[3:0]),
	.W2MID(Tile_X7Y4_W2BEG[7:0]),
	.W2END(Tile_X7Y4_W2BEGb[7:0]),
	.WW4END(Tile_X7Y4_WW4BEG[15:0]),
	.W6END(Tile_X7Y4_W6BEG[11:0]),
	.N1BEG(Tile_X6Y4_N1BEG[3:0]),
	.N2BEG(Tile_X6Y4_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y4_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y4_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y4_NN4BEG[15:0]),
	.Co(Tile_X6Y4_Co[0:0]),
	.E1BEG(Tile_X6Y4_E1BEG[3:0]),
	.E2BEG(Tile_X6Y4_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y4_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y4_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y4_E6BEG[11:0]),
	.S1BEG(Tile_X6Y4_S1BEG[3:0]),
	.S2BEG(Tile_X6Y4_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y4_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y4_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y4_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y4_W1BEG[3:0]),
	.W2BEG(Tile_X6Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y4_FrameData_O), 
	.FrameData_O(Tile_X6Y4_FrameData_O), 
	.FrameStrobe(Tile_X6Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y4_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y4_E_CPU_IO (
	.E1END(Tile_X6Y4_E1BEG[3:0]),
	.E2MID(Tile_X6Y4_E2BEG[7:0]),
	.E2END(Tile_X6Y4_E2BEGb[7:0]),
	.EE4END(Tile_X6Y4_EE4BEG[15:0]),
	.E6END(Tile_X6Y4_E6BEG[11:0]),
	.W1BEG(Tile_X7Y4_W1BEG[3:0]),
	.W2BEG(Tile_X7Y4_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y4_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y4_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y4_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y4_OPA_I0),
	.OPA_I1(Tile_X7Y4_OPA_I1),
	.OPA_I2(Tile_X7Y4_OPA_I2),
	.OPA_I3(Tile_X7Y4_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y4_OPB_I0),
	.OPB_I1(Tile_X7Y4_OPB_I1),
	.OPB_I2(Tile_X7Y4_OPB_I2),
	.OPB_I3(Tile_X7Y4_OPB_I3),
	.RES0_O0(Tile_X7Y4_RES0_O0),
	.RES0_O1(Tile_X7Y4_RES0_O1),
	.RES0_O2(Tile_X7Y4_RES0_O2),
	.RES0_O3(Tile_X7Y4_RES0_O3),
	.RES1_O0(Tile_X7Y4_RES1_O0),
	.RES1_O1(Tile_X7Y4_RES1_O1),
	.RES1_O2(Tile_X7Y4_RES1_O2),
	.RES1_O3(Tile_X7Y4_RES1_O3),
	.RES2_O0(Tile_X7Y4_RES2_O0),
	.RES2_O1(Tile_X7Y4_RES2_O1),
	.RES2_O2(Tile_X7Y4_RES2_O2),
	.RES2_O3(Tile_X7Y4_RES2_O3),
	.FrameData(Tile_X6Y4_FrameData_O), 
	.FrameData_O(Tile_X7Y4_FrameData_O), 
	.FrameStrobe(Tile_X7Y5_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y4_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y5_W_CPU_IO (
	.W1END(Tile_X1Y5_W1BEG[3:0]),
	.W2MID(Tile_X1Y5_W2BEG[7:0]),
	.W2END(Tile_X1Y5_W2BEGb[7:0]),
	.WW4END(Tile_X1Y5_WW4BEG[15:0]),
	.W6END(Tile_X1Y5_W6BEG[11:0]),
	.E1BEG(Tile_X0Y5_E1BEG[3:0]),
	.E2BEG(Tile_X0Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y5_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y5_OPA_I0),
	.OPA_I1(Tile_X0Y5_OPA_I1),
	.OPA_I2(Tile_X0Y5_OPA_I2),
	.OPA_I3(Tile_X0Y5_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y5_OPB_I0),
	.OPB_I1(Tile_X0Y5_OPB_I1),
	.OPB_I2(Tile_X0Y5_OPB_I2),
	.OPB_I3(Tile_X0Y5_OPB_I3),
	.RES0_O0(Tile_X0Y5_RES0_O0),
	.RES0_O1(Tile_X0Y5_RES0_O1),
	.RES0_O2(Tile_X0Y5_RES0_O2),
	.RES0_O3(Tile_X0Y5_RES0_O3),
	.RES1_O0(Tile_X0Y5_RES1_O0),
	.RES1_O1(Tile_X0Y5_RES1_O1),
	.RES1_O2(Tile_X0Y5_RES1_O2),
	.RES1_O3(Tile_X0Y5_RES1_O3),
	.RES2_O0(Tile_X0Y5_RES2_O0),
	.RES2_O1(Tile_X0Y5_RES2_O1),
	.RES2_O2(Tile_X0Y5_RES2_O2),
	.RES2_O3(Tile_X0Y5_RES2_O3),
	.FrameData(Tile_Y5_FrameData), 
	.FrameData_O(Tile_X0Y5_FrameData_O), 
	.FrameStrobe(Tile_X0Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y5_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y5_LUT4AB (
	.N1END(Tile_X2Y6_N1BEG[3:0]),
	.N2MID(Tile_X2Y6_N2BEG[7:0]),
	.N2END(Tile_X2Y6_N2BEGb[7:0]),
	.N4END(Tile_X2Y6_N4BEG[15:0]),
	.NN4END(Tile_X2Y6_NN4BEG[15:0]),
	.Ci(Tile_X2Y6_Co[0:0]),
	.E1END(Tile_X1Y5_E1BEG[3:0]),
	.E2MID(Tile_X1Y5_E2BEG[7:0]),
	.E2END(Tile_X1Y5_E2BEGb[7:0]),
	.EE4END(Tile_X1Y5_EE4BEG[15:0]),
	.E6END(Tile_X1Y5_E6BEG[11:0]),
	.S1END(Tile_X2Y4_S1BEG[3:0]),
	.S2MID(Tile_X2Y4_S2BEG[7:0]),
	.S2END(Tile_X2Y4_S2BEGb[7:0]),
	.S4END(Tile_X2Y4_S4BEG[15:0]),
	.SS4END(Tile_X2Y4_SS4BEG[15:0]),
	.W1END(Tile_X3Y5_W1BEG[3:0]),
	.W2MID(Tile_X3Y5_W2BEG[7:0]),
	.W2END(Tile_X3Y5_W2BEGb[7:0]),
	.WW4END(Tile_X3Y5_WW4BEG[15:0]),
	.W6END(Tile_X3Y5_W6BEG[11:0]),
	.N1BEG(Tile_X2Y5_N1BEG[3:0]),
	.N2BEG(Tile_X2Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y5_NN4BEG[15:0]),
	.Co(Tile_X2Y5_Co[0:0]),
	.E1BEG(Tile_X2Y5_E1BEG[3:0]),
	.E2BEG(Tile_X2Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y5_E6BEG[11:0]),
	.S1BEG(Tile_X2Y5_S1BEG[3:0]),
	.S2BEG(Tile_X2Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y5_W1BEG[3:0]),
	.W2BEG(Tile_X2Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y5_FrameData_O), 
	.FrameData_O(Tile_X2Y5_FrameData_O), 
	.FrameStrobe(Tile_X2Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y5_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y5_LUT4AB (
	.N1END(Tile_X3Y6_N1BEG[3:0]),
	.N2MID(Tile_X3Y6_N2BEG[7:0]),
	.N2END(Tile_X3Y6_N2BEGb[7:0]),
	.N4END(Tile_X3Y6_N4BEG[15:0]),
	.NN4END(Tile_X3Y6_NN4BEG[15:0]),
	.Ci(Tile_X3Y6_Co[0:0]),
	.E1END(Tile_X2Y5_E1BEG[3:0]),
	.E2MID(Tile_X2Y5_E2BEG[7:0]),
	.E2END(Tile_X2Y5_E2BEGb[7:0]),
	.EE4END(Tile_X2Y5_EE4BEG[15:0]),
	.E6END(Tile_X2Y5_E6BEG[11:0]),
	.S1END(Tile_X3Y4_S1BEG[3:0]),
	.S2MID(Tile_X3Y4_S2BEG[7:0]),
	.S2END(Tile_X3Y4_S2BEGb[7:0]),
	.S4END(Tile_X3Y4_S4BEG[15:0]),
	.SS4END(Tile_X3Y4_SS4BEG[15:0]),
	.W1END(Tile_X4Y5_W1BEG[3:0]),
	.W2MID(Tile_X4Y5_W2BEG[7:0]),
	.W2END(Tile_X4Y5_W2BEGb[7:0]),
	.WW4END(Tile_X4Y5_WW4BEG[15:0]),
	.W6END(Tile_X4Y5_W6BEG[11:0]),
	.N1BEG(Tile_X3Y5_N1BEG[3:0]),
	.N2BEG(Tile_X3Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y5_NN4BEG[15:0]),
	.Co(Tile_X3Y5_Co[0:0]),
	.E1BEG(Tile_X3Y5_E1BEG[3:0]),
	.E2BEG(Tile_X3Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y5_E6BEG[11:0]),
	.S1BEG(Tile_X3Y5_S1BEG[3:0]),
	.S2BEG(Tile_X3Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y5_W1BEG[3:0]),
	.W2BEG(Tile_X3Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y5_FrameData_O), 
	.FrameData_O(Tile_X3Y5_FrameData_O), 
	.FrameStrobe(Tile_X3Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y5_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y5_LUT4AB (
	.N1END(Tile_X4Y6_N1BEG[3:0]),
	.N2MID(Tile_X4Y6_N2BEG[7:0]),
	.N2END(Tile_X4Y6_N2BEGb[7:0]),
	.N4END(Tile_X4Y6_N4BEG[15:0]),
	.NN4END(Tile_X4Y6_NN4BEG[15:0]),
	.Ci(Tile_X4Y6_Co[0:0]),
	.E1END(Tile_X3Y5_E1BEG[3:0]),
	.E2MID(Tile_X3Y5_E2BEG[7:0]),
	.E2END(Tile_X3Y5_E2BEGb[7:0]),
	.EE4END(Tile_X3Y5_EE4BEG[15:0]),
	.E6END(Tile_X3Y5_E6BEG[11:0]),
	.S1END(Tile_X4Y4_S1BEG[3:0]),
	.S2MID(Tile_X4Y4_S2BEG[7:0]),
	.S2END(Tile_X4Y4_S2BEGb[7:0]),
	.S4END(Tile_X4Y4_S4BEG[15:0]),
	.SS4END(Tile_X4Y4_SS4BEG[15:0]),
	.W1END(Tile_X5Y5_W1BEG[3:0]),
	.W2MID(Tile_X5Y5_W2BEG[7:0]),
	.W2END(Tile_X5Y5_W2BEGb[7:0]),
	.WW4END(Tile_X5Y5_WW4BEG[15:0]),
	.W6END(Tile_X5Y5_W6BEG[11:0]),
	.N1BEG(Tile_X4Y5_N1BEG[3:0]),
	.N2BEG(Tile_X4Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y5_NN4BEG[15:0]),
	.Co(Tile_X4Y5_Co[0:0]),
	.E1BEG(Tile_X4Y5_E1BEG[3:0]),
	.E2BEG(Tile_X4Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y5_E6BEG[11:0]),
	.S1BEG(Tile_X4Y5_S1BEG[3:0]),
	.S2BEG(Tile_X4Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y5_W1BEG[3:0]),
	.W2BEG(Tile_X4Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y5_FrameData_O), 
	.FrameData_O(Tile_X4Y5_FrameData_O), 
	.FrameStrobe(Tile_X4Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y5_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y5_LUT4AB (
	.N1END(Tile_X6Y6_N1BEG[3:0]),
	.N2MID(Tile_X6Y6_N2BEG[7:0]),
	.N2END(Tile_X6Y6_N2BEGb[7:0]),
	.N4END(Tile_X6Y6_N4BEG[15:0]),
	.NN4END(Tile_X6Y6_NN4BEG[15:0]),
	.Ci(Tile_X6Y6_Co[0:0]),
	.E1END(Tile_X5Y5_E1BEG[3:0]),
	.E2MID(Tile_X5Y5_E2BEG[7:0]),
	.E2END(Tile_X5Y5_E2BEGb[7:0]),
	.EE4END(Tile_X5Y5_EE4BEG[15:0]),
	.E6END(Tile_X5Y5_E6BEG[11:0]),
	.S1END(Tile_X6Y4_S1BEG[3:0]),
	.S2MID(Tile_X6Y4_S2BEG[7:0]),
	.S2END(Tile_X6Y4_S2BEGb[7:0]),
	.S4END(Tile_X6Y4_S4BEG[15:0]),
	.SS4END(Tile_X6Y4_SS4BEG[15:0]),
	.W1END(Tile_X7Y5_W1BEG[3:0]),
	.W2MID(Tile_X7Y5_W2BEG[7:0]),
	.W2END(Tile_X7Y5_W2BEGb[7:0]),
	.WW4END(Tile_X7Y5_WW4BEG[15:0]),
	.W6END(Tile_X7Y5_W6BEG[11:0]),
	.N1BEG(Tile_X6Y5_N1BEG[3:0]),
	.N2BEG(Tile_X6Y5_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y5_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y5_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y5_NN4BEG[15:0]),
	.Co(Tile_X6Y5_Co[0:0]),
	.E1BEG(Tile_X6Y5_E1BEG[3:0]),
	.E2BEG(Tile_X6Y5_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y5_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y5_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y5_E6BEG[11:0]),
	.S1BEG(Tile_X6Y5_S1BEG[3:0]),
	.S2BEG(Tile_X6Y5_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y5_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y5_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y5_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y5_W1BEG[3:0]),
	.W2BEG(Tile_X6Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y5_FrameData_O), 
	.FrameData_O(Tile_X6Y5_FrameData_O), 
	.FrameStrobe(Tile_X6Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y5_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y5_E_CPU_IO (
	.E1END(Tile_X6Y5_E1BEG[3:0]),
	.E2MID(Tile_X6Y5_E2BEG[7:0]),
	.E2END(Tile_X6Y5_E2BEGb[7:0]),
	.EE4END(Tile_X6Y5_EE4BEG[15:0]),
	.E6END(Tile_X6Y5_E6BEG[11:0]),
	.W1BEG(Tile_X7Y5_W1BEG[3:0]),
	.W2BEG(Tile_X7Y5_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y5_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y5_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y5_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y5_OPA_I0),
	.OPA_I1(Tile_X7Y5_OPA_I1),
	.OPA_I2(Tile_X7Y5_OPA_I2),
	.OPA_I3(Tile_X7Y5_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y5_OPB_I0),
	.OPB_I1(Tile_X7Y5_OPB_I1),
	.OPB_I2(Tile_X7Y5_OPB_I2),
	.OPB_I3(Tile_X7Y5_OPB_I3),
	.RES0_O0(Tile_X7Y5_RES0_O0),
	.RES0_O1(Tile_X7Y5_RES0_O1),
	.RES0_O2(Tile_X7Y5_RES0_O2),
	.RES0_O3(Tile_X7Y5_RES0_O3),
	.RES1_O0(Tile_X7Y5_RES1_O0),
	.RES1_O1(Tile_X7Y5_RES1_O1),
	.RES1_O2(Tile_X7Y5_RES1_O2),
	.RES1_O3(Tile_X7Y5_RES1_O3),
	.RES2_O0(Tile_X7Y5_RES2_O0),
	.RES2_O1(Tile_X7Y5_RES2_O1),
	.RES2_O2(Tile_X7Y5_RES2_O2),
	.RES2_O3(Tile_X7Y5_RES2_O3),
	.FrameData(Tile_X6Y5_FrameData_O), 
	.FrameData_O(Tile_X7Y5_FrameData_O), 
	.FrameStrobe(Tile_X7Y6_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y5_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y6_W_CPU_IO (
	.W1END(Tile_X1Y6_W1BEG[3:0]),
	.W2MID(Tile_X1Y6_W2BEG[7:0]),
	.W2END(Tile_X1Y6_W2BEGb[7:0]),
	.WW4END(Tile_X1Y6_WW4BEG[15:0]),
	.W6END(Tile_X1Y6_W6BEG[11:0]),
	.E1BEG(Tile_X0Y6_E1BEG[3:0]),
	.E2BEG(Tile_X0Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y6_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y6_OPA_I0),
	.OPA_I1(Tile_X0Y6_OPA_I1),
	.OPA_I2(Tile_X0Y6_OPA_I2),
	.OPA_I3(Tile_X0Y6_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y6_OPB_I0),
	.OPB_I1(Tile_X0Y6_OPB_I1),
	.OPB_I2(Tile_X0Y6_OPB_I2),
	.OPB_I3(Tile_X0Y6_OPB_I3),
	.RES0_O0(Tile_X0Y6_RES0_O0),
	.RES0_O1(Tile_X0Y6_RES0_O1),
	.RES0_O2(Tile_X0Y6_RES0_O2),
	.RES0_O3(Tile_X0Y6_RES0_O3),
	.RES1_O0(Tile_X0Y6_RES1_O0),
	.RES1_O1(Tile_X0Y6_RES1_O1),
	.RES1_O2(Tile_X0Y6_RES1_O2),
	.RES1_O3(Tile_X0Y6_RES1_O3),
	.RES2_O0(Tile_X0Y6_RES2_O0),
	.RES2_O1(Tile_X0Y6_RES2_O1),
	.RES2_O2(Tile_X0Y6_RES2_O2),
	.RES2_O3(Tile_X0Y6_RES2_O3),
	.FrameData(Tile_Y6_FrameData), 
	.FrameData_O(Tile_X0Y6_FrameData_O), 
	.FrameStrobe(Tile_X0Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y6_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y6_LUT4AB (
	.N1END(Tile_X2Y7_N1BEG[3:0]),
	.N2MID(Tile_X2Y7_N2BEG[7:0]),
	.N2END(Tile_X2Y7_N2BEGb[7:0]),
	.N4END(Tile_X2Y7_N4BEG[15:0]),
	.NN4END(Tile_X2Y7_NN4BEG[15:0]),
	.Ci(Tile_X2Y7_Co[0:0]),
	.E1END(Tile_X1Y6_E1BEG[3:0]),
	.E2MID(Tile_X1Y6_E2BEG[7:0]),
	.E2END(Tile_X1Y6_E2BEGb[7:0]),
	.EE4END(Tile_X1Y6_EE4BEG[15:0]),
	.E6END(Tile_X1Y6_E6BEG[11:0]),
	.S1END(Tile_X2Y5_S1BEG[3:0]),
	.S2MID(Tile_X2Y5_S2BEG[7:0]),
	.S2END(Tile_X2Y5_S2BEGb[7:0]),
	.S4END(Tile_X2Y5_S4BEG[15:0]),
	.SS4END(Tile_X2Y5_SS4BEG[15:0]),
	.W1END(Tile_X3Y6_W1BEG[3:0]),
	.W2MID(Tile_X3Y6_W2BEG[7:0]),
	.W2END(Tile_X3Y6_W2BEGb[7:0]),
	.WW4END(Tile_X3Y6_WW4BEG[15:0]),
	.W6END(Tile_X3Y6_W6BEG[11:0]),
	.N1BEG(Tile_X2Y6_N1BEG[3:0]),
	.N2BEG(Tile_X2Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y6_NN4BEG[15:0]),
	.Co(Tile_X2Y6_Co[0:0]),
	.E1BEG(Tile_X2Y6_E1BEG[3:0]),
	.E2BEG(Tile_X2Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y6_E6BEG[11:0]),
	.S1BEG(Tile_X2Y6_S1BEG[3:0]),
	.S2BEG(Tile_X2Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y6_W1BEG[3:0]),
	.W2BEG(Tile_X2Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y6_FrameData_O), 
	.FrameData_O(Tile_X2Y6_FrameData_O), 
	.FrameStrobe(Tile_X2Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y6_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y6_LUT4AB (
	.N1END(Tile_X3Y7_N1BEG[3:0]),
	.N2MID(Tile_X3Y7_N2BEG[7:0]),
	.N2END(Tile_X3Y7_N2BEGb[7:0]),
	.N4END(Tile_X3Y7_N4BEG[15:0]),
	.NN4END(Tile_X3Y7_NN4BEG[15:0]),
	.Ci(Tile_X3Y7_Co[0:0]),
	.E1END(Tile_X2Y6_E1BEG[3:0]),
	.E2MID(Tile_X2Y6_E2BEG[7:0]),
	.E2END(Tile_X2Y6_E2BEGb[7:0]),
	.EE4END(Tile_X2Y6_EE4BEG[15:0]),
	.E6END(Tile_X2Y6_E6BEG[11:0]),
	.S1END(Tile_X3Y5_S1BEG[3:0]),
	.S2MID(Tile_X3Y5_S2BEG[7:0]),
	.S2END(Tile_X3Y5_S2BEGb[7:0]),
	.S4END(Tile_X3Y5_S4BEG[15:0]),
	.SS4END(Tile_X3Y5_SS4BEG[15:0]),
	.W1END(Tile_X4Y6_W1BEG[3:0]),
	.W2MID(Tile_X4Y6_W2BEG[7:0]),
	.W2END(Tile_X4Y6_W2BEGb[7:0]),
	.WW4END(Tile_X4Y6_WW4BEG[15:0]),
	.W6END(Tile_X4Y6_W6BEG[11:0]),
	.N1BEG(Tile_X3Y6_N1BEG[3:0]),
	.N2BEG(Tile_X3Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y6_NN4BEG[15:0]),
	.Co(Tile_X3Y6_Co[0:0]),
	.E1BEG(Tile_X3Y6_E1BEG[3:0]),
	.E2BEG(Tile_X3Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y6_E6BEG[11:0]),
	.S1BEG(Tile_X3Y6_S1BEG[3:0]),
	.S2BEG(Tile_X3Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y6_W1BEG[3:0]),
	.W2BEG(Tile_X3Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y6_FrameData_O), 
	.FrameData_O(Tile_X3Y6_FrameData_O), 
	.FrameStrobe(Tile_X3Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y6_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y6_LUT4AB (
	.N1END(Tile_X4Y7_N1BEG[3:0]),
	.N2MID(Tile_X4Y7_N2BEG[7:0]),
	.N2END(Tile_X4Y7_N2BEGb[7:0]),
	.N4END(Tile_X4Y7_N4BEG[15:0]),
	.NN4END(Tile_X4Y7_NN4BEG[15:0]),
	.Ci(Tile_X4Y7_Co[0:0]),
	.E1END(Tile_X3Y6_E1BEG[3:0]),
	.E2MID(Tile_X3Y6_E2BEG[7:0]),
	.E2END(Tile_X3Y6_E2BEGb[7:0]),
	.EE4END(Tile_X3Y6_EE4BEG[15:0]),
	.E6END(Tile_X3Y6_E6BEG[11:0]),
	.S1END(Tile_X4Y5_S1BEG[3:0]),
	.S2MID(Tile_X4Y5_S2BEG[7:0]),
	.S2END(Tile_X4Y5_S2BEGb[7:0]),
	.S4END(Tile_X4Y5_S4BEG[15:0]),
	.SS4END(Tile_X4Y5_SS4BEG[15:0]),
	.W1END(Tile_X5Y6_W1BEG[3:0]),
	.W2MID(Tile_X5Y6_W2BEG[7:0]),
	.W2END(Tile_X5Y6_W2BEGb[7:0]),
	.WW4END(Tile_X5Y6_WW4BEG[15:0]),
	.W6END(Tile_X5Y6_W6BEG[11:0]),
	.N1BEG(Tile_X4Y6_N1BEG[3:0]),
	.N2BEG(Tile_X4Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y6_NN4BEG[15:0]),
	.Co(Tile_X4Y6_Co[0:0]),
	.E1BEG(Tile_X4Y6_E1BEG[3:0]),
	.E2BEG(Tile_X4Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y6_E6BEG[11:0]),
	.S1BEG(Tile_X4Y6_S1BEG[3:0]),
	.S2BEG(Tile_X4Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y6_W1BEG[3:0]),
	.W2BEG(Tile_X4Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y6_FrameData_O), 
	.FrameData_O(Tile_X4Y6_FrameData_O), 
	.FrameStrobe(Tile_X4Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y6_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y6_LUT4AB (
	.N1END(Tile_X6Y7_N1BEG[3:0]),
	.N2MID(Tile_X6Y7_N2BEG[7:0]),
	.N2END(Tile_X6Y7_N2BEGb[7:0]),
	.N4END(Tile_X6Y7_N4BEG[15:0]),
	.NN4END(Tile_X6Y7_NN4BEG[15:0]),
	.Ci(Tile_X6Y7_Co[0:0]),
	.E1END(Tile_X5Y6_E1BEG[3:0]),
	.E2MID(Tile_X5Y6_E2BEG[7:0]),
	.E2END(Tile_X5Y6_E2BEGb[7:0]),
	.EE4END(Tile_X5Y6_EE4BEG[15:0]),
	.E6END(Tile_X5Y6_E6BEG[11:0]),
	.S1END(Tile_X6Y5_S1BEG[3:0]),
	.S2MID(Tile_X6Y5_S2BEG[7:0]),
	.S2END(Tile_X6Y5_S2BEGb[7:0]),
	.S4END(Tile_X6Y5_S4BEG[15:0]),
	.SS4END(Tile_X6Y5_SS4BEG[15:0]),
	.W1END(Tile_X7Y6_W1BEG[3:0]),
	.W2MID(Tile_X7Y6_W2BEG[7:0]),
	.W2END(Tile_X7Y6_W2BEGb[7:0]),
	.WW4END(Tile_X7Y6_WW4BEG[15:0]),
	.W6END(Tile_X7Y6_W6BEG[11:0]),
	.N1BEG(Tile_X6Y6_N1BEG[3:0]),
	.N2BEG(Tile_X6Y6_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y6_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y6_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y6_NN4BEG[15:0]),
	.Co(Tile_X6Y6_Co[0:0]),
	.E1BEG(Tile_X6Y6_E1BEG[3:0]),
	.E2BEG(Tile_X6Y6_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y6_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y6_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y6_E6BEG[11:0]),
	.S1BEG(Tile_X6Y6_S1BEG[3:0]),
	.S2BEG(Tile_X6Y6_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y6_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y6_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y6_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y6_W1BEG[3:0]),
	.W2BEG(Tile_X6Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y6_FrameData_O), 
	.FrameData_O(Tile_X6Y6_FrameData_O), 
	.FrameStrobe(Tile_X6Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y6_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y6_E_CPU_IO (
	.E1END(Tile_X6Y6_E1BEG[3:0]),
	.E2MID(Tile_X6Y6_E2BEG[7:0]),
	.E2END(Tile_X6Y6_E2BEGb[7:0]),
	.EE4END(Tile_X6Y6_EE4BEG[15:0]),
	.E6END(Tile_X6Y6_E6BEG[11:0]),
	.W1BEG(Tile_X7Y6_W1BEG[3:0]),
	.W2BEG(Tile_X7Y6_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y6_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y6_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y6_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y6_OPA_I0),
	.OPA_I1(Tile_X7Y6_OPA_I1),
	.OPA_I2(Tile_X7Y6_OPA_I2),
	.OPA_I3(Tile_X7Y6_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y6_OPB_I0),
	.OPB_I1(Tile_X7Y6_OPB_I1),
	.OPB_I2(Tile_X7Y6_OPB_I2),
	.OPB_I3(Tile_X7Y6_OPB_I3),
	.RES0_O0(Tile_X7Y6_RES0_O0),
	.RES0_O1(Tile_X7Y6_RES0_O1),
	.RES0_O2(Tile_X7Y6_RES0_O2),
	.RES0_O3(Tile_X7Y6_RES0_O3),
	.RES1_O0(Tile_X7Y6_RES1_O0),
	.RES1_O1(Tile_X7Y6_RES1_O1),
	.RES1_O2(Tile_X7Y6_RES1_O2),
	.RES1_O3(Tile_X7Y6_RES1_O3),
	.RES2_O0(Tile_X7Y6_RES2_O0),
	.RES2_O1(Tile_X7Y6_RES2_O1),
	.RES2_O2(Tile_X7Y6_RES2_O2),
	.RES2_O3(Tile_X7Y6_RES2_O3),
	.FrameData(Tile_X6Y6_FrameData_O), 
	.FrameData_O(Tile_X7Y6_FrameData_O), 
	.FrameStrobe(Tile_X7Y7_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y6_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y7_W_CPU_IO (
	.W1END(Tile_X1Y7_W1BEG[3:0]),
	.W2MID(Tile_X1Y7_W2BEG[7:0]),
	.W2END(Tile_X1Y7_W2BEGb[7:0]),
	.WW4END(Tile_X1Y7_WW4BEG[15:0]),
	.W6END(Tile_X1Y7_W6BEG[11:0]),
	.E1BEG(Tile_X0Y7_E1BEG[3:0]),
	.E2BEG(Tile_X0Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y7_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y7_OPA_I0),
	.OPA_I1(Tile_X0Y7_OPA_I1),
	.OPA_I2(Tile_X0Y7_OPA_I2),
	.OPA_I3(Tile_X0Y7_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y7_OPB_I0),
	.OPB_I1(Tile_X0Y7_OPB_I1),
	.OPB_I2(Tile_X0Y7_OPB_I2),
	.OPB_I3(Tile_X0Y7_OPB_I3),
	.RES0_O0(Tile_X0Y7_RES0_O0),
	.RES0_O1(Tile_X0Y7_RES0_O1),
	.RES0_O2(Tile_X0Y7_RES0_O2),
	.RES0_O3(Tile_X0Y7_RES0_O3),
	.RES1_O0(Tile_X0Y7_RES1_O0),
	.RES1_O1(Tile_X0Y7_RES1_O1),
	.RES1_O2(Tile_X0Y7_RES1_O2),
	.RES1_O3(Tile_X0Y7_RES1_O3),
	.RES2_O0(Tile_X0Y7_RES2_O0),
	.RES2_O1(Tile_X0Y7_RES2_O1),
	.RES2_O2(Tile_X0Y7_RES2_O2),
	.RES2_O3(Tile_X0Y7_RES2_O3),
	.FrameData(Tile_Y7_FrameData), 
	.FrameData_O(Tile_X0Y7_FrameData_O), 
	.FrameStrobe(Tile_X0Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y7_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y7_LUT4AB (
	.N1END(Tile_X2Y8_N1BEG[3:0]),
	.N2MID(Tile_X2Y8_N2BEG[7:0]),
	.N2END(Tile_X2Y8_N2BEGb[7:0]),
	.N4END(Tile_X2Y8_N4BEG[15:0]),
	.NN4END(Tile_X2Y8_NN4BEG[15:0]),
	.Ci(Tile_X2Y8_Co[0:0]),
	.E1END(Tile_X1Y7_E1BEG[3:0]),
	.E2MID(Tile_X1Y7_E2BEG[7:0]),
	.E2END(Tile_X1Y7_E2BEGb[7:0]),
	.EE4END(Tile_X1Y7_EE4BEG[15:0]),
	.E6END(Tile_X1Y7_E6BEG[11:0]),
	.S1END(Tile_X2Y6_S1BEG[3:0]),
	.S2MID(Tile_X2Y6_S2BEG[7:0]),
	.S2END(Tile_X2Y6_S2BEGb[7:0]),
	.S4END(Tile_X2Y6_S4BEG[15:0]),
	.SS4END(Tile_X2Y6_SS4BEG[15:0]),
	.W1END(Tile_X3Y7_W1BEG[3:0]),
	.W2MID(Tile_X3Y7_W2BEG[7:0]),
	.W2END(Tile_X3Y7_W2BEGb[7:0]),
	.WW4END(Tile_X3Y7_WW4BEG[15:0]),
	.W6END(Tile_X3Y7_W6BEG[11:0]),
	.N1BEG(Tile_X2Y7_N1BEG[3:0]),
	.N2BEG(Tile_X2Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y7_NN4BEG[15:0]),
	.Co(Tile_X2Y7_Co[0:0]),
	.E1BEG(Tile_X2Y7_E1BEG[3:0]),
	.E2BEG(Tile_X2Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y7_E6BEG[11:0]),
	.S1BEG(Tile_X2Y7_S1BEG[3:0]),
	.S2BEG(Tile_X2Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y7_W1BEG[3:0]),
	.W2BEG(Tile_X2Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y7_FrameData_O), 
	.FrameData_O(Tile_X2Y7_FrameData_O), 
	.FrameStrobe(Tile_X2Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y7_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y7_LUT4AB (
	.N1END(Tile_X3Y8_N1BEG[3:0]),
	.N2MID(Tile_X3Y8_N2BEG[7:0]),
	.N2END(Tile_X3Y8_N2BEGb[7:0]),
	.N4END(Tile_X3Y8_N4BEG[15:0]),
	.NN4END(Tile_X3Y8_NN4BEG[15:0]),
	.Ci(Tile_X3Y8_Co[0:0]),
	.E1END(Tile_X2Y7_E1BEG[3:0]),
	.E2MID(Tile_X2Y7_E2BEG[7:0]),
	.E2END(Tile_X2Y7_E2BEGb[7:0]),
	.EE4END(Tile_X2Y7_EE4BEG[15:0]),
	.E6END(Tile_X2Y7_E6BEG[11:0]),
	.S1END(Tile_X3Y6_S1BEG[3:0]),
	.S2MID(Tile_X3Y6_S2BEG[7:0]),
	.S2END(Tile_X3Y6_S2BEGb[7:0]),
	.S4END(Tile_X3Y6_S4BEG[15:0]),
	.SS4END(Tile_X3Y6_SS4BEG[15:0]),
	.W1END(Tile_X4Y7_W1BEG[3:0]),
	.W2MID(Tile_X4Y7_W2BEG[7:0]),
	.W2END(Tile_X4Y7_W2BEGb[7:0]),
	.WW4END(Tile_X4Y7_WW4BEG[15:0]),
	.W6END(Tile_X4Y7_W6BEG[11:0]),
	.N1BEG(Tile_X3Y7_N1BEG[3:0]),
	.N2BEG(Tile_X3Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y7_NN4BEG[15:0]),
	.Co(Tile_X3Y7_Co[0:0]),
	.E1BEG(Tile_X3Y7_E1BEG[3:0]),
	.E2BEG(Tile_X3Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y7_E6BEG[11:0]),
	.S1BEG(Tile_X3Y7_S1BEG[3:0]),
	.S2BEG(Tile_X3Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y7_W1BEG[3:0]),
	.W2BEG(Tile_X3Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y7_FrameData_O), 
	.FrameData_O(Tile_X3Y7_FrameData_O), 
	.FrameStrobe(Tile_X3Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y7_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y7_LUT4AB (
	.N1END(Tile_X4Y8_N1BEG[3:0]),
	.N2MID(Tile_X4Y8_N2BEG[7:0]),
	.N2END(Tile_X4Y8_N2BEGb[7:0]),
	.N4END(Tile_X4Y8_N4BEG[15:0]),
	.NN4END(Tile_X4Y8_NN4BEG[15:0]),
	.Ci(Tile_X4Y8_Co[0:0]),
	.E1END(Tile_X3Y7_E1BEG[3:0]),
	.E2MID(Tile_X3Y7_E2BEG[7:0]),
	.E2END(Tile_X3Y7_E2BEGb[7:0]),
	.EE4END(Tile_X3Y7_EE4BEG[15:0]),
	.E6END(Tile_X3Y7_E6BEG[11:0]),
	.S1END(Tile_X4Y6_S1BEG[3:0]),
	.S2MID(Tile_X4Y6_S2BEG[7:0]),
	.S2END(Tile_X4Y6_S2BEGb[7:0]),
	.S4END(Tile_X4Y6_S4BEG[15:0]),
	.SS4END(Tile_X4Y6_SS4BEG[15:0]),
	.W1END(Tile_X5Y7_W1BEG[3:0]),
	.W2MID(Tile_X5Y7_W2BEG[7:0]),
	.W2END(Tile_X5Y7_W2BEGb[7:0]),
	.WW4END(Tile_X5Y7_WW4BEG[15:0]),
	.W6END(Tile_X5Y7_W6BEG[11:0]),
	.N1BEG(Tile_X4Y7_N1BEG[3:0]),
	.N2BEG(Tile_X4Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y7_NN4BEG[15:0]),
	.Co(Tile_X4Y7_Co[0:0]),
	.E1BEG(Tile_X4Y7_E1BEG[3:0]),
	.E2BEG(Tile_X4Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y7_E6BEG[11:0]),
	.S1BEG(Tile_X4Y7_S1BEG[3:0]),
	.S2BEG(Tile_X4Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y7_W1BEG[3:0]),
	.W2BEG(Tile_X4Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y7_FrameData_O), 
	.FrameData_O(Tile_X4Y7_FrameData_O), 
	.FrameStrobe(Tile_X4Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y7_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y7_LUT4AB (
	.N1END(Tile_X6Y8_N1BEG[3:0]),
	.N2MID(Tile_X6Y8_N2BEG[7:0]),
	.N2END(Tile_X6Y8_N2BEGb[7:0]),
	.N4END(Tile_X6Y8_N4BEG[15:0]),
	.NN4END(Tile_X6Y8_NN4BEG[15:0]),
	.Ci(Tile_X6Y8_Co[0:0]),
	.E1END(Tile_X5Y7_E1BEG[3:0]),
	.E2MID(Tile_X5Y7_E2BEG[7:0]),
	.E2END(Tile_X5Y7_E2BEGb[7:0]),
	.EE4END(Tile_X5Y7_EE4BEG[15:0]),
	.E6END(Tile_X5Y7_E6BEG[11:0]),
	.S1END(Tile_X6Y6_S1BEG[3:0]),
	.S2MID(Tile_X6Y6_S2BEG[7:0]),
	.S2END(Tile_X6Y6_S2BEGb[7:0]),
	.S4END(Tile_X6Y6_S4BEG[15:0]),
	.SS4END(Tile_X6Y6_SS4BEG[15:0]),
	.W1END(Tile_X7Y7_W1BEG[3:0]),
	.W2MID(Tile_X7Y7_W2BEG[7:0]),
	.W2END(Tile_X7Y7_W2BEGb[7:0]),
	.WW4END(Tile_X7Y7_WW4BEG[15:0]),
	.W6END(Tile_X7Y7_W6BEG[11:0]),
	.N1BEG(Tile_X6Y7_N1BEG[3:0]),
	.N2BEG(Tile_X6Y7_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y7_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y7_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y7_NN4BEG[15:0]),
	.Co(Tile_X6Y7_Co[0:0]),
	.E1BEG(Tile_X6Y7_E1BEG[3:0]),
	.E2BEG(Tile_X6Y7_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y7_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y7_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y7_E6BEG[11:0]),
	.S1BEG(Tile_X6Y7_S1BEG[3:0]),
	.S2BEG(Tile_X6Y7_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y7_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y7_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y7_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y7_W1BEG[3:0]),
	.W2BEG(Tile_X6Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y7_FrameData_O), 
	.FrameData_O(Tile_X6Y7_FrameData_O), 
	.FrameStrobe(Tile_X6Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y7_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y7_E_CPU_IO (
	.E1END(Tile_X6Y7_E1BEG[3:0]),
	.E2MID(Tile_X6Y7_E2BEG[7:0]),
	.E2END(Tile_X6Y7_E2BEGb[7:0]),
	.EE4END(Tile_X6Y7_EE4BEG[15:0]),
	.E6END(Tile_X6Y7_E6BEG[11:0]),
	.W1BEG(Tile_X7Y7_W1BEG[3:0]),
	.W2BEG(Tile_X7Y7_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y7_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y7_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y7_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y7_OPA_I0),
	.OPA_I1(Tile_X7Y7_OPA_I1),
	.OPA_I2(Tile_X7Y7_OPA_I2),
	.OPA_I3(Tile_X7Y7_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y7_OPB_I0),
	.OPB_I1(Tile_X7Y7_OPB_I1),
	.OPB_I2(Tile_X7Y7_OPB_I2),
	.OPB_I3(Tile_X7Y7_OPB_I3),
	.RES0_O0(Tile_X7Y7_RES0_O0),
	.RES0_O1(Tile_X7Y7_RES0_O1),
	.RES0_O2(Tile_X7Y7_RES0_O2),
	.RES0_O3(Tile_X7Y7_RES0_O3),
	.RES1_O0(Tile_X7Y7_RES1_O0),
	.RES1_O1(Tile_X7Y7_RES1_O1),
	.RES1_O2(Tile_X7Y7_RES1_O2),
	.RES1_O3(Tile_X7Y7_RES1_O3),
	.RES2_O0(Tile_X7Y7_RES2_O0),
	.RES2_O1(Tile_X7Y7_RES2_O1),
	.RES2_O2(Tile_X7Y7_RES2_O2),
	.RES2_O3(Tile_X7Y7_RES2_O3),
	.FrameData(Tile_X6Y7_FrameData_O), 
	.FrameData_O(Tile_X7Y7_FrameData_O), 
	.FrameStrobe(Tile_X7Y8_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y7_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y8_W_CPU_IO (
	.W1END(Tile_X1Y8_W1BEG[3:0]),
	.W2MID(Tile_X1Y8_W2BEG[7:0]),
	.W2END(Tile_X1Y8_W2BEGb[7:0]),
	.WW4END(Tile_X1Y8_WW4BEG[15:0]),
	.W6END(Tile_X1Y8_W6BEG[11:0]),
	.E1BEG(Tile_X0Y8_E1BEG[3:0]),
	.E2BEG(Tile_X0Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y8_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y8_OPA_I0),
	.OPA_I1(Tile_X0Y8_OPA_I1),
	.OPA_I2(Tile_X0Y8_OPA_I2),
	.OPA_I3(Tile_X0Y8_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y8_OPB_I0),
	.OPB_I1(Tile_X0Y8_OPB_I1),
	.OPB_I2(Tile_X0Y8_OPB_I2),
	.OPB_I3(Tile_X0Y8_OPB_I3),
	.RES0_O0(Tile_X0Y8_RES0_O0),
	.RES0_O1(Tile_X0Y8_RES0_O1),
	.RES0_O2(Tile_X0Y8_RES0_O2),
	.RES0_O3(Tile_X0Y8_RES0_O3),
	.RES1_O0(Tile_X0Y8_RES1_O0),
	.RES1_O1(Tile_X0Y8_RES1_O1),
	.RES1_O2(Tile_X0Y8_RES1_O2),
	.RES1_O3(Tile_X0Y8_RES1_O3),
	.RES2_O0(Tile_X0Y8_RES2_O0),
	.RES2_O1(Tile_X0Y8_RES2_O1),
	.RES2_O2(Tile_X0Y8_RES2_O2),
	.RES2_O3(Tile_X0Y8_RES2_O3),
	.FrameData(Tile_Y8_FrameData), 
	.FrameData_O(Tile_X0Y8_FrameData_O), 
	.FrameStrobe(Tile_X0Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y8_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y8_LUT4AB (
	.N1END(Tile_X2Y9_N1BEG[3:0]),
	.N2MID(Tile_X2Y9_N2BEG[7:0]),
	.N2END(Tile_X2Y9_N2BEGb[7:0]),
	.N4END(Tile_X2Y9_N4BEG[15:0]),
	.NN4END(Tile_X2Y9_NN4BEG[15:0]),
	.Ci(Tile_X2Y9_Co[0:0]),
	.E1END(Tile_X1Y8_E1BEG[3:0]),
	.E2MID(Tile_X1Y8_E2BEG[7:0]),
	.E2END(Tile_X1Y8_E2BEGb[7:0]),
	.EE4END(Tile_X1Y8_EE4BEG[15:0]),
	.E6END(Tile_X1Y8_E6BEG[11:0]),
	.S1END(Tile_X2Y7_S1BEG[3:0]),
	.S2MID(Tile_X2Y7_S2BEG[7:0]),
	.S2END(Tile_X2Y7_S2BEGb[7:0]),
	.S4END(Tile_X2Y7_S4BEG[15:0]),
	.SS4END(Tile_X2Y7_SS4BEG[15:0]),
	.W1END(Tile_X3Y8_W1BEG[3:0]),
	.W2MID(Tile_X3Y8_W2BEG[7:0]),
	.W2END(Tile_X3Y8_W2BEGb[7:0]),
	.WW4END(Tile_X3Y8_WW4BEG[15:0]),
	.W6END(Tile_X3Y8_W6BEG[11:0]),
	.N1BEG(Tile_X2Y8_N1BEG[3:0]),
	.N2BEG(Tile_X2Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y8_NN4BEG[15:0]),
	.Co(Tile_X2Y8_Co[0:0]),
	.E1BEG(Tile_X2Y8_E1BEG[3:0]),
	.E2BEG(Tile_X2Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y8_E6BEG[11:0]),
	.S1BEG(Tile_X2Y8_S1BEG[3:0]),
	.S2BEG(Tile_X2Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y8_W1BEG[3:0]),
	.W2BEG(Tile_X2Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y8_FrameData_O), 
	.FrameData_O(Tile_X2Y8_FrameData_O), 
	.FrameStrobe(Tile_X2Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y8_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y8_LUT4AB (
	.N1END(Tile_X3Y9_N1BEG[3:0]),
	.N2MID(Tile_X3Y9_N2BEG[7:0]),
	.N2END(Tile_X3Y9_N2BEGb[7:0]),
	.N4END(Tile_X3Y9_N4BEG[15:0]),
	.NN4END(Tile_X3Y9_NN4BEG[15:0]),
	.Ci(Tile_X3Y9_Co[0:0]),
	.E1END(Tile_X2Y8_E1BEG[3:0]),
	.E2MID(Tile_X2Y8_E2BEG[7:0]),
	.E2END(Tile_X2Y8_E2BEGb[7:0]),
	.EE4END(Tile_X2Y8_EE4BEG[15:0]),
	.E6END(Tile_X2Y8_E6BEG[11:0]),
	.S1END(Tile_X3Y7_S1BEG[3:0]),
	.S2MID(Tile_X3Y7_S2BEG[7:0]),
	.S2END(Tile_X3Y7_S2BEGb[7:0]),
	.S4END(Tile_X3Y7_S4BEG[15:0]),
	.SS4END(Tile_X3Y7_SS4BEG[15:0]),
	.W1END(Tile_X4Y8_W1BEG[3:0]),
	.W2MID(Tile_X4Y8_W2BEG[7:0]),
	.W2END(Tile_X4Y8_W2BEGb[7:0]),
	.WW4END(Tile_X4Y8_WW4BEG[15:0]),
	.W6END(Tile_X4Y8_W6BEG[11:0]),
	.N1BEG(Tile_X3Y8_N1BEG[3:0]),
	.N2BEG(Tile_X3Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y8_NN4BEG[15:0]),
	.Co(Tile_X3Y8_Co[0:0]),
	.E1BEG(Tile_X3Y8_E1BEG[3:0]),
	.E2BEG(Tile_X3Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y8_E6BEG[11:0]),
	.S1BEG(Tile_X3Y8_S1BEG[3:0]),
	.S2BEG(Tile_X3Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y8_W1BEG[3:0]),
	.W2BEG(Tile_X3Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y8_FrameData_O), 
	.FrameData_O(Tile_X3Y8_FrameData_O), 
	.FrameStrobe(Tile_X3Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y8_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y8_LUT4AB (
	.N1END(Tile_X4Y9_N1BEG[3:0]),
	.N2MID(Tile_X4Y9_N2BEG[7:0]),
	.N2END(Tile_X4Y9_N2BEGb[7:0]),
	.N4END(Tile_X4Y9_N4BEG[15:0]),
	.NN4END(Tile_X4Y9_NN4BEG[15:0]),
	.Ci(Tile_X4Y9_Co[0:0]),
	.E1END(Tile_X3Y8_E1BEG[3:0]),
	.E2MID(Tile_X3Y8_E2BEG[7:0]),
	.E2END(Tile_X3Y8_E2BEGb[7:0]),
	.EE4END(Tile_X3Y8_EE4BEG[15:0]),
	.E6END(Tile_X3Y8_E6BEG[11:0]),
	.S1END(Tile_X4Y7_S1BEG[3:0]),
	.S2MID(Tile_X4Y7_S2BEG[7:0]),
	.S2END(Tile_X4Y7_S2BEGb[7:0]),
	.S4END(Tile_X4Y7_S4BEG[15:0]),
	.SS4END(Tile_X4Y7_SS4BEG[15:0]),
	.W1END(Tile_X5Y8_W1BEG[3:0]),
	.W2MID(Tile_X5Y8_W2BEG[7:0]),
	.W2END(Tile_X5Y8_W2BEGb[7:0]),
	.WW4END(Tile_X5Y8_WW4BEG[15:0]),
	.W6END(Tile_X5Y8_W6BEG[11:0]),
	.N1BEG(Tile_X4Y8_N1BEG[3:0]),
	.N2BEG(Tile_X4Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y8_NN4BEG[15:0]),
	.Co(Tile_X4Y8_Co[0:0]),
	.E1BEG(Tile_X4Y8_E1BEG[3:0]),
	.E2BEG(Tile_X4Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y8_E6BEG[11:0]),
	.S1BEG(Tile_X4Y8_S1BEG[3:0]),
	.S2BEG(Tile_X4Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y8_W1BEG[3:0]),
	.W2BEG(Tile_X4Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y8_FrameData_O), 
	.FrameData_O(Tile_X4Y8_FrameData_O), 
	.FrameStrobe(Tile_X4Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y8_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y8_LUT4AB (
	.N1END(Tile_X6Y9_N1BEG[3:0]),
	.N2MID(Tile_X6Y9_N2BEG[7:0]),
	.N2END(Tile_X6Y9_N2BEGb[7:0]),
	.N4END(Tile_X6Y9_N4BEG[15:0]),
	.NN4END(Tile_X6Y9_NN4BEG[15:0]),
	.Ci(Tile_X6Y9_Co[0:0]),
	.E1END(Tile_X5Y8_E1BEG[3:0]),
	.E2MID(Tile_X5Y8_E2BEG[7:0]),
	.E2END(Tile_X5Y8_E2BEGb[7:0]),
	.EE4END(Tile_X5Y8_EE4BEG[15:0]),
	.E6END(Tile_X5Y8_E6BEG[11:0]),
	.S1END(Tile_X6Y7_S1BEG[3:0]),
	.S2MID(Tile_X6Y7_S2BEG[7:0]),
	.S2END(Tile_X6Y7_S2BEGb[7:0]),
	.S4END(Tile_X6Y7_S4BEG[15:0]),
	.SS4END(Tile_X6Y7_SS4BEG[15:0]),
	.W1END(Tile_X7Y8_W1BEG[3:0]),
	.W2MID(Tile_X7Y8_W2BEG[7:0]),
	.W2END(Tile_X7Y8_W2BEGb[7:0]),
	.WW4END(Tile_X7Y8_WW4BEG[15:0]),
	.W6END(Tile_X7Y8_W6BEG[11:0]),
	.N1BEG(Tile_X6Y8_N1BEG[3:0]),
	.N2BEG(Tile_X6Y8_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y8_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y8_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y8_NN4BEG[15:0]),
	.Co(Tile_X6Y8_Co[0:0]),
	.E1BEG(Tile_X6Y8_E1BEG[3:0]),
	.E2BEG(Tile_X6Y8_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y8_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y8_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y8_E6BEG[11:0]),
	.S1BEG(Tile_X6Y8_S1BEG[3:0]),
	.S2BEG(Tile_X6Y8_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y8_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y8_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y8_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y8_W1BEG[3:0]),
	.W2BEG(Tile_X6Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y8_FrameData_O), 
	.FrameData_O(Tile_X6Y8_FrameData_O), 
	.FrameStrobe(Tile_X6Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y8_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y8_E_CPU_IO (
	.E1END(Tile_X6Y8_E1BEG[3:0]),
	.E2MID(Tile_X6Y8_E2BEG[7:0]),
	.E2END(Tile_X6Y8_E2BEGb[7:0]),
	.EE4END(Tile_X6Y8_EE4BEG[15:0]),
	.E6END(Tile_X6Y8_E6BEG[11:0]),
	.W1BEG(Tile_X7Y8_W1BEG[3:0]),
	.W2BEG(Tile_X7Y8_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y8_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y8_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y8_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y8_OPA_I0),
	.OPA_I1(Tile_X7Y8_OPA_I1),
	.OPA_I2(Tile_X7Y8_OPA_I2),
	.OPA_I3(Tile_X7Y8_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y8_OPB_I0),
	.OPB_I1(Tile_X7Y8_OPB_I1),
	.OPB_I2(Tile_X7Y8_OPB_I2),
	.OPB_I3(Tile_X7Y8_OPB_I3),
	.RES0_O0(Tile_X7Y8_RES0_O0),
	.RES0_O1(Tile_X7Y8_RES0_O1),
	.RES0_O2(Tile_X7Y8_RES0_O2),
	.RES0_O3(Tile_X7Y8_RES0_O3),
	.RES1_O0(Tile_X7Y8_RES1_O0),
	.RES1_O1(Tile_X7Y8_RES1_O1),
	.RES1_O2(Tile_X7Y8_RES1_O2),
	.RES1_O3(Tile_X7Y8_RES1_O3),
	.RES2_O0(Tile_X7Y8_RES2_O0),
	.RES2_O1(Tile_X7Y8_RES2_O1),
	.RES2_O2(Tile_X7Y8_RES2_O2),
	.RES2_O3(Tile_X7Y8_RES2_O3),
	.FrameData(Tile_X6Y8_FrameData_O), 
	.FrameData_O(Tile_X7Y8_FrameData_O), 
	.FrameStrobe(Tile_X7Y9_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y8_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y9_W_CPU_IO (
	.W1END(Tile_X1Y9_W1BEG[3:0]),
	.W2MID(Tile_X1Y9_W2BEG[7:0]),
	.W2END(Tile_X1Y9_W2BEGb[7:0]),
	.WW4END(Tile_X1Y9_WW4BEG[15:0]),
	.W6END(Tile_X1Y9_W6BEG[11:0]),
	.E1BEG(Tile_X0Y9_E1BEG[3:0]),
	.E2BEG(Tile_X0Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y9_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y9_OPA_I0),
	.OPA_I1(Tile_X0Y9_OPA_I1),
	.OPA_I2(Tile_X0Y9_OPA_I2),
	.OPA_I3(Tile_X0Y9_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y9_OPB_I0),
	.OPB_I1(Tile_X0Y9_OPB_I1),
	.OPB_I2(Tile_X0Y9_OPB_I2),
	.OPB_I3(Tile_X0Y9_OPB_I3),
	.RES0_O0(Tile_X0Y9_RES0_O0),
	.RES0_O1(Tile_X0Y9_RES0_O1),
	.RES0_O2(Tile_X0Y9_RES0_O2),
	.RES0_O3(Tile_X0Y9_RES0_O3),
	.RES1_O0(Tile_X0Y9_RES1_O0),
	.RES1_O1(Tile_X0Y9_RES1_O1),
	.RES1_O2(Tile_X0Y9_RES1_O2),
	.RES1_O3(Tile_X0Y9_RES1_O3),
	.RES2_O0(Tile_X0Y9_RES2_O0),
	.RES2_O1(Tile_X0Y9_RES2_O1),
	.RES2_O2(Tile_X0Y9_RES2_O2),
	.RES2_O3(Tile_X0Y9_RES2_O3),
	.FrameData(Tile_Y9_FrameData), 
	.FrameData_O(Tile_X0Y9_FrameData_O), 
	.FrameStrobe(Tile_X0Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X0Y9_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y9_LUT4AB (
	.N1END(Tile_X2Y10_N1BEG[3:0]),
	.N2MID(Tile_X2Y10_N2BEG[7:0]),
	.N2END(Tile_X2Y10_N2BEGb[7:0]),
	.N4END(Tile_X2Y10_N4BEG[15:0]),
	.NN4END(Tile_X2Y10_NN4BEG[15:0]),
	.Ci(Tile_X2Y10_Co[0:0]),
	.E1END(Tile_X1Y9_E1BEG[3:0]),
	.E2MID(Tile_X1Y9_E2BEG[7:0]),
	.E2END(Tile_X1Y9_E2BEGb[7:0]),
	.EE4END(Tile_X1Y9_EE4BEG[15:0]),
	.E6END(Tile_X1Y9_E6BEG[11:0]),
	.S1END(Tile_X2Y8_S1BEG[3:0]),
	.S2MID(Tile_X2Y8_S2BEG[7:0]),
	.S2END(Tile_X2Y8_S2BEGb[7:0]),
	.S4END(Tile_X2Y8_S4BEG[15:0]),
	.SS4END(Tile_X2Y8_SS4BEG[15:0]),
	.W1END(Tile_X3Y9_W1BEG[3:0]),
	.W2MID(Tile_X3Y9_W2BEG[7:0]),
	.W2END(Tile_X3Y9_W2BEGb[7:0]),
	.WW4END(Tile_X3Y9_WW4BEG[15:0]),
	.W6END(Tile_X3Y9_W6BEG[11:0]),
	.N1BEG(Tile_X2Y9_N1BEG[3:0]),
	.N2BEG(Tile_X2Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y9_NN4BEG[15:0]),
	.Co(Tile_X2Y9_Co[0:0]),
	.E1BEG(Tile_X2Y9_E1BEG[3:0]),
	.E2BEG(Tile_X2Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y9_E6BEG[11:0]),
	.S1BEG(Tile_X2Y9_S1BEG[3:0]),
	.S2BEG(Tile_X2Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y9_W1BEG[3:0]),
	.W2BEG(Tile_X2Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y9_FrameData_O), 
	.FrameData_O(Tile_X2Y9_FrameData_O), 
	.FrameStrobe(Tile_X2Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y9_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y9_LUT4AB (
	.N1END(Tile_X3Y10_N1BEG[3:0]),
	.N2MID(Tile_X3Y10_N2BEG[7:0]),
	.N2END(Tile_X3Y10_N2BEGb[7:0]),
	.N4END(Tile_X3Y10_N4BEG[15:0]),
	.NN4END(Tile_X3Y10_NN4BEG[15:0]),
	.Ci(Tile_X3Y10_Co[0:0]),
	.E1END(Tile_X2Y9_E1BEG[3:0]),
	.E2MID(Tile_X2Y9_E2BEG[7:0]),
	.E2END(Tile_X2Y9_E2BEGb[7:0]),
	.EE4END(Tile_X2Y9_EE4BEG[15:0]),
	.E6END(Tile_X2Y9_E6BEG[11:0]),
	.S1END(Tile_X3Y8_S1BEG[3:0]),
	.S2MID(Tile_X3Y8_S2BEG[7:0]),
	.S2END(Tile_X3Y8_S2BEGb[7:0]),
	.S4END(Tile_X3Y8_S4BEG[15:0]),
	.SS4END(Tile_X3Y8_SS4BEG[15:0]),
	.W1END(Tile_X4Y9_W1BEG[3:0]),
	.W2MID(Tile_X4Y9_W2BEG[7:0]),
	.W2END(Tile_X4Y9_W2BEGb[7:0]),
	.WW4END(Tile_X4Y9_WW4BEG[15:0]),
	.W6END(Tile_X4Y9_W6BEG[11:0]),
	.N1BEG(Tile_X3Y9_N1BEG[3:0]),
	.N2BEG(Tile_X3Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y9_NN4BEG[15:0]),
	.Co(Tile_X3Y9_Co[0:0]),
	.E1BEG(Tile_X3Y9_E1BEG[3:0]),
	.E2BEG(Tile_X3Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y9_E6BEG[11:0]),
	.S1BEG(Tile_X3Y9_S1BEG[3:0]),
	.S2BEG(Tile_X3Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y9_W1BEG[3:0]),
	.W2BEG(Tile_X3Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y9_FrameData_O), 
	.FrameData_O(Tile_X3Y9_FrameData_O), 
	.FrameStrobe(Tile_X3Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y9_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y9_LUT4AB (
	.N1END(Tile_X4Y10_N1BEG[3:0]),
	.N2MID(Tile_X4Y10_N2BEG[7:0]),
	.N2END(Tile_X4Y10_N2BEGb[7:0]),
	.N4END(Tile_X4Y10_N4BEG[15:0]),
	.NN4END(Tile_X4Y10_NN4BEG[15:0]),
	.Ci(Tile_X4Y10_Co[0:0]),
	.E1END(Tile_X3Y9_E1BEG[3:0]),
	.E2MID(Tile_X3Y9_E2BEG[7:0]),
	.E2END(Tile_X3Y9_E2BEGb[7:0]),
	.EE4END(Tile_X3Y9_EE4BEG[15:0]),
	.E6END(Tile_X3Y9_E6BEG[11:0]),
	.S1END(Tile_X4Y8_S1BEG[3:0]),
	.S2MID(Tile_X4Y8_S2BEG[7:0]),
	.S2END(Tile_X4Y8_S2BEGb[7:0]),
	.S4END(Tile_X4Y8_S4BEG[15:0]),
	.SS4END(Tile_X4Y8_SS4BEG[15:0]),
	.W1END(Tile_X5Y9_W1BEG[3:0]),
	.W2MID(Tile_X5Y9_W2BEG[7:0]),
	.W2END(Tile_X5Y9_W2BEGb[7:0]),
	.WW4END(Tile_X5Y9_WW4BEG[15:0]),
	.W6END(Tile_X5Y9_W6BEG[11:0]),
	.N1BEG(Tile_X4Y9_N1BEG[3:0]),
	.N2BEG(Tile_X4Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y9_NN4BEG[15:0]),
	.Co(Tile_X4Y9_Co[0:0]),
	.E1BEG(Tile_X4Y9_E1BEG[3:0]),
	.E2BEG(Tile_X4Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y9_E6BEG[11:0]),
	.S1BEG(Tile_X4Y9_S1BEG[3:0]),
	.S2BEG(Tile_X4Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y9_W1BEG[3:0]),
	.W2BEG(Tile_X4Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y9_FrameData_O), 
	.FrameData_O(Tile_X4Y9_FrameData_O), 
	.FrameStrobe(Tile_X4Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y9_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y9_LUT4AB (
	.N1END(Tile_X6Y10_N1BEG[3:0]),
	.N2MID(Tile_X6Y10_N2BEG[7:0]),
	.N2END(Tile_X6Y10_N2BEGb[7:0]),
	.N4END(Tile_X6Y10_N4BEG[15:0]),
	.NN4END(Tile_X6Y10_NN4BEG[15:0]),
	.Ci(Tile_X6Y10_Co[0:0]),
	.E1END(Tile_X5Y9_E1BEG[3:0]),
	.E2MID(Tile_X5Y9_E2BEG[7:0]),
	.E2END(Tile_X5Y9_E2BEGb[7:0]),
	.EE4END(Tile_X5Y9_EE4BEG[15:0]),
	.E6END(Tile_X5Y9_E6BEG[11:0]),
	.S1END(Tile_X6Y8_S1BEG[3:0]),
	.S2MID(Tile_X6Y8_S2BEG[7:0]),
	.S2END(Tile_X6Y8_S2BEGb[7:0]),
	.S4END(Tile_X6Y8_S4BEG[15:0]),
	.SS4END(Tile_X6Y8_SS4BEG[15:0]),
	.W1END(Tile_X7Y9_W1BEG[3:0]),
	.W2MID(Tile_X7Y9_W2BEG[7:0]),
	.W2END(Tile_X7Y9_W2BEGb[7:0]),
	.WW4END(Tile_X7Y9_WW4BEG[15:0]),
	.W6END(Tile_X7Y9_W6BEG[11:0]),
	.N1BEG(Tile_X6Y9_N1BEG[3:0]),
	.N2BEG(Tile_X6Y9_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y9_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y9_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y9_NN4BEG[15:0]),
	.Co(Tile_X6Y9_Co[0:0]),
	.E1BEG(Tile_X6Y9_E1BEG[3:0]),
	.E2BEG(Tile_X6Y9_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y9_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y9_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y9_E6BEG[11:0]),
	.S1BEG(Tile_X6Y9_S1BEG[3:0]),
	.S2BEG(Tile_X6Y9_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y9_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y9_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y9_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y9_W1BEG[3:0]),
	.W2BEG(Tile_X6Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y9_FrameData_O), 
	.FrameData_O(Tile_X6Y9_FrameData_O), 
	.FrameStrobe(Tile_X6Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y9_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y9_E_CPU_IO (
	.E1END(Tile_X6Y9_E1BEG[3:0]),
	.E2MID(Tile_X6Y9_E2BEG[7:0]),
	.E2END(Tile_X6Y9_E2BEGb[7:0]),
	.EE4END(Tile_X6Y9_EE4BEG[15:0]),
	.E6END(Tile_X6Y9_E6BEG[11:0]),
	.W1BEG(Tile_X7Y9_W1BEG[3:0]),
	.W2BEG(Tile_X7Y9_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y9_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y9_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y9_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y9_OPA_I0),
	.OPA_I1(Tile_X7Y9_OPA_I1),
	.OPA_I2(Tile_X7Y9_OPA_I2),
	.OPA_I3(Tile_X7Y9_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y9_OPB_I0),
	.OPB_I1(Tile_X7Y9_OPB_I1),
	.OPB_I2(Tile_X7Y9_OPB_I2),
	.OPB_I3(Tile_X7Y9_OPB_I3),
	.RES0_O0(Tile_X7Y9_RES0_O0),
	.RES0_O1(Tile_X7Y9_RES0_O1),
	.RES0_O2(Tile_X7Y9_RES0_O2),
	.RES0_O3(Tile_X7Y9_RES0_O3),
	.RES1_O0(Tile_X7Y9_RES1_O0),
	.RES1_O1(Tile_X7Y9_RES1_O1),
	.RES1_O2(Tile_X7Y9_RES1_O2),
	.RES1_O3(Tile_X7Y9_RES1_O3),
	.RES2_O0(Tile_X7Y9_RES2_O0),
	.RES2_O1(Tile_X7Y9_RES2_O1),
	.RES2_O2(Tile_X7Y9_RES2_O2),
	.RES2_O3(Tile_X7Y9_RES2_O3),
	.FrameData(Tile_X6Y9_FrameData_O), 
	.FrameData_O(Tile_X7Y9_FrameData_O), 
	.FrameStrobe(Tile_X7Y10_FrameStrobe_O),
	.FrameStrobe_O(Tile_X7Y9_FrameStrobe_O)
	);

	W_CPU_IO Tile_X0Y10_W_CPU_IO (
	.W1END(Tile_X1Y10_W1BEG[3:0]),
	.W2MID(Tile_X1Y10_W2BEG[7:0]),
	.W2END(Tile_X1Y10_W2BEGb[7:0]),
	.WW4END(Tile_X1Y10_WW4BEG[15:0]),
	.W6END(Tile_X1Y10_W6BEG[11:0]),
	.E1BEG(Tile_X0Y10_E1BEG[3:0]),
	.E2BEG(Tile_X0Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X0Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X0Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X0Y10_E6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X0Y10_OPA_I0),
	.OPA_I1(Tile_X0Y10_OPA_I1),
	.OPA_I2(Tile_X0Y10_OPA_I2),
	.OPA_I3(Tile_X0Y10_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X0Y10_OPB_I0),
	.OPB_I1(Tile_X0Y10_OPB_I1),
	.OPB_I2(Tile_X0Y10_OPB_I2),
	.OPB_I3(Tile_X0Y10_OPB_I3),
	.RES0_O0(Tile_X0Y10_RES0_O0),
	.RES0_O1(Tile_X0Y10_RES0_O1),
	.RES0_O2(Tile_X0Y10_RES0_O2),
	.RES0_O3(Tile_X0Y10_RES0_O3),
	.RES1_O0(Tile_X0Y10_RES1_O0),
	.RES1_O1(Tile_X0Y10_RES1_O1),
	.RES1_O2(Tile_X0Y10_RES1_O2),
	.RES1_O3(Tile_X0Y10_RES1_O3),
	.RES2_O0(Tile_X0Y10_RES2_O0),
	.RES2_O1(Tile_X0Y10_RES2_O1),
	.RES2_O2(Tile_X0Y10_RES2_O2),
	.RES2_O3(Tile_X0Y10_RES2_O3),
	.FrameData(Tile_Y10_FrameData), 
	.FrameData_O(Tile_X0Y10_FrameData_O), 
	.FrameStrobe(Tile_X0_FrameStrobe),
	.FrameStrobe_O(Tile_X0Y10_FrameStrobe_O)
	);


	LUT4AB Tile_X2Y10_LUT4AB (
	.N1END(Tile_X2Y11_N1BEG[3:0]),
	.N2MID(Tile_X2Y11_N2BEG[7:0]),
	.N2END(Tile_X2Y11_N2BEGb[7:0]),
	.N4END(Tile_X2Y11_N4BEG[15:0]),
	.NN4END(Tile_X2Y11_NN4BEG[15:0]),
	.Ci(Tile_X2Y11_Co[0:0]),
	.E1END(Tile_X1Y10_E1BEG[3:0]),
	.E2MID(Tile_X1Y10_E2BEG[7:0]),
	.E2END(Tile_X1Y10_E2BEGb[7:0]),
	.EE4END(Tile_X1Y10_EE4BEG[15:0]),
	.E6END(Tile_X1Y10_E6BEG[11:0]),
	.S1END(Tile_X2Y9_S1BEG[3:0]),
	.S2MID(Tile_X2Y9_S2BEG[7:0]),
	.S2END(Tile_X2Y9_S2BEGb[7:0]),
	.S4END(Tile_X2Y9_S4BEG[15:0]),
	.SS4END(Tile_X2Y9_SS4BEG[15:0]),
	.W1END(Tile_X3Y10_W1BEG[3:0]),
	.W2MID(Tile_X3Y10_W2BEG[7:0]),
	.W2END(Tile_X3Y10_W2BEGb[7:0]),
	.WW4END(Tile_X3Y10_WW4BEG[15:0]),
	.W6END(Tile_X3Y10_W6BEG[11:0]),
	.N1BEG(Tile_X2Y10_N1BEG[3:0]),
	.N2BEG(Tile_X2Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y10_NN4BEG[15:0]),
	.Co(Tile_X2Y10_Co[0:0]),
	.E1BEG(Tile_X2Y10_E1BEG[3:0]),
	.E2BEG(Tile_X2Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X2Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X2Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X2Y10_E6BEG[11:0]),
	.S1BEG(Tile_X2Y10_S1BEG[3:0]),
	.S2BEG(Tile_X2Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X2Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X2Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X2Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X2Y10_W1BEG[3:0]),
	.W2BEG(Tile_X2Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X2Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X2Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X2Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X1Y10_FrameData_O), 
	.FrameData_O(Tile_X2Y10_FrameData_O), 
	.FrameStrobe(Tile_X2Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X2Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X3Y10_LUT4AB (
	.N1END(Tile_X3Y11_N1BEG[3:0]),
	.N2MID(Tile_X3Y11_N2BEG[7:0]),
	.N2END(Tile_X3Y11_N2BEGb[7:0]),
	.N4END(Tile_X3Y11_N4BEG[15:0]),
	.NN4END(Tile_X3Y11_NN4BEG[15:0]),
	.Ci(Tile_X3Y11_Co[0:0]),
	.E1END(Tile_X2Y10_E1BEG[3:0]),
	.E2MID(Tile_X2Y10_E2BEG[7:0]),
	.E2END(Tile_X2Y10_E2BEGb[7:0]),
	.EE4END(Tile_X2Y10_EE4BEG[15:0]),
	.E6END(Tile_X2Y10_E6BEG[11:0]),
	.S1END(Tile_X3Y9_S1BEG[3:0]),
	.S2MID(Tile_X3Y9_S2BEG[7:0]),
	.S2END(Tile_X3Y9_S2BEGb[7:0]),
	.S4END(Tile_X3Y9_S4BEG[15:0]),
	.SS4END(Tile_X3Y9_SS4BEG[15:0]),
	.W1END(Tile_X4Y10_W1BEG[3:0]),
	.W2MID(Tile_X4Y10_W2BEG[7:0]),
	.W2END(Tile_X4Y10_W2BEGb[7:0]),
	.WW4END(Tile_X4Y10_WW4BEG[15:0]),
	.W6END(Tile_X4Y10_W6BEG[11:0]),
	.N1BEG(Tile_X3Y10_N1BEG[3:0]),
	.N2BEG(Tile_X3Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y10_NN4BEG[15:0]),
	.Co(Tile_X3Y10_Co[0:0]),
	.E1BEG(Tile_X3Y10_E1BEG[3:0]),
	.E2BEG(Tile_X3Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X3Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X3Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X3Y10_E6BEG[11:0]),
	.S1BEG(Tile_X3Y10_S1BEG[3:0]),
	.S2BEG(Tile_X3Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X3Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X3Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X3Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X3Y10_W1BEG[3:0]),
	.W2BEG(Tile_X3Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X3Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X3Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X3Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X2Y10_FrameData_O), 
	.FrameData_O(Tile_X3Y10_FrameData_O), 
	.FrameStrobe(Tile_X3Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X3Y10_FrameStrobe_O)
	);

	LUT4AB Tile_X4Y10_LUT4AB (
	.N1END(Tile_X4Y11_N1BEG[3:0]),
	.N2MID(Tile_X4Y11_N2BEG[7:0]),
	.N2END(Tile_X4Y11_N2BEGb[7:0]),
	.N4END(Tile_X4Y11_N4BEG[15:0]),
	.NN4END(Tile_X4Y11_NN4BEG[15:0]),
	.Ci(Tile_X4Y11_Co[0:0]),
	.E1END(Tile_X3Y10_E1BEG[3:0]),
	.E2MID(Tile_X3Y10_E2BEG[7:0]),
	.E2END(Tile_X3Y10_E2BEGb[7:0]),
	.EE4END(Tile_X3Y10_EE4BEG[15:0]),
	.E6END(Tile_X3Y10_E6BEG[11:0]),
	.S1END(Tile_X4Y9_S1BEG[3:0]),
	.S2MID(Tile_X4Y9_S2BEG[7:0]),
	.S2END(Tile_X4Y9_S2BEGb[7:0]),
	.S4END(Tile_X4Y9_S4BEG[15:0]),
	.SS4END(Tile_X4Y9_SS4BEG[15:0]),
	.W1END(Tile_X5Y10_W1BEG[3:0]),
	.W2MID(Tile_X5Y10_W2BEG[7:0]),
	.W2END(Tile_X5Y10_W2BEGb[7:0]),
	.WW4END(Tile_X5Y10_WW4BEG[15:0]),
	.W6END(Tile_X5Y10_W6BEG[11:0]),
	.N1BEG(Tile_X4Y10_N1BEG[3:0]),
	.N2BEG(Tile_X4Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y10_NN4BEG[15:0]),
	.Co(Tile_X4Y10_Co[0:0]),
	.E1BEG(Tile_X4Y10_E1BEG[3:0]),
	.E2BEG(Tile_X4Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X4Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X4Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X4Y10_E6BEG[11:0]),
	.S1BEG(Tile_X4Y10_S1BEG[3:0]),
	.S2BEG(Tile_X4Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X4Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X4Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X4Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X4Y10_W1BEG[3:0]),
	.W2BEG(Tile_X4Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X4Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X4Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X4Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X3Y10_FrameData_O), 
	.FrameData_O(Tile_X4Y10_FrameData_O), 
	.FrameStrobe(Tile_X4Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X4Y10_FrameStrobe_O)
	);


	LUT4AB Tile_X6Y10_LUT4AB (
	.N1END(Tile_X6Y11_N1BEG[3:0]),
	.N2MID(Tile_X6Y11_N2BEG[7:0]),
	.N2END(Tile_X6Y11_N2BEGb[7:0]),
	.N4END(Tile_X6Y11_N4BEG[15:0]),
	.NN4END(Tile_X6Y11_NN4BEG[15:0]),
	.Ci(Tile_X6Y11_Co[0:0]),
	.E1END(Tile_X5Y10_E1BEG[3:0]),
	.E2MID(Tile_X5Y10_E2BEG[7:0]),
	.E2END(Tile_X5Y10_E2BEGb[7:0]),
	.EE4END(Tile_X5Y10_EE4BEG[15:0]),
	.E6END(Tile_X5Y10_E6BEG[11:0]),
	.S1END(Tile_X6Y9_S1BEG[3:0]),
	.S2MID(Tile_X6Y9_S2BEG[7:0]),
	.S2END(Tile_X6Y9_S2BEGb[7:0]),
	.S4END(Tile_X6Y9_S4BEG[15:0]),
	.SS4END(Tile_X6Y9_SS4BEG[15:0]),
	.W1END(Tile_X7Y10_W1BEG[3:0]),
	.W2MID(Tile_X7Y10_W2BEG[7:0]),
	.W2END(Tile_X7Y10_W2BEGb[7:0]),
	.WW4END(Tile_X7Y10_WW4BEG[15:0]),
	.W6END(Tile_X7Y10_W6BEG[11:0]),
	.N1BEG(Tile_X6Y10_N1BEG[3:0]),
	.N2BEG(Tile_X6Y10_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y10_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y10_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y10_NN4BEG[15:0]),
	.Co(Tile_X6Y10_Co[0:0]),
	.E1BEG(Tile_X6Y10_E1BEG[3:0]),
	.E2BEG(Tile_X6Y10_E2BEG[7:0]),
	.E2BEGb(Tile_X6Y10_E2BEGb[7:0]),
	.EE4BEG(Tile_X6Y10_EE4BEG[15:0]),
	.E6BEG(Tile_X6Y10_E6BEG[11:0]),
	.S1BEG(Tile_X6Y10_S1BEG[3:0]),
	.S2BEG(Tile_X6Y10_S2BEG[7:0]),
	.S2BEGb(Tile_X6Y10_S2BEGb[7:0]),
	.S4BEG(Tile_X6Y10_S4BEG[15:0]),
	.SS4BEG(Tile_X6Y10_SS4BEG[15:0]),
	.W1BEG(Tile_X6Y10_W1BEG[3:0]),
	.W2BEG(Tile_X6Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X6Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X6Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X6Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.UserCLK(UserCLK),
	.FrameData(Tile_X5Y10_FrameData_O), 
	.FrameData_O(Tile_X6Y10_FrameData_O), 
	.FrameStrobe(Tile_X6Y11_FrameStrobe_O),
	.FrameStrobe_O(Tile_X6Y10_FrameStrobe_O)
	);

	E_CPU_IO Tile_X7Y10_E_CPU_IO (
	.E1END(Tile_X6Y10_E1BEG[3:0]),
	.E2MID(Tile_X6Y10_E2BEG[7:0]),
	.E2END(Tile_X6Y10_E2BEGb[7:0]),
	.EE4END(Tile_X6Y10_EE4BEG[15:0]),
	.E6END(Tile_X6Y10_E6BEG[11:0]),
	.W1BEG(Tile_X7Y10_W1BEG[3:0]),
	.W2BEG(Tile_X7Y10_W2BEG[7:0]),
	.W2BEGb(Tile_X7Y10_W2BEGb[7:0]),
	.WW4BEG(Tile_X7Y10_WW4BEG[15:0]),
	.W6BEG(Tile_X7Y10_W6BEG[11:0]),
	//tile IO port which gets directly connected to top-level tile module
	.OPA_I0(Tile_X7Y10_OPA_I0),
	.OPA_I1(Tile_X7Y10_OPA_I1),
	.OPA_I2(Tile_X7Y10_OPA_I2),
	.OPA_I3(Tile_X7Y10_OPA_I3),
	.UserCLK(UserCLK),
	.OPB_I0(Tile_X7Y10_OPB_I0),
	.OPB_I1(Tile_X7Y10_OPB_I1),
	.OPB_I2(Tile_X7Y10_OPB_I2),
	.OPB_I3(Tile_X7Y10_OPB_I3),
	.RES0_O0(Tile_X7Y10_RES0_O0),
	.RES0_O1(Tile_X7Y10_RES0_O1),
	.RES0_O2(Tile_X7Y10_RES0_O2),
	.RES0_O3(Tile_X7Y10_RES0_O3),
	.RES1_O0(Tile_X7Y10_RES1_O0),
	.RES1_O1(Tile_X7Y10_RES1_O1),
	.RES1_O2(Tile_X7Y10_RES1_O2),
	.RES1_O3(Tile_X7Y10_RES1_O3),
	.RES2_O0(Tile_X7Y10_RES2_O0),
	.RES2_O1(Tile_X7Y10_RES2_O1),
	.RES2_O2(Tile_X7Y10_RES2_O2),
	.RES2_O3(Tile_X7Y10_RES2_O3),
	.FrameData(Tile_X6Y10_FrameData_O), 
	.FrameData_O(Tile_X7Y10_FrameData_O), 
	.FrameStrobe(Tile_X7_FrameStrobe),
	.FrameStrobe_O(Tile_X7Y10_FrameStrobe_O)
	);

	S_term_DSP Tile_X1Y11_S_term_DSP (
	.S1END(Tile_X1Y10_S1BEG[3:0]),
	.S2MID(Tile_X1Y10_S2BEG[7:0]),
	.S2END(Tile_X1Y10_S2BEGb[7:0]),
	.S4END(Tile_X1Y10_S4BEG[15:0]),
	.SS4END(Tile_X1Y10_SS4BEG[15:0]),
	.N1BEG(Tile_X1Y11_N1BEG[3:0]),
	.N2BEG(Tile_X1Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X1Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X1Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X1Y11_NN4BEG[15:0]),
	.FrameData(Tile_Y11_FrameData), 
	.FrameData_O(Tile_X1Y11_FrameData_O), 
	.FrameStrobe(Tile_X1_FrameStrobe),
	.FrameStrobe_O(Tile_X1Y11_FrameStrobe_O)
	);

	S_term_single Tile_X2Y11_S_term_single (
	.S1END(Tile_X2Y10_S1BEG[3:0]),
	.S2MID(Tile_X2Y10_S2BEG[7:0]),
	.S2END(Tile_X2Y10_S2BEGb[7:0]),
	.S4END(Tile_X2Y10_S4BEG[15:0]),
	.SS4END(Tile_X2Y10_SS4BEG[15:0]),
	.N1BEG(Tile_X2Y11_N1BEG[3:0]),
	.N2BEG(Tile_X2Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X2Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X2Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X2Y11_NN4BEG[15:0]),
	.Co(Tile_X2Y11_Co[0:0]),
	.FrameData(Tile_X1Y11_FrameData_O), 
	.FrameData_O(Tile_X2Y11_FrameData_O), 
	.FrameStrobe(Tile_X2_FrameStrobe),
	.FrameStrobe_O(Tile_X2Y11_FrameStrobe_O)
	);

	S_term_single Tile_X3Y11_S_term_single (
	.S1END(Tile_X3Y10_S1BEG[3:0]),
	.S2MID(Tile_X3Y10_S2BEG[7:0]),
	.S2END(Tile_X3Y10_S2BEGb[7:0]),
	.S4END(Tile_X3Y10_S4BEG[15:0]),
	.SS4END(Tile_X3Y10_SS4BEG[15:0]),
	.N1BEG(Tile_X3Y11_N1BEG[3:0]),
	.N2BEG(Tile_X3Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X3Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X3Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X3Y11_NN4BEG[15:0]),
	.Co(Tile_X3Y11_Co[0:0]),
	.FrameData(Tile_X2Y11_FrameData_O), 
	.FrameData_O(Tile_X3Y11_FrameData_O), 
	.FrameStrobe(Tile_X3_FrameStrobe),
	.FrameStrobe_O(Tile_X3Y11_FrameStrobe_O)
	);

	S_term_single Tile_X4Y11_S_term_single (
	.S1END(Tile_X4Y10_S1BEG[3:0]),
	.S2MID(Tile_X4Y10_S2BEG[7:0]),
	.S2END(Tile_X4Y10_S2BEGb[7:0]),
	.S4END(Tile_X4Y10_S4BEG[15:0]),
	.SS4END(Tile_X4Y10_SS4BEG[15:0]),
	.N1BEG(Tile_X4Y11_N1BEG[3:0]),
	.N2BEG(Tile_X4Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X4Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X4Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X4Y11_NN4BEG[15:0]),
	.Co(Tile_X4Y11_Co[0:0]),
	.FrameData(Tile_X3Y11_FrameData_O), 
	.FrameData_O(Tile_X4Y11_FrameData_O), 
	.FrameStrobe(Tile_X4_FrameStrobe),
	.FrameStrobe_O(Tile_X4Y11_FrameStrobe_O)
	);

	S_term_DSP Tile_X5Y11_S_term_DSP (
	.S1END(Tile_X5Y10_S1BEG[3:0]),
	.S2MID(Tile_X5Y10_S2BEG[7:0]),
	.S2END(Tile_X5Y10_S2BEGb[7:0]),
	.S4END(Tile_X5Y10_S4BEG[15:0]),
	.SS4END(Tile_X5Y10_SS4BEG[15:0]),
	.N1BEG(Tile_X5Y11_N1BEG[3:0]),
	.N2BEG(Tile_X5Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X5Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X5Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X5Y11_NN4BEG[15:0]),
	.FrameData(Tile_X4Y11_FrameData_O), 
	.FrameData_O(Tile_X5Y11_FrameData_O), 
	.FrameStrobe(Tile_X5_FrameStrobe),
	.FrameStrobe_O(Tile_X5Y11_FrameStrobe_O)
	);

	S_term_single Tile_X6Y11_S_term_single (
	.S1END(Tile_X6Y10_S1BEG[3:0]),
	.S2MID(Tile_X6Y10_S2BEG[7:0]),
	.S2END(Tile_X6Y10_S2BEGb[7:0]),
	.S4END(Tile_X6Y10_S4BEG[15:0]),
	.SS4END(Tile_X6Y10_SS4BEG[15:0]),
	.N1BEG(Tile_X6Y11_N1BEG[3:0]),
	.N2BEG(Tile_X6Y11_N2BEG[7:0]),
	.N2BEGb(Tile_X6Y11_N2BEGb[7:0]),
	.N4BEG(Tile_X6Y11_N4BEG[15:0]),
	.NN4BEG(Tile_X6Y11_NN4BEG[15:0]),
	.Co(Tile_X6Y11_Co[0:0]),
	.FrameData(Tile_X5Y11_FrameData_O), 
	.FrameData_O(Tile_X6Y11_FrameData_O), 
	.FrameStrobe(Tile_X6_FrameStrobe),
	.FrameStrobe_O(Tile_X6Y11_FrameStrobe_O)
	);


	DSP Tile_X1Y1_X1Y2_DSP_tile (
	.top_E1END(Tile_X0Y1_E1BEG[3:0]),
	.top_E2MID(Tile_X0Y1_E2BEG[7:0]),
	.top_E2END(Tile_X0Y1_E2BEGb[7:0]),
	.top_EE4END(Tile_X0Y1_EE4BEG[15:0]),
	.top_E6END(Tile_X0Y1_E6BEG[11:0]),
	.top_S1END(Tile_X1Y0_S1BEG[3:0]),
	.top_S2MID(Tile_X1Y0_S2BEG[7:0]),
	.top_S2END(Tile_X1Y0_S2BEGb[7:0]),
	.top_S4END(Tile_X1Y0_S4BEG[15:0]),
	.top_SS4END(Tile_X1Y0_SS4BEG[15:0]),
	.top_W1END(Tile_X2Y1_W1BEG[3:0]),
	.top_W2MID(Tile_X2Y1_W2BEG[7:0]),
	.top_W2END(Tile_X2Y1_W2BEGb[7:0]),
	.top_WW4END(Tile_X2Y1_WW4BEG[15:0]),
	.top_W6END(Tile_X2Y1_W6BEG[11:0]),
	.top_N1BEG(Tile_X1Y1_N1BEG[3:0]),
	.top_N2BEG(Tile_X1Y1_N2BEG[7:0]),
	.top_N2BEGb(Tile_X1Y1_N2BEGb[7:0]),
	.top_N4BEG(Tile_X1Y1_N4BEG[15:0]),
	.top_NN4BEG(Tile_X1Y1_NN4BEG[15:0]),
	.top_E1BEG(Tile_X1Y1_E1BEG[3:0]),
	.top_E2BEG(Tile_X1Y1_E2BEG[7:0]),
	.top_E2BEGb(Tile_X1Y1_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X1Y1_EE4BEG[15:0]),
	.top_E6BEG(Tile_X1Y1_E6BEG[11:0]),
	.top_W1BEG(Tile_X1Y1_W1BEG[3:0]),
	.top_W2BEG(Tile_X1Y1_W2BEG[7:0]),
	.top_W2BEGb(Tile_X1Y1_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X1Y1_WW4BEG[15:0]),
	.top_W6BEG(Tile_X1Y1_W6BEG[11:0]),
	.top_FrameData(Tile_X0Y1_FrameData_O),
	.top_FrameData_O(Tile_X1Y1_FrameData_O),
	.FrameStrobe_O(Tile_X1Y1_FrameStrobe_O),
	.bot_N1END(Tile_X1Y3_N1BEG[3:0]),
	.bot_N2MID(Tile_X1Y3_N2BEG[7:0]),
	.bot_N2END(Tile_X1Y3_N2BEGb[7:0]),
	.bot_N4END(Tile_X1Y3_N4BEG[15:0]),
	.bot_NN4END(Tile_X1Y3_NN4BEG[15:0]),
	.bot_E1END(Tile_X0Y2_E1BEG[3:0]),
	.bot_E2MID(Tile_X0Y2_E2BEG[7:0]),
	.bot_E2END(Tile_X0Y2_E2BEGb[7:0]),
	.bot_EE4END(Tile_X0Y2_EE4BEG[15:0]),
	.bot_E6END(Tile_X0Y2_E6BEG[11:0]),
	.bot_W1END(Tile_X2Y2_W1BEG[3:0]),
	.bot_W2MID(Tile_X2Y2_W2BEG[7:0]),
	.bot_W2END(Tile_X2Y2_W2BEGb[7:0]),
	.bot_WW4END(Tile_X2Y2_WW4BEG[15:0]),
	.bot_W6END(Tile_X2Y2_W6BEG[11:0]),
	.bot_E1BEG(Tile_X1Y2_E1BEG[3:0]),
	.bot_E2BEG(Tile_X1Y2_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X1Y2_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X1Y2_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X1Y2_E6BEG[11:0]),
	.bot_S1BEG(Tile_X1Y2_S1BEG[3:0]),
	.bot_S2BEG(Tile_X1Y2_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X1Y2_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X1Y2_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X1Y2_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X1Y2_W1BEG[3:0]),
	.bot_W2BEG(Tile_X1Y2_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X1Y2_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X1Y2_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X1Y2_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X0Y2_FrameData_O),
	.bot_FrameData_O(Tile_X1Y2_FrameData_O),
	.FrameStrobe(Tile_X1Y3_FrameStrobe_O)
	);

	DSP Tile_X5Y1_X5Y2_DSP_tile (
	.top_E1END(Tile_X4Y1_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y1_E2BEG[7:0]),
	.top_E2END(Tile_X4Y1_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y1_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y1_E6BEG[11:0]),
	.top_S1END(Tile_X5Y0_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y0_S2BEG[7:0]),
	.top_S2END(Tile_X5Y0_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y0_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y0_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y1_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y1_W2BEG[7:0]),
	.top_W2END(Tile_X6Y1_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y1_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y1_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y1_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y1_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y1_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y1_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y1_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y1_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y1_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y1_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y1_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y1_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y1_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y1_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y1_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y1_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y1_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y1_FrameData_O),
	.top_FrameData_O(Tile_X5Y1_FrameData_O),
	.FrameStrobe_O(Tile_X5Y1_FrameStrobe_O),
	.bot_N1END(Tile_X5Y3_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y3_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y3_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y3_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y3_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y2_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y2_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y2_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y2_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y2_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y2_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y2_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y2_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y2_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y2_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y2_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y2_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y2_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y2_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y2_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y2_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y2_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y2_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y2_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y2_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y2_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y2_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y2_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y2_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y2_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X4Y2_FrameData_O),
	.bot_FrameData_O(Tile_X5Y2_FrameData_O),
	.FrameStrobe(Tile_X5Y3_FrameStrobe_O)
	);

	DSP Tile_X1Y3_X1Y4_DSP_tile (
	.top_E1END(Tile_X0Y3_E1BEG[3:0]),
	.top_E2MID(Tile_X0Y3_E2BEG[7:0]),
	.top_E2END(Tile_X0Y3_E2BEGb[7:0]),
	.top_EE4END(Tile_X0Y3_EE4BEG[15:0]),
	.top_E6END(Tile_X0Y3_E6BEG[11:0]),
	.top_S1END(Tile_X1Y2_S1BEG[3:0]),
	.top_S2MID(Tile_X1Y2_S2BEG[7:0]),
	.top_S2END(Tile_X1Y2_S2BEGb[7:0]),
	.top_S4END(Tile_X1Y2_S4BEG[15:0]),
	.top_SS4END(Tile_X1Y2_SS4BEG[15:0]),
	.top_W1END(Tile_X2Y3_W1BEG[3:0]),
	.top_W2MID(Tile_X2Y3_W2BEG[7:0]),
	.top_W2END(Tile_X2Y3_W2BEGb[7:0]),
	.top_WW4END(Tile_X2Y3_WW4BEG[15:0]),
	.top_W6END(Tile_X2Y3_W6BEG[11:0]),
	.top_N1BEG(Tile_X1Y3_N1BEG[3:0]),
	.top_N2BEG(Tile_X1Y3_N2BEG[7:0]),
	.top_N2BEGb(Tile_X1Y3_N2BEGb[7:0]),
	.top_N4BEG(Tile_X1Y3_N4BEG[15:0]),
	.top_NN4BEG(Tile_X1Y3_NN4BEG[15:0]),
	.top_E1BEG(Tile_X1Y3_E1BEG[3:0]),
	.top_E2BEG(Tile_X1Y3_E2BEG[7:0]),
	.top_E2BEGb(Tile_X1Y3_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X1Y3_EE4BEG[15:0]),
	.top_E6BEG(Tile_X1Y3_E6BEG[11:0]),
	.top_W1BEG(Tile_X1Y3_W1BEG[3:0]),
	.top_W2BEG(Tile_X1Y3_W2BEG[7:0]),
	.top_W2BEGb(Tile_X1Y3_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X1Y3_WW4BEG[15:0]),
	.top_W6BEG(Tile_X1Y3_W6BEG[11:0]),
	.top_FrameData(Tile_X0Y3_FrameData_O),
	.top_FrameData_O(Tile_X1Y3_FrameData_O),
	.FrameStrobe_O(Tile_X1Y3_FrameStrobe_O),
	.bot_N1END(Tile_X1Y5_N1BEG[3:0]),
	.bot_N2MID(Tile_X1Y5_N2BEG[7:0]),
	.bot_N2END(Tile_X1Y5_N2BEGb[7:0]),
	.bot_N4END(Tile_X1Y5_N4BEG[15:0]),
	.bot_NN4END(Tile_X1Y5_NN4BEG[15:0]),
	.bot_E1END(Tile_X0Y4_E1BEG[3:0]),
	.bot_E2MID(Tile_X0Y4_E2BEG[7:0]),
	.bot_E2END(Tile_X0Y4_E2BEGb[7:0]),
	.bot_EE4END(Tile_X0Y4_EE4BEG[15:0]),
	.bot_E6END(Tile_X0Y4_E6BEG[11:0]),
	.bot_W1END(Tile_X2Y4_W1BEG[3:0]),
	.bot_W2MID(Tile_X2Y4_W2BEG[7:0]),
	.bot_W2END(Tile_X2Y4_W2BEGb[7:0]),
	.bot_WW4END(Tile_X2Y4_WW4BEG[15:0]),
	.bot_W6END(Tile_X2Y4_W6BEG[11:0]),
	.bot_E1BEG(Tile_X1Y4_E1BEG[3:0]),
	.bot_E2BEG(Tile_X1Y4_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X1Y4_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X1Y4_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X1Y4_E6BEG[11:0]),
	.bot_S1BEG(Tile_X1Y4_S1BEG[3:0]),
	.bot_S2BEG(Tile_X1Y4_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X1Y4_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X1Y4_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X1Y4_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X1Y4_W1BEG[3:0]),
	.bot_W2BEG(Tile_X1Y4_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X1Y4_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X1Y4_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X1Y4_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X0Y4_FrameData_O),
	.bot_FrameData_O(Tile_X1Y4_FrameData_O),
	.FrameStrobe(Tile_X1Y5_FrameStrobe_O)
	);

	DSP Tile_X5Y3_X5Y4_DSP_tile (
	.top_E1END(Tile_X4Y3_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y3_E2BEG[7:0]),
	.top_E2END(Tile_X4Y3_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y3_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y3_E6BEG[11:0]),
	.top_S1END(Tile_X5Y2_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y2_S2BEG[7:0]),
	.top_S2END(Tile_X5Y2_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y2_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y2_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y3_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y3_W2BEG[7:0]),
	.top_W2END(Tile_X6Y3_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y3_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y3_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y3_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y3_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y3_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y3_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y3_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y3_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y3_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y3_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y3_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y3_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y3_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y3_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y3_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y3_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y3_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y3_FrameData_O),
	.top_FrameData_O(Tile_X5Y3_FrameData_O),
	.FrameStrobe_O(Tile_X5Y3_FrameStrobe_O),
	.bot_N1END(Tile_X5Y5_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y5_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y5_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y5_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y5_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y4_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y4_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y4_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y4_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y4_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y4_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y4_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y4_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y4_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y4_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y4_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y4_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y4_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y4_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y4_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y4_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y4_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y4_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y4_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y4_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y4_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y4_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y4_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y4_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y4_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X4Y4_FrameData_O),
	.bot_FrameData_O(Tile_X5Y4_FrameData_O),
	.FrameStrobe(Tile_X5Y5_FrameStrobe_O)
	);

	DSP Tile_X1Y5_X1Y6_DSP_tile (
	.top_E1END(Tile_X0Y5_E1BEG[3:0]),
	.top_E2MID(Tile_X0Y5_E2BEG[7:0]),
	.top_E2END(Tile_X0Y5_E2BEGb[7:0]),
	.top_EE4END(Tile_X0Y5_EE4BEG[15:0]),
	.top_E6END(Tile_X0Y5_E6BEG[11:0]),
	.top_S1END(Tile_X1Y4_S1BEG[3:0]),
	.top_S2MID(Tile_X1Y4_S2BEG[7:0]),
	.top_S2END(Tile_X1Y4_S2BEGb[7:0]),
	.top_S4END(Tile_X1Y4_S4BEG[15:0]),
	.top_SS4END(Tile_X1Y4_SS4BEG[15:0]),
	.top_W1END(Tile_X2Y5_W1BEG[3:0]),
	.top_W2MID(Tile_X2Y5_W2BEG[7:0]),
	.top_W2END(Tile_X2Y5_W2BEGb[7:0]),
	.top_WW4END(Tile_X2Y5_WW4BEG[15:0]),
	.top_W6END(Tile_X2Y5_W6BEG[11:0]),
	.top_N1BEG(Tile_X1Y5_N1BEG[3:0]),
	.top_N2BEG(Tile_X1Y5_N2BEG[7:0]),
	.top_N2BEGb(Tile_X1Y5_N2BEGb[7:0]),
	.top_N4BEG(Tile_X1Y5_N4BEG[15:0]),
	.top_NN4BEG(Tile_X1Y5_NN4BEG[15:0]),
	.top_E1BEG(Tile_X1Y5_E1BEG[3:0]),
	.top_E2BEG(Tile_X1Y5_E2BEG[7:0]),
	.top_E2BEGb(Tile_X1Y5_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X1Y5_EE4BEG[15:0]),
	.top_E6BEG(Tile_X1Y5_E6BEG[11:0]),
	.top_W1BEG(Tile_X1Y5_W1BEG[3:0]),
	.top_W2BEG(Tile_X1Y5_W2BEG[7:0]),
	.top_W2BEGb(Tile_X1Y5_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X1Y5_WW4BEG[15:0]),
	.top_W6BEG(Tile_X1Y5_W6BEG[11:0]),
	.top_FrameData(Tile_X0Y5_FrameData_O),
	.top_FrameData_O(Tile_X1Y5_FrameData_O),
	.FrameStrobe_O(Tile_X1Y5_FrameStrobe_O),
	.bot_N1END(Tile_X1Y7_N1BEG[3:0]),
	.bot_N2MID(Tile_X1Y7_N2BEG[7:0]),
	.bot_N2END(Tile_X1Y7_N2BEGb[7:0]),
	.bot_N4END(Tile_X1Y7_N4BEG[15:0]),
	.bot_NN4END(Tile_X1Y7_NN4BEG[15:0]),
	.bot_E1END(Tile_X0Y6_E1BEG[3:0]),
	.bot_E2MID(Tile_X0Y6_E2BEG[7:0]),
	.bot_E2END(Tile_X0Y6_E2BEGb[7:0]),
	.bot_EE4END(Tile_X0Y6_EE4BEG[15:0]),
	.bot_E6END(Tile_X0Y6_E6BEG[11:0]),
	.bot_W1END(Tile_X2Y6_W1BEG[3:0]),
	.bot_W2MID(Tile_X2Y6_W2BEG[7:0]),
	.bot_W2END(Tile_X2Y6_W2BEGb[7:0]),
	.bot_WW4END(Tile_X2Y6_WW4BEG[15:0]),
	.bot_W6END(Tile_X2Y6_W6BEG[11:0]),
	.bot_E1BEG(Tile_X1Y6_E1BEG[3:0]),
	.bot_E2BEG(Tile_X1Y6_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X1Y6_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X1Y6_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X1Y6_E6BEG[11:0]),
	.bot_S1BEG(Tile_X1Y6_S1BEG[3:0]),
	.bot_S2BEG(Tile_X1Y6_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X1Y6_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X1Y6_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X1Y6_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X1Y6_W1BEG[3:0]),
	.bot_W2BEG(Tile_X1Y6_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X1Y6_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X1Y6_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X1Y6_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X0Y6_FrameData_O),
	.bot_FrameData_O(Tile_X1Y6_FrameData_O),
	.FrameStrobe(Tile_X1Y7_FrameStrobe_O)
	);

	DSP Tile_X5Y5_X5Y6_DSP_tile (
	.top_E1END(Tile_X4Y5_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y5_E2BEG[7:0]),
	.top_E2END(Tile_X4Y5_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y5_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y5_E6BEG[11:0]),
	.top_S1END(Tile_X5Y4_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y4_S2BEG[7:0]),
	.top_S2END(Tile_X5Y4_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y4_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y4_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y5_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y5_W2BEG[7:0]),
	.top_W2END(Tile_X6Y5_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y5_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y5_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y5_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y5_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y5_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y5_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y5_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y5_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y5_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y5_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y5_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y5_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y5_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y5_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y5_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y5_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y5_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y5_FrameData_O),
	.top_FrameData_O(Tile_X5Y5_FrameData_O),
	.FrameStrobe_O(Tile_X5Y5_FrameStrobe_O),
	.bot_N1END(Tile_X5Y7_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y7_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y7_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y7_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y7_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y6_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y6_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y6_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y6_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y6_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y6_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y6_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y6_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y6_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y6_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y6_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y6_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y6_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y6_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y6_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y6_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y6_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y6_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y6_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y6_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y6_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y6_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y6_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y6_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y6_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X4Y6_FrameData_O),
	.bot_FrameData_O(Tile_X5Y6_FrameData_O),
	.FrameStrobe(Tile_X5Y7_FrameStrobe_O)
	);

	DSP Tile_X1Y7_X1Y8_DSP_tile (
	.top_E1END(Tile_X0Y7_E1BEG[3:0]),
	.top_E2MID(Tile_X0Y7_E2BEG[7:0]),
	.top_E2END(Tile_X0Y7_E2BEGb[7:0]),
	.top_EE4END(Tile_X0Y7_EE4BEG[15:0]),
	.top_E6END(Tile_X0Y7_E6BEG[11:0]),
	.top_S1END(Tile_X1Y6_S1BEG[3:0]),
	.top_S2MID(Tile_X1Y6_S2BEG[7:0]),
	.top_S2END(Tile_X1Y6_S2BEGb[7:0]),
	.top_S4END(Tile_X1Y6_S4BEG[15:0]),
	.top_SS4END(Tile_X1Y6_SS4BEG[15:0]),
	.top_W1END(Tile_X2Y7_W1BEG[3:0]),
	.top_W2MID(Tile_X2Y7_W2BEG[7:0]),
	.top_W2END(Tile_X2Y7_W2BEGb[7:0]),
	.top_WW4END(Tile_X2Y7_WW4BEG[15:0]),
	.top_W6END(Tile_X2Y7_W6BEG[11:0]),
	.top_N1BEG(Tile_X1Y7_N1BEG[3:0]),
	.top_N2BEG(Tile_X1Y7_N2BEG[7:0]),
	.top_N2BEGb(Tile_X1Y7_N2BEGb[7:0]),
	.top_N4BEG(Tile_X1Y7_N4BEG[15:0]),
	.top_NN4BEG(Tile_X1Y7_NN4BEG[15:0]),
	.top_E1BEG(Tile_X1Y7_E1BEG[3:0]),
	.top_E2BEG(Tile_X1Y7_E2BEG[7:0]),
	.top_E2BEGb(Tile_X1Y7_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X1Y7_EE4BEG[15:0]),
	.top_E6BEG(Tile_X1Y7_E6BEG[11:0]),
	.top_W1BEG(Tile_X1Y7_W1BEG[3:0]),
	.top_W2BEG(Tile_X1Y7_W2BEG[7:0]),
	.top_W2BEGb(Tile_X1Y7_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X1Y7_WW4BEG[15:0]),
	.top_W6BEG(Tile_X1Y7_W6BEG[11:0]),
	.top_FrameData(Tile_X0Y7_FrameData_O),
	.top_FrameData_O(Tile_X1Y7_FrameData_O),
	.FrameStrobe_O(Tile_X1Y7_FrameStrobe_O),
	.bot_N1END(Tile_X1Y9_N1BEG[3:0]),
	.bot_N2MID(Tile_X1Y9_N2BEG[7:0]),
	.bot_N2END(Tile_X1Y9_N2BEGb[7:0]),
	.bot_N4END(Tile_X1Y9_N4BEG[15:0]),
	.bot_NN4END(Tile_X1Y9_NN4BEG[15:0]),
	.bot_E1END(Tile_X0Y8_E1BEG[3:0]),
	.bot_E2MID(Tile_X0Y8_E2BEG[7:0]),
	.bot_E2END(Tile_X0Y8_E2BEGb[7:0]),
	.bot_EE4END(Tile_X0Y8_EE4BEG[15:0]),
	.bot_E6END(Tile_X0Y8_E6BEG[11:0]),
	.bot_W1END(Tile_X2Y8_W1BEG[3:0]),
	.bot_W2MID(Tile_X2Y8_W2BEG[7:0]),
	.bot_W2END(Tile_X2Y8_W2BEGb[7:0]),
	.bot_WW4END(Tile_X2Y8_WW4BEG[15:0]),
	.bot_W6END(Tile_X2Y8_W6BEG[11:0]),
	.bot_E1BEG(Tile_X1Y8_E1BEG[3:0]),
	.bot_E2BEG(Tile_X1Y8_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X1Y8_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X1Y8_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X1Y8_E6BEG[11:0]),
	.bot_S1BEG(Tile_X1Y8_S1BEG[3:0]),
	.bot_S2BEG(Tile_X1Y8_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X1Y8_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X1Y8_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X1Y8_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X1Y8_W1BEG[3:0]),
	.bot_W2BEG(Tile_X1Y8_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X1Y8_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X1Y8_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X1Y8_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X0Y8_FrameData_O),
	.bot_FrameData_O(Tile_X1Y8_FrameData_O),
	.FrameStrobe(Tile_X1Y9_FrameStrobe_O)
	);

	DSP Tile_X5Y7_X5Y8_DSP_tile (
	.top_E1END(Tile_X4Y7_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y7_E2BEG[7:0]),
	.top_E2END(Tile_X4Y7_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y7_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y7_E6BEG[11:0]),
	.top_S1END(Tile_X5Y6_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y6_S2BEG[7:0]),
	.top_S2END(Tile_X5Y6_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y6_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y6_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y7_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y7_W2BEG[7:0]),
	.top_W2END(Tile_X6Y7_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y7_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y7_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y7_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y7_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y7_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y7_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y7_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y7_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y7_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y7_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y7_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y7_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y7_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y7_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y7_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y7_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y7_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y7_FrameData_O),
	.top_FrameData_O(Tile_X5Y7_FrameData_O),
	.FrameStrobe_O(Tile_X5Y7_FrameStrobe_O),
	.bot_N1END(Tile_X5Y9_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y9_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y9_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y9_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y9_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y8_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y8_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y8_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y8_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y8_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y8_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y8_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y8_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y8_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y8_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y8_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y8_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y8_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y8_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y8_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y8_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y8_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y8_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y8_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y8_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y8_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y8_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y8_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y8_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y8_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X4Y8_FrameData_O),
	.bot_FrameData_O(Tile_X5Y8_FrameData_O),
	.FrameStrobe(Tile_X5Y9_FrameStrobe_O)
	);

	DSP Tile_X1Y9_X1Y10_DSP_tile (
	.top_E1END(Tile_X0Y9_E1BEG[3:0]),
	.top_E2MID(Tile_X0Y9_E2BEG[7:0]),
	.top_E2END(Tile_X0Y9_E2BEGb[7:0]),
	.top_EE4END(Tile_X0Y9_EE4BEG[15:0]),
	.top_E6END(Tile_X0Y9_E6BEG[11:0]),
	.top_S1END(Tile_X1Y8_S1BEG[3:0]),
	.top_S2MID(Tile_X1Y8_S2BEG[7:0]),
	.top_S2END(Tile_X1Y8_S2BEGb[7:0]),
	.top_S4END(Tile_X1Y8_S4BEG[15:0]),
	.top_SS4END(Tile_X1Y8_SS4BEG[15:0]),
	.top_W1END(Tile_X2Y9_W1BEG[3:0]),
	.top_W2MID(Tile_X2Y9_W2BEG[7:0]),
	.top_W2END(Tile_X2Y9_W2BEGb[7:0]),
	.top_WW4END(Tile_X2Y9_WW4BEG[15:0]),
	.top_W6END(Tile_X2Y9_W6BEG[11:0]),
	.top_N1BEG(Tile_X1Y9_N1BEG[3:0]),
	.top_N2BEG(Tile_X1Y9_N2BEG[7:0]),
	.top_N2BEGb(Tile_X1Y9_N2BEGb[7:0]),
	.top_N4BEG(Tile_X1Y9_N4BEG[15:0]),
	.top_NN4BEG(Tile_X1Y9_NN4BEG[15:0]),
	.top_E1BEG(Tile_X1Y9_E1BEG[3:0]),
	.top_E2BEG(Tile_X1Y9_E2BEG[7:0]),
	.top_E2BEGb(Tile_X1Y9_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X1Y9_EE4BEG[15:0]),
	.top_E6BEG(Tile_X1Y9_E6BEG[11:0]),
	.top_W1BEG(Tile_X1Y9_W1BEG[3:0]),
	.top_W2BEG(Tile_X1Y9_W2BEG[7:0]),
	.top_W2BEGb(Tile_X1Y9_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X1Y9_WW4BEG[15:0]),
	.top_W6BEG(Tile_X1Y9_W6BEG[11:0]),
	.top_FrameData(Tile_X0Y9_FrameData_O),
	.top_FrameData_O(Tile_X1Y9_FrameData_O),
	.FrameStrobe_O(Tile_X1Y9_FrameStrobe_O),
	.bot_N1END(Tile_X1Y11_N1BEG[3:0]),
	.bot_N2MID(Tile_X1Y11_N2BEG[7:0]),
	.bot_N2END(Tile_X1Y11_N2BEGb[7:0]),
	.bot_N4END(Tile_X1Y11_N4BEG[15:0]),
	.bot_NN4END(Tile_X1Y11_NN4BEG[15:0]),
	.bot_E1END(Tile_X0Y10_E1BEG[3:0]),
	.bot_E2MID(Tile_X0Y10_E2BEG[7:0]),
	.bot_E2END(Tile_X0Y10_E2BEGb[7:0]),
	.bot_EE4END(Tile_X0Y10_EE4BEG[15:0]),
	.bot_E6END(Tile_X0Y10_E6BEG[11:0]),
	.bot_W1END(Tile_X2Y10_W1BEG[3:0]),
	.bot_W2MID(Tile_X2Y10_W2BEG[7:0]),
	.bot_W2END(Tile_X2Y10_W2BEGb[7:0]),
	.bot_WW4END(Tile_X2Y10_WW4BEG[15:0]),
	.bot_W6END(Tile_X2Y10_W6BEG[11:0]),
	.bot_E1BEG(Tile_X1Y10_E1BEG[3:0]),
	.bot_E2BEG(Tile_X1Y10_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X1Y10_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X1Y10_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X1Y10_E6BEG[11:0]),
	.bot_S1BEG(Tile_X1Y10_S1BEG[3:0]),
	.bot_S2BEG(Tile_X1Y10_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X1Y10_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X1Y10_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X1Y10_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X1Y10_W1BEG[3:0]),
	.bot_W2BEG(Tile_X1Y10_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X1Y10_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X1Y10_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X1Y10_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X0Y10_FrameData_O),
	.bot_FrameData_O(Tile_X1Y10_FrameData_O),
	.FrameStrobe(Tile_X1Y11_FrameStrobe_O)
	);

	DSP Tile_X5Y9_X5Y10_DSP_tile (
	.top_E1END(Tile_X4Y9_E1BEG[3:0]),
	.top_E2MID(Tile_X4Y9_E2BEG[7:0]),
	.top_E2END(Tile_X4Y9_E2BEGb[7:0]),
	.top_EE4END(Tile_X4Y9_EE4BEG[15:0]),
	.top_E6END(Tile_X4Y9_E6BEG[11:0]),
	.top_S1END(Tile_X5Y8_S1BEG[3:0]),
	.top_S2MID(Tile_X5Y8_S2BEG[7:0]),
	.top_S2END(Tile_X5Y8_S2BEGb[7:0]),
	.top_S4END(Tile_X5Y8_S4BEG[15:0]),
	.top_SS4END(Tile_X5Y8_SS4BEG[15:0]),
	.top_W1END(Tile_X6Y9_W1BEG[3:0]),
	.top_W2MID(Tile_X6Y9_W2BEG[7:0]),
	.top_W2END(Tile_X6Y9_W2BEGb[7:0]),
	.top_WW4END(Tile_X6Y9_WW4BEG[15:0]),
	.top_W6END(Tile_X6Y9_W6BEG[11:0]),
	.top_N1BEG(Tile_X5Y9_N1BEG[3:0]),
	.top_N2BEG(Tile_X5Y9_N2BEG[7:0]),
	.top_N2BEGb(Tile_X5Y9_N2BEGb[7:0]),
	.top_N4BEG(Tile_X5Y9_N4BEG[15:0]),
	.top_NN4BEG(Tile_X5Y9_NN4BEG[15:0]),
	.top_E1BEG(Tile_X5Y9_E1BEG[3:0]),
	.top_E2BEG(Tile_X5Y9_E2BEG[7:0]),
	.top_E2BEGb(Tile_X5Y9_E2BEGb[7:0]),
	.top_EE4BEG(Tile_X5Y9_EE4BEG[15:0]),
	.top_E6BEG(Tile_X5Y9_E6BEG[11:0]),
	.top_W1BEG(Tile_X5Y9_W1BEG[3:0]),
	.top_W2BEG(Tile_X5Y9_W2BEG[7:0]),
	.top_W2BEGb(Tile_X5Y9_W2BEGb[7:0]),
	.top_WW4BEG(Tile_X5Y9_WW4BEG[15:0]),
	.top_W6BEG(Tile_X5Y9_W6BEG[11:0]),
	.top_FrameData(Tile_X4Y9_FrameData_O),
	.top_FrameData_O(Tile_X5Y9_FrameData_O),
	.FrameStrobe_O(Tile_X5Y9_FrameStrobe_O),
	.bot_N1END(Tile_X5Y11_N1BEG[3:0]),
	.bot_N2MID(Tile_X5Y11_N2BEG[7:0]),
	.bot_N2END(Tile_X5Y11_N2BEGb[7:0]),
	.bot_N4END(Tile_X5Y11_N4BEG[15:0]),
	.bot_NN4END(Tile_X5Y11_NN4BEG[15:0]),
	.bot_E1END(Tile_X4Y10_E1BEG[3:0]),
	.bot_E2MID(Tile_X4Y10_E2BEG[7:0]),
	.bot_E2END(Tile_X4Y10_E2BEGb[7:0]),
	.bot_EE4END(Tile_X4Y10_EE4BEG[15:0]),
	.bot_E6END(Tile_X4Y10_E6BEG[11:0]),
	.bot_W1END(Tile_X6Y10_W1BEG[3:0]),
	.bot_W2MID(Tile_X6Y10_W2BEG[7:0]),
	.bot_W2END(Tile_X6Y10_W2BEGb[7:0]),
	.bot_WW4END(Tile_X6Y10_WW4BEG[15:0]),
	.bot_W6END(Tile_X6Y10_W6BEG[11:0]),
	.bot_E1BEG(Tile_X5Y10_E1BEG[3:0]),
	.bot_E2BEG(Tile_X5Y10_E2BEG[7:0]),
	.bot_E2BEGb(Tile_X5Y10_E2BEGb[7:0]),
	.bot_EE4BEG(Tile_X5Y10_EE4BEG[15:0]),
	.bot_E6BEG(Tile_X5Y10_E6BEG[11:0]),
	.bot_S1BEG(Tile_X5Y10_S1BEG[3:0]),
	.bot_S2BEG(Tile_X5Y10_S2BEG[7:0]),
	.bot_S2BEGb(Tile_X5Y10_S2BEGb[7:0]),
	.bot_S4BEG(Tile_X5Y10_S4BEG[15:0]),
	.bot_SS4BEG(Tile_X5Y10_SS4BEG[15:0]),
	.bot_W1BEG(Tile_X5Y10_W1BEG[3:0]),
	.bot_W2BEG(Tile_X5Y10_W2BEG[7:0]),
	.bot_W2BEGb(Tile_X5Y10_W2BEGb[7:0]),
	.bot_WW4BEG(Tile_X5Y10_WW4BEG[15:0]),
	.bot_W6BEG(Tile_X5Y10_W6BEG[11:0]),
	.UserCLK(UserCLK),
	.bot_FrameData(Tile_X4Y10_FrameData_O),
	.bot_FrameData_O(Tile_X5Y10_FrameData_O),
	.FrameStrobe(Tile_X5Y11_FrameStrobe_O)
	);

endmodule
