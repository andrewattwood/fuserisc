magic
tech sky130A
magscale 1 2
timestamp 1623936842
<< obsli1 >>
rect 1104 2159 238740 239377
<< obsm1 >>
rect 474 1776 238740 239488
<< metal2 >>
rect 1398 241210 1454 242010
rect 4158 241210 4214 242010
rect 6918 241210 6974 242010
rect 10138 241210 10194 242010
rect 12898 241210 12954 242010
rect 15658 241210 15714 242010
rect 18418 241210 18474 242010
rect 21178 241210 21234 242010
rect 23938 241210 23994 242010
rect 26698 241210 26754 242010
rect 29458 241210 29514 242010
rect 32218 241210 32274 242010
rect 34978 241210 35034 242010
rect 37738 241210 37794 242010
rect 40498 241210 40554 242010
rect 43258 241210 43314 242010
rect 46018 241210 46074 242010
rect 48778 241210 48834 242010
rect 51538 241210 51594 242010
rect 54298 241210 54354 242010
rect 57058 241210 57114 242010
rect 59818 241210 59874 242010
rect 62578 241210 62634 242010
rect 65338 241210 65394 242010
rect 68558 241210 68614 242010
rect 71318 241210 71374 242010
rect 74078 241210 74134 242010
rect 76838 241210 76894 242010
rect 79598 241210 79654 242010
rect 82358 241210 82414 242010
rect 85118 241210 85174 242010
rect 87878 241210 87934 242010
rect 90638 241210 90694 242010
rect 93398 241210 93454 242010
rect 96158 241210 96214 242010
rect 98918 241210 98974 242010
rect 101678 241210 101734 242010
rect 104438 241210 104494 242010
rect 107198 241210 107254 242010
rect 109958 241210 110014 242010
rect 112718 241210 112774 242010
rect 115478 241210 115534 242010
rect 118238 241210 118294 242010
rect 120998 241210 121054 242010
rect 123758 241210 123814 242010
rect 126978 241210 127034 242010
rect 129738 241210 129794 242010
rect 132498 241210 132554 242010
rect 135258 241210 135314 242010
rect 138018 241210 138074 242010
rect 140778 241210 140834 242010
rect 143538 241210 143594 242010
rect 146298 241210 146354 242010
rect 149058 241210 149114 242010
rect 151818 241210 151874 242010
rect 154578 241210 154634 242010
rect 157338 241210 157394 242010
rect 160098 241210 160154 242010
rect 162858 241210 162914 242010
rect 165618 241210 165674 242010
rect 168378 241210 168434 242010
rect 171138 241210 171194 242010
rect 173898 241210 173954 242010
rect 176658 241210 176714 242010
rect 179418 241210 179474 242010
rect 182638 241210 182694 242010
rect 185398 241210 185454 242010
rect 188158 241210 188214 242010
rect 190918 241210 190974 242010
rect 193678 241210 193734 242010
rect 196438 241210 196494 242010
rect 199198 241210 199254 242010
rect 201958 241210 202014 242010
rect 204718 241210 204774 242010
rect 207478 241210 207534 242010
rect 210238 241210 210294 242010
rect 212998 241210 213054 242010
rect 215758 241210 215814 242010
rect 218518 241210 218574 242010
rect 221278 241210 221334 242010
rect 224038 241210 224094 242010
rect 226798 241210 226854 242010
rect 229558 241210 229614 242010
rect 232318 241210 232374 242010
rect 235078 241210 235134 242010
rect 237838 241210 237894 242010
rect 478 0 534 800
rect 3238 0 3294 800
rect 5998 0 6054 800
rect 8758 0 8814 800
rect 11518 0 11574 800
rect 14278 0 14334 800
rect 17038 0 17094 800
rect 19798 0 19854 800
rect 22558 0 22614 800
rect 25318 0 25374 800
rect 28078 0 28134 800
rect 30838 0 30894 800
rect 33598 0 33654 800
rect 36358 0 36414 800
rect 39118 0 39174 800
rect 41878 0 41934 800
rect 44638 0 44694 800
rect 47398 0 47454 800
rect 50158 0 50214 800
rect 52918 0 52974 800
rect 55678 0 55734 800
rect 58898 0 58954 800
rect 61658 0 61714 800
rect 64418 0 64474 800
rect 67178 0 67234 800
rect 69938 0 69994 800
rect 72698 0 72754 800
rect 75458 0 75514 800
rect 78218 0 78274 800
rect 80978 0 81034 800
rect 83738 0 83794 800
rect 86498 0 86554 800
rect 89258 0 89314 800
rect 92018 0 92074 800
rect 94778 0 94834 800
rect 97538 0 97594 800
rect 100298 0 100354 800
rect 103058 0 103114 800
rect 105818 0 105874 800
rect 108578 0 108634 800
rect 111338 0 111394 800
rect 114098 0 114154 800
rect 117318 0 117374 800
rect 120078 0 120134 800
rect 122838 0 122894 800
rect 125598 0 125654 800
rect 128358 0 128414 800
rect 131118 0 131174 800
rect 133878 0 133934 800
rect 136638 0 136694 800
rect 139398 0 139454 800
rect 142158 0 142214 800
rect 144918 0 144974 800
rect 147678 0 147734 800
rect 150438 0 150494 800
rect 153198 0 153254 800
rect 155958 0 156014 800
rect 158718 0 158774 800
rect 161478 0 161534 800
rect 164238 0 164294 800
rect 166998 0 167054 800
rect 169758 0 169814 800
rect 172978 0 173034 800
rect 175738 0 175794 800
rect 178498 0 178554 800
rect 181258 0 181314 800
rect 184018 0 184074 800
rect 186778 0 186834 800
rect 189538 0 189594 800
rect 192298 0 192354 800
rect 195058 0 195114 800
rect 197818 0 197874 800
rect 200578 0 200634 800
rect 203338 0 203394 800
rect 206098 0 206154 800
rect 208858 0 208914 800
rect 211618 0 211674 800
rect 214378 0 214434 800
rect 217138 0 217194 800
rect 219898 0 219954 800
rect 222658 0 222714 800
rect 225418 0 225474 800
rect 228178 0 228234 800
rect 231398 0 231454 800
rect 234158 0 234214 800
rect 236918 0 236974 800
<< obsm2 >>
rect 480 241154 1342 241210
rect 1510 241154 4102 241210
rect 4270 241154 6862 241210
rect 7030 241154 10082 241210
rect 10250 241154 12842 241210
rect 13010 241154 15602 241210
rect 15770 241154 18362 241210
rect 18530 241154 21122 241210
rect 21290 241154 23882 241210
rect 24050 241154 26642 241210
rect 26810 241154 29402 241210
rect 29570 241154 32162 241210
rect 32330 241154 34922 241210
rect 35090 241154 37682 241210
rect 37850 241154 40442 241210
rect 40610 241154 43202 241210
rect 43370 241154 45962 241210
rect 46130 241154 48722 241210
rect 48890 241154 51482 241210
rect 51650 241154 54242 241210
rect 54410 241154 57002 241210
rect 57170 241154 59762 241210
rect 59930 241154 62522 241210
rect 62690 241154 65282 241210
rect 65450 241154 68502 241210
rect 68670 241154 71262 241210
rect 71430 241154 74022 241210
rect 74190 241154 76782 241210
rect 76950 241154 79542 241210
rect 79710 241154 82302 241210
rect 82470 241154 85062 241210
rect 85230 241154 87822 241210
rect 87990 241154 90582 241210
rect 90750 241154 93342 241210
rect 93510 241154 96102 241210
rect 96270 241154 98862 241210
rect 99030 241154 101622 241210
rect 101790 241154 104382 241210
rect 104550 241154 107142 241210
rect 107310 241154 109902 241210
rect 110070 241154 112662 241210
rect 112830 241154 115422 241210
rect 115590 241154 118182 241210
rect 118350 241154 120942 241210
rect 121110 241154 123702 241210
rect 123870 241154 126922 241210
rect 127090 241154 129682 241210
rect 129850 241154 132442 241210
rect 132610 241154 135202 241210
rect 135370 241154 137962 241210
rect 138130 241154 140722 241210
rect 140890 241154 143482 241210
rect 143650 241154 146242 241210
rect 146410 241154 149002 241210
rect 149170 241154 151762 241210
rect 151930 241154 154522 241210
rect 154690 241154 157282 241210
rect 157450 241154 160042 241210
rect 160210 241154 162802 241210
rect 162970 241154 165562 241210
rect 165730 241154 168322 241210
rect 168490 241154 171082 241210
rect 171250 241154 173842 241210
rect 174010 241154 176602 241210
rect 176770 241154 179362 241210
rect 179530 241154 182582 241210
rect 182750 241154 185342 241210
rect 185510 241154 188102 241210
rect 188270 241154 190862 241210
rect 191030 241154 193622 241210
rect 193790 241154 196382 241210
rect 196550 241154 199142 241210
rect 199310 241154 201902 241210
rect 202070 241154 204662 241210
rect 204830 241154 207422 241210
rect 207590 241154 210182 241210
rect 210350 241154 212942 241210
rect 213110 241154 215702 241210
rect 215870 241154 218462 241210
rect 218630 241154 221222 241210
rect 221390 241154 223982 241210
rect 224150 241154 226742 241210
rect 226910 241154 229502 241210
rect 229670 241154 232262 241210
rect 232430 241154 235022 241210
rect 235190 241154 237782 241210
rect 237950 241154 238078 241210
rect 480 856 238078 241154
rect 590 711 3182 856
rect 3350 711 5942 856
rect 6110 711 8702 856
rect 8870 711 11462 856
rect 11630 711 14222 856
rect 14390 711 16982 856
rect 17150 711 19742 856
rect 19910 711 22502 856
rect 22670 711 25262 856
rect 25430 711 28022 856
rect 28190 711 30782 856
rect 30950 711 33542 856
rect 33710 711 36302 856
rect 36470 711 39062 856
rect 39230 711 41822 856
rect 41990 711 44582 856
rect 44750 711 47342 856
rect 47510 711 50102 856
rect 50270 711 52862 856
rect 53030 711 55622 856
rect 55790 711 58842 856
rect 59010 711 61602 856
rect 61770 711 64362 856
rect 64530 711 67122 856
rect 67290 711 69882 856
rect 70050 711 72642 856
rect 72810 711 75402 856
rect 75570 711 78162 856
rect 78330 711 80922 856
rect 81090 711 83682 856
rect 83850 711 86442 856
rect 86610 711 89202 856
rect 89370 711 91962 856
rect 92130 711 94722 856
rect 94890 711 97482 856
rect 97650 711 100242 856
rect 100410 711 103002 856
rect 103170 711 105762 856
rect 105930 711 108522 856
rect 108690 711 111282 856
rect 111450 711 114042 856
rect 114210 711 117262 856
rect 117430 711 120022 856
rect 120190 711 122782 856
rect 122950 711 125542 856
rect 125710 711 128302 856
rect 128470 711 131062 856
rect 131230 711 133822 856
rect 133990 711 136582 856
rect 136750 711 139342 856
rect 139510 711 142102 856
rect 142270 711 144862 856
rect 145030 711 147622 856
rect 147790 711 150382 856
rect 150550 711 153142 856
rect 153310 711 155902 856
rect 156070 711 158662 856
rect 158830 711 161422 856
rect 161590 711 164182 856
rect 164350 711 166942 856
rect 167110 711 169702 856
rect 169870 711 172922 856
rect 173090 711 175682 856
rect 175850 711 178442 856
rect 178610 711 181202 856
rect 181370 711 183962 856
rect 184130 711 186722 856
rect 186890 711 189482 856
rect 189650 711 192242 856
rect 192410 711 195002 856
rect 195170 711 197762 856
rect 197930 711 200522 856
rect 200690 711 203282 856
rect 203450 711 206042 856
rect 206210 711 208802 856
rect 208970 711 211562 856
rect 211730 711 214322 856
rect 214490 711 217082 856
rect 217250 711 219842 856
rect 220010 711 222602 856
rect 222770 711 225362 856
rect 225530 711 228122 856
rect 228290 711 231342 856
rect 231510 711 234102 856
rect 234270 711 236862 856
rect 237030 711 238078 856
<< metal3 >>
rect 0 238688 800 238808
rect 239066 238688 239866 238808
rect 0 234608 800 234728
rect 239066 234608 239866 234728
rect 0 230528 800 230648
rect 239066 230528 239866 230648
rect 0 226448 800 226568
rect 239066 226448 239866 226568
rect 0 222368 800 222488
rect 239066 222368 239866 222488
rect 0 218288 800 218408
rect 239066 218288 239866 218408
rect 0 214208 800 214328
rect 239066 214208 239866 214328
rect 0 210128 800 210248
rect 239066 210128 239866 210248
rect 0 206048 800 206168
rect 239066 206048 239866 206168
rect 0 201968 800 202088
rect 239066 201968 239866 202088
rect 0 197888 800 198008
rect 239066 197888 239866 198008
rect 0 193808 800 193928
rect 239066 193808 239866 193928
rect 0 189728 800 189848
rect 239066 189728 239866 189848
rect 0 185648 800 185768
rect 239066 185648 239866 185768
rect 0 181568 800 181688
rect 239066 181568 239866 181688
rect 0 177488 800 177608
rect 239066 177488 239866 177608
rect 0 173408 800 173528
rect 239066 173408 239866 173528
rect 239066 169328 239866 169448
rect 0 168648 800 168768
rect 239066 165248 239866 165368
rect 0 164568 800 164688
rect 239066 161168 239866 161288
rect 0 160488 800 160608
rect 239066 157088 239866 157208
rect 0 156408 800 156528
rect 0 152328 800 152448
rect 239066 152328 239866 152448
rect 0 148248 800 148368
rect 239066 148248 239866 148368
rect 0 144168 800 144288
rect 239066 144168 239866 144288
rect 0 140088 800 140208
rect 239066 140088 239866 140208
rect 0 136008 800 136128
rect 239066 136008 239866 136128
rect 0 131928 800 132048
rect 239066 131928 239866 132048
rect 0 127848 800 127968
rect 239066 127848 239866 127968
rect 0 123768 800 123888
rect 239066 123768 239866 123888
rect 0 119688 800 119808
rect 239066 119688 239866 119808
rect 0 115608 800 115728
rect 239066 115608 239866 115728
rect 0 111528 800 111648
rect 239066 111528 239866 111648
rect 0 107448 800 107568
rect 239066 107448 239866 107568
rect 0 103368 800 103488
rect 239066 103368 239866 103488
rect 0 99288 800 99408
rect 239066 99288 239866 99408
rect 0 95208 800 95328
rect 239066 95208 239866 95328
rect 0 91128 800 91248
rect 239066 91128 239866 91248
rect 0 87048 800 87168
rect 239066 87048 239866 87168
rect 239066 82968 239866 83088
rect 0 82288 800 82408
rect 239066 78888 239866 79008
rect 0 78208 800 78328
rect 239066 74808 239866 74928
rect 0 74128 800 74248
rect 0 70048 800 70168
rect 239066 70048 239866 70168
rect 0 65968 800 66088
rect 239066 65968 239866 66088
rect 0 61888 800 62008
rect 239066 61888 239866 62008
rect 0 57808 800 57928
rect 239066 57808 239866 57928
rect 0 53728 800 53848
rect 239066 53728 239866 53848
rect 0 49648 800 49768
rect 239066 49648 239866 49768
rect 0 45568 800 45688
rect 239066 45568 239866 45688
rect 0 41488 800 41608
rect 239066 41488 239866 41608
rect 0 37408 800 37528
rect 239066 37408 239866 37528
rect 0 33328 800 33448
rect 239066 33328 239866 33448
rect 0 29248 800 29368
rect 239066 29248 239866 29368
rect 0 25168 800 25288
rect 239066 25168 239866 25288
rect 0 21088 800 21208
rect 239066 21088 239866 21208
rect 0 17008 800 17128
rect 239066 17008 239866 17128
rect 0 12928 800 13048
rect 239066 12928 239866 13048
rect 0 8848 800 8968
rect 239066 8848 239866 8968
rect 0 4768 800 4888
rect 239066 4768 239866 4888
rect 239066 688 239866 808
<< obsm3 >>
rect 800 238888 239066 239597
rect 880 238608 238986 238888
rect 800 234808 239066 238608
rect 880 234528 238986 234808
rect 800 230728 239066 234528
rect 880 230448 238986 230728
rect 800 226648 239066 230448
rect 880 226368 238986 226648
rect 800 222568 239066 226368
rect 880 222288 238986 222568
rect 800 218488 239066 222288
rect 880 218208 238986 218488
rect 800 214408 239066 218208
rect 880 214128 238986 214408
rect 800 210328 239066 214128
rect 880 210048 238986 210328
rect 800 206248 239066 210048
rect 880 205968 238986 206248
rect 800 202168 239066 205968
rect 880 201888 238986 202168
rect 800 198088 239066 201888
rect 880 197808 238986 198088
rect 800 194008 239066 197808
rect 880 193728 238986 194008
rect 800 189928 239066 193728
rect 880 189648 238986 189928
rect 800 185848 239066 189648
rect 880 185568 238986 185848
rect 800 181768 239066 185568
rect 880 181488 238986 181768
rect 800 177688 239066 181488
rect 880 177408 238986 177688
rect 800 173608 239066 177408
rect 880 173328 238986 173608
rect 800 169528 239066 173328
rect 800 169248 238986 169528
rect 800 168848 239066 169248
rect 880 168568 239066 168848
rect 800 165448 239066 168568
rect 800 165168 238986 165448
rect 800 164768 239066 165168
rect 880 164488 239066 164768
rect 800 161368 239066 164488
rect 800 161088 238986 161368
rect 800 160688 239066 161088
rect 880 160408 239066 160688
rect 800 157288 239066 160408
rect 800 157008 238986 157288
rect 800 156608 239066 157008
rect 880 156328 239066 156608
rect 800 152528 239066 156328
rect 880 152248 238986 152528
rect 800 148448 239066 152248
rect 880 148168 238986 148448
rect 800 144368 239066 148168
rect 880 144088 238986 144368
rect 800 140288 239066 144088
rect 880 140008 238986 140288
rect 800 136208 239066 140008
rect 880 135928 238986 136208
rect 800 132128 239066 135928
rect 880 131848 238986 132128
rect 800 128048 239066 131848
rect 880 127768 238986 128048
rect 800 123968 239066 127768
rect 880 123688 238986 123968
rect 800 119888 239066 123688
rect 880 119608 238986 119888
rect 800 115808 239066 119608
rect 880 115528 238986 115808
rect 800 111728 239066 115528
rect 880 111448 238986 111728
rect 800 107648 239066 111448
rect 880 107368 238986 107648
rect 800 103568 239066 107368
rect 880 103288 238986 103568
rect 800 99488 239066 103288
rect 880 99208 238986 99488
rect 800 95408 239066 99208
rect 880 95128 238986 95408
rect 800 91328 239066 95128
rect 880 91048 238986 91328
rect 800 87248 239066 91048
rect 880 86968 238986 87248
rect 800 83168 239066 86968
rect 800 82888 238986 83168
rect 800 82488 239066 82888
rect 880 82208 239066 82488
rect 800 79088 239066 82208
rect 800 78808 238986 79088
rect 800 78408 239066 78808
rect 880 78128 239066 78408
rect 800 75008 239066 78128
rect 800 74728 238986 75008
rect 800 74328 239066 74728
rect 880 74048 239066 74328
rect 800 70248 239066 74048
rect 880 69968 238986 70248
rect 800 66168 239066 69968
rect 880 65888 238986 66168
rect 800 62088 239066 65888
rect 880 61808 238986 62088
rect 800 58008 239066 61808
rect 880 57728 238986 58008
rect 800 53928 239066 57728
rect 880 53648 238986 53928
rect 800 49848 239066 53648
rect 880 49568 238986 49848
rect 800 45768 239066 49568
rect 880 45488 238986 45768
rect 800 41688 239066 45488
rect 880 41408 238986 41688
rect 800 37608 239066 41408
rect 880 37328 238986 37608
rect 800 33528 239066 37328
rect 880 33248 238986 33528
rect 800 29448 239066 33248
rect 880 29168 238986 29448
rect 800 25368 239066 29168
rect 880 25088 238986 25368
rect 800 21288 239066 25088
rect 880 21008 238986 21288
rect 800 17208 239066 21008
rect 880 16928 238986 17208
rect 800 13128 239066 16928
rect 880 12848 238986 13128
rect 800 9048 239066 12848
rect 880 8768 238986 9048
rect 800 4968 239066 8768
rect 880 4688 238986 4968
rect 800 888 239066 4688
rect 800 715 238986 888
<< metal4 >>
rect 4208 2128 4528 239408
rect 9208 2128 9528 239408
rect 14208 2128 14528 239408
rect 19208 2128 19528 239408
rect 24208 2128 24528 239408
rect 29208 2128 29528 239408
rect 34208 218452 34528 239408
rect 39208 218452 39528 239408
rect 44208 218452 44528 239408
rect 49208 218452 49528 239408
rect 54208 218452 54528 239408
rect 59208 218452 59528 239408
rect 64208 218452 64528 239408
rect 69208 218452 69528 239408
rect 74208 218452 74528 239408
rect 79208 218452 79528 239408
rect 84208 218452 84528 239408
rect 89208 218452 89528 239408
rect 94208 218452 94528 239408
rect 99208 218452 99528 239408
rect 104208 218452 104528 239408
rect 109208 218452 109528 239408
rect 114208 218452 114528 239408
rect 119208 218452 119528 239408
rect 124208 218452 124528 239408
rect 129208 218452 129528 239408
rect 34208 2128 34528 137048
rect 39208 2128 39528 137048
rect 44208 2128 44528 137048
rect 49208 2128 49528 137048
rect 54208 2128 54528 137048
rect 59208 2128 59528 137048
rect 64208 2128 64528 137048
rect 69208 2128 69528 137048
rect 74208 2128 74528 137048
rect 79208 2128 79528 137048
rect 84208 2128 84528 137048
rect 89208 2128 89528 137048
rect 94208 2128 94528 137048
rect 99208 2128 99528 137048
rect 104208 2128 104528 137048
rect 109208 2128 109528 137048
rect 114208 2128 114528 137048
rect 119208 2128 119528 137048
rect 124208 2128 124528 137048
rect 129208 2128 129528 137048
rect 134208 2128 134528 239408
rect 139208 2128 139528 239408
rect 144208 2128 144528 239408
rect 149208 2128 149528 239408
rect 154208 2128 154528 239408
rect 159208 2128 159528 239408
rect 164208 2128 164528 239408
rect 169208 2128 169528 239408
rect 174208 2128 174528 239408
rect 179208 2128 179528 239408
rect 184208 2128 184528 239408
rect 189208 2128 189528 239408
rect 194208 2128 194528 239408
rect 199208 2128 199528 239408
rect 204208 2128 204528 239408
rect 209208 2128 209528 239408
rect 214208 2128 214528 239408
rect 219208 2128 219528 239408
rect 224208 2128 224528 239408
rect 229208 2128 229528 239408
rect 234208 2128 234528 239408
<< obsm4 >>
rect 33731 239488 171245 239597
rect 33731 218372 34128 239488
rect 34608 218372 39128 239488
rect 39608 218372 44128 239488
rect 44608 218372 49128 239488
rect 49608 218372 54128 239488
rect 54608 218372 59128 239488
rect 59608 218372 64128 239488
rect 64608 218372 69128 239488
rect 69608 218372 74128 239488
rect 74608 218372 79128 239488
rect 79608 218372 84128 239488
rect 84608 218372 89128 239488
rect 89608 218372 94128 239488
rect 94608 218372 99128 239488
rect 99608 218372 104128 239488
rect 104608 218372 109128 239488
rect 109608 218372 114128 239488
rect 114608 218372 119128 239488
rect 119608 218372 124128 239488
rect 124608 218372 129128 239488
rect 129608 218372 134128 239488
rect 33731 137128 134128 218372
rect 33731 2048 34128 137128
rect 34608 2048 39128 137128
rect 39608 2048 44128 137128
rect 44608 2048 49128 137128
rect 49608 2048 54128 137128
rect 54608 2048 59128 137128
rect 59608 2048 64128 137128
rect 64608 2048 69128 137128
rect 69608 2048 74128 137128
rect 74608 2048 79128 137128
rect 79608 2048 84128 137128
rect 84608 2048 89128 137128
rect 89608 2048 94128 137128
rect 94608 2048 99128 137128
rect 99608 2048 104128 137128
rect 104608 2048 109128 137128
rect 109608 2048 114128 137128
rect 114608 2048 119128 137128
rect 119608 2048 124128 137128
rect 124608 2048 129128 137128
rect 129608 2048 134128 137128
rect 134608 2048 139128 239488
rect 139608 2048 144128 239488
rect 144608 2048 149128 239488
rect 149608 2048 154128 239488
rect 154608 2048 159128 239488
rect 159608 2048 164128 239488
rect 164608 2048 169128 239488
rect 169608 2048 171245 239488
rect 33731 1667 171245 2048
<< metal5 >>
rect 1104 235068 238740 235388
rect 1104 219750 238740 220070
rect 1104 204432 238740 204752
rect 1104 189114 238740 189434
rect 1104 173796 238740 174116
rect 1104 158478 238740 158798
rect 1104 143160 238740 143480
rect 1104 127842 238740 128162
rect 1104 112524 238740 112844
rect 1104 97206 238740 97526
rect 1104 81888 238740 82208
rect 1104 66570 238740 66890
rect 1104 51252 238740 51572
rect 1104 35934 238740 36254
rect 1104 20616 238740 20936
rect 1104 5298 238740 5618
<< labels >>
rlabel metal2 s 29458 241210 29514 242010 6 clk_i
port 1 nsew signal input
rlabel metal3 s 239066 185648 239866 185768 6 debug_req_i
port 2 nsew signal input
rlabel metal2 s 232318 241210 232374 242010 6 eFPGA_delay_o[0]
port 3 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 eFPGA_delay_o[1]
port 4 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 eFPGA_delay_o[2]
port 5 nsew signal output
rlabel metal2 s 171138 241210 171194 242010 6 eFPGA_delay_o[3]
port 6 nsew signal output
rlabel metal2 s 87878 241210 87934 242010 6 eFPGA_en_o
port 7 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 eFPGA_fpga_done_i
port 8 nsew signal input
rlabel metal3 s 239066 177488 239866 177608 6 eFPGA_operand_a_o[0]
port 9 nsew signal output
rlabel metal3 s 239066 65968 239866 66088 6 eFPGA_operand_a_o[10]
port 10 nsew signal output
rlabel metal3 s 0 230528 800 230648 6 eFPGA_operand_a_o[11]
port 11 nsew signal output
rlabel metal2 s 146298 241210 146354 242010 6 eFPGA_operand_a_o[12]
port 12 nsew signal output
rlabel metal2 s 101678 241210 101734 242010 6 eFPGA_operand_a_o[13]
port 13 nsew signal output
rlabel metal3 s 239066 107448 239866 107568 6 eFPGA_operand_a_o[14]
port 14 nsew signal output
rlabel metal3 s 0 193808 800 193928 6 eFPGA_operand_a_o[15]
port 15 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 eFPGA_operand_a_o[16]
port 16 nsew signal output
rlabel metal3 s 239066 123768 239866 123888 6 eFPGA_operand_a_o[17]
port 17 nsew signal output
rlabel metal2 s 1398 241210 1454 242010 6 eFPGA_operand_a_o[18]
port 18 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 eFPGA_operand_a_o[19]
port 19 nsew signal output
rlabel metal2 s 15658 241210 15714 242010 6 eFPGA_operand_a_o[1]
port 20 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 eFPGA_operand_a_o[20]
port 21 nsew signal output
rlabel metal3 s 239066 161168 239866 161288 6 eFPGA_operand_a_o[21]
port 22 nsew signal output
rlabel metal3 s 239066 37408 239866 37528 6 eFPGA_operand_a_o[22]
port 23 nsew signal output
rlabel metal3 s 239066 140088 239866 140208 6 eFPGA_operand_a_o[23]
port 24 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 eFPGA_operand_a_o[24]
port 25 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 eFPGA_operand_a_o[25]
port 26 nsew signal output
rlabel metal3 s 239066 17008 239866 17128 6 eFPGA_operand_a_o[26]
port 27 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 eFPGA_operand_a_o[27]
port 28 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 eFPGA_operand_a_o[28]
port 29 nsew signal output
rlabel metal2 s 165618 241210 165674 242010 6 eFPGA_operand_a_o[29]
port 30 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 eFPGA_operand_a_o[2]
port 31 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 eFPGA_operand_a_o[30]
port 32 nsew signal output
rlabel metal2 s 18418 241210 18474 242010 6 eFPGA_operand_a_o[31]
port 33 nsew signal output
rlabel metal2 s 179418 241210 179474 242010 6 eFPGA_operand_a_o[3]
port 34 nsew signal output
rlabel metal2 s 40498 241210 40554 242010 6 eFPGA_operand_a_o[4]
port 35 nsew signal output
rlabel metal2 s 221278 241210 221334 242010 6 eFPGA_operand_a_o[5]
port 36 nsew signal output
rlabel metal2 s 93398 241210 93454 242010 6 eFPGA_operand_a_o[6]
port 37 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 eFPGA_operand_a_o[7]
port 38 nsew signal output
rlabel metal2 s 157338 241210 157394 242010 6 eFPGA_operand_a_o[8]
port 39 nsew signal output
rlabel metal2 s 109958 241210 110014 242010 6 eFPGA_operand_a_o[9]
port 40 nsew signal output
rlabel metal2 s 189538 0 189594 800 6 eFPGA_operand_b_o[0]
port 41 nsew signal output
rlabel metal3 s 239066 87048 239866 87168 6 eFPGA_operand_b_o[10]
port 42 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 eFPGA_operand_b_o[11]
port 43 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 eFPGA_operand_b_o[12]
port 44 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 eFPGA_operand_b_o[13]
port 45 nsew signal output
rlabel metal2 s 4158 241210 4214 242010 6 eFPGA_operand_b_o[14]
port 46 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 eFPGA_operand_b_o[15]
port 47 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 eFPGA_operand_b_o[16]
port 48 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 eFPGA_operand_b_o[17]
port 49 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 eFPGA_operand_b_o[18]
port 50 nsew signal output
rlabel metal2 s 234158 0 234214 800 6 eFPGA_operand_b_o[19]
port 51 nsew signal output
rlabel metal2 s 196438 241210 196494 242010 6 eFPGA_operand_b_o[1]
port 52 nsew signal output
rlabel metal2 s 85118 241210 85174 242010 6 eFPGA_operand_b_o[20]
port 53 nsew signal output
rlabel metal2 s 96158 241210 96214 242010 6 eFPGA_operand_b_o[21]
port 54 nsew signal output
rlabel metal2 s 229558 241210 229614 242010 6 eFPGA_operand_b_o[22]
port 55 nsew signal output
rlabel metal3 s 239066 234608 239866 234728 6 eFPGA_operand_b_o[23]
port 56 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 eFPGA_operand_b_o[24]
port 57 nsew signal output
rlabel metal2 s 126978 241210 127034 242010 6 eFPGA_operand_b_o[25]
port 58 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 eFPGA_operand_b_o[26]
port 59 nsew signal output
rlabel metal3 s 239066 181568 239866 181688 6 eFPGA_operand_b_o[27]
port 60 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 eFPGA_operand_b_o[28]
port 61 nsew signal output
rlabel metal3 s 239066 165248 239866 165368 6 eFPGA_operand_b_o[29]
port 62 nsew signal output
rlabel metal2 s 57058 241210 57114 242010 6 eFPGA_operand_b_o[2]
port 63 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 eFPGA_operand_b_o[30]
port 64 nsew signal output
rlabel metal3 s 239066 70048 239866 70168 6 eFPGA_operand_b_o[31]
port 65 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 eFPGA_operand_b_o[3]
port 66 nsew signal output
rlabel metal3 s 0 181568 800 181688 6 eFPGA_operand_b_o[4]
port 67 nsew signal output
rlabel metal3 s 239066 111528 239866 111648 6 eFPGA_operand_b_o[5]
port 68 nsew signal output
rlabel metal2 s 154578 241210 154634 242010 6 eFPGA_operand_b_o[6]
port 69 nsew signal output
rlabel metal2 s 204718 241210 204774 242010 6 eFPGA_operand_b_o[7]
port 70 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 eFPGA_operand_b_o[8]
port 71 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 eFPGA_operand_b_o[9]
port 72 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 eFPGA_operator_o[0]
port 73 nsew signal output
rlabel metal2 s 21178 241210 21234 242010 6 eFPGA_operator_o[1]
port 74 nsew signal output
rlabel metal2 s 34978 241210 35034 242010 6 eFPGA_result_a_i[0]
port 75 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 eFPGA_result_a_i[10]
port 76 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 eFPGA_result_a_i[11]
port 77 nsew signal input
rlabel metal3 s 0 214208 800 214328 6 eFPGA_result_a_i[12]
port 78 nsew signal input
rlabel metal3 s 239066 218288 239866 218408 6 eFPGA_result_a_i[13]
port 79 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 eFPGA_result_a_i[14]
port 80 nsew signal input
rlabel metal3 s 239066 61888 239866 62008 6 eFPGA_result_a_i[15]
port 81 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 eFPGA_result_a_i[16]
port 82 nsew signal input
rlabel metal2 s 182638 241210 182694 242010 6 eFPGA_result_a_i[17]
port 83 nsew signal input
rlabel metal2 s 54298 241210 54354 242010 6 eFPGA_result_a_i[18]
port 84 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 eFPGA_result_a_i[19]
port 85 nsew signal input
rlabel metal3 s 239066 173408 239866 173528 6 eFPGA_result_a_i[1]
port 86 nsew signal input
rlabel metal2 s 201958 241210 202014 242010 6 eFPGA_result_a_i[20]
port 87 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 eFPGA_result_a_i[21]
port 88 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 eFPGA_result_a_i[22]
port 89 nsew signal input
rlabel metal3 s 239066 21088 239866 21208 6 eFPGA_result_a_i[23]
port 90 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 eFPGA_result_a_i[24]
port 91 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 eFPGA_result_a_i[25]
port 92 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 eFPGA_result_a_i[26]
port 93 nsew signal input
rlabel metal2 s 65338 241210 65394 242010 6 eFPGA_result_a_i[27]
port 94 nsew signal input
rlabel metal3 s 0 197888 800 198008 6 eFPGA_result_a_i[28]
port 95 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 eFPGA_result_a_i[29]
port 96 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 eFPGA_result_a_i[2]
port 97 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 eFPGA_result_a_i[30]
port 98 nsew signal input
rlabel metal2 s 115478 241210 115534 242010 6 eFPGA_result_a_i[31]
port 99 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 eFPGA_result_a_i[3]
port 100 nsew signal input
rlabel metal2 s 188158 241210 188214 242010 6 eFPGA_result_a_i[4]
port 101 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 eFPGA_result_a_i[5]
port 102 nsew signal input
rlabel metal3 s 0 210128 800 210248 6 eFPGA_result_a_i[6]
port 103 nsew signal input
rlabel metal3 s 239066 136008 239866 136128 6 eFPGA_result_a_i[7]
port 104 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 eFPGA_result_a_i[8]
port 105 nsew signal input
rlabel metal2 s 215758 241210 215814 242010 6 eFPGA_result_a_i[9]
port 106 nsew signal input
rlabel metal2 s 46018 241210 46074 242010 6 eFPGA_result_b_i[0]
port 107 nsew signal input
rlabel metal3 s 239066 33328 239866 33448 6 eFPGA_result_b_i[10]
port 108 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 eFPGA_result_b_i[11]
port 109 nsew signal input
rlabel metal2 s 199198 241210 199254 242010 6 eFPGA_result_b_i[12]
port 110 nsew signal input
rlabel metal3 s 239066 103368 239866 103488 6 eFPGA_result_b_i[13]
port 111 nsew signal input
rlabel metal2 s 98918 241210 98974 242010 6 eFPGA_result_b_i[14]
port 112 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 eFPGA_result_b_i[15]
port 113 nsew signal input
rlabel metal3 s 239066 230528 239866 230648 6 eFPGA_result_b_i[16]
port 114 nsew signal input
rlabel metal2 s 62578 241210 62634 242010 6 eFPGA_result_b_i[17]
port 115 nsew signal input
rlabel metal3 s 239066 25168 239866 25288 6 eFPGA_result_b_i[18]
port 116 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 eFPGA_result_b_i[19]
port 117 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 eFPGA_result_b_i[1]
port 118 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 eFPGA_result_b_i[20]
port 119 nsew signal input
rlabel metal2 s 90638 241210 90694 242010 6 eFPGA_result_b_i[21]
port 120 nsew signal input
rlabel metal3 s 0 238688 800 238808 6 eFPGA_result_b_i[22]
port 121 nsew signal input
rlabel metal3 s 239066 222368 239866 222488 6 eFPGA_result_b_i[23]
port 122 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 eFPGA_result_b_i[24]
port 123 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 eFPGA_result_b_i[25]
port 124 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 eFPGA_result_b_i[26]
port 125 nsew signal input
rlabel metal2 s 190918 241210 190974 242010 6 eFPGA_result_b_i[27]
port 126 nsew signal input
rlabel metal3 s 239066 115608 239866 115728 6 eFPGA_result_b_i[28]
port 127 nsew signal input
rlabel metal3 s 239066 193808 239866 193928 6 eFPGA_result_b_i[29]
port 128 nsew signal input
rlabel metal3 s 239066 201968 239866 202088 6 eFPGA_result_b_i[2]
port 129 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 eFPGA_result_b_i[30]
port 130 nsew signal input
rlabel metal2 s 10138 241210 10194 242010 6 eFPGA_result_b_i[31]
port 131 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 eFPGA_result_b_i[3]
port 132 nsew signal input
rlabel metal3 s 239066 8848 239866 8968 6 eFPGA_result_b_i[4]
port 133 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 eFPGA_result_b_i[5]
port 134 nsew signal input
rlabel metal2 s 181258 0 181314 800 6 eFPGA_result_b_i[6]
port 135 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 eFPGA_result_b_i[7]
port 136 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 eFPGA_result_b_i[8]
port 137 nsew signal input
rlabel metal3 s 0 226448 800 226568 6 eFPGA_result_b_i[9]
port 138 nsew signal input
rlabel metal2 s 132498 241210 132554 242010 6 eFPGA_result_c_i[0]
port 139 nsew signal input
rlabel metal2 s 176658 241210 176714 242010 6 eFPGA_result_c_i[10]
port 140 nsew signal input
rlabel metal2 s 68558 241210 68614 242010 6 eFPGA_result_c_i[11]
port 141 nsew signal input
rlabel metal2 s 162858 241210 162914 242010 6 eFPGA_result_c_i[12]
port 142 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 eFPGA_result_c_i[13]
port 143 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 eFPGA_result_c_i[14]
port 144 nsew signal input
rlabel metal2 s 168378 241210 168434 242010 6 eFPGA_result_c_i[15]
port 145 nsew signal input
rlabel metal2 s 140778 241210 140834 242010 6 eFPGA_result_c_i[16]
port 146 nsew signal input
rlabel metal2 s 23938 241210 23994 242010 6 eFPGA_result_c_i[17]
port 147 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 eFPGA_result_c_i[18]
port 148 nsew signal input
rlabel metal3 s 239066 119688 239866 119808 6 eFPGA_result_c_i[19]
port 149 nsew signal input
rlabel metal3 s 239066 148248 239866 148368 6 eFPGA_result_c_i[1]
port 150 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 eFPGA_result_c_i[20]
port 151 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 eFPGA_result_c_i[21]
port 152 nsew signal input
rlabel metal2 s 226798 241210 226854 242010 6 eFPGA_result_c_i[22]
port 153 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 eFPGA_result_c_i[23]
port 154 nsew signal input
rlabel metal3 s 239066 169328 239866 169448 6 eFPGA_result_c_i[24]
port 155 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 eFPGA_result_c_i[25]
port 156 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 eFPGA_result_c_i[26]
port 157 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 eFPGA_result_c_i[27]
port 158 nsew signal input
rlabel metal2 s 160098 241210 160154 242010 6 eFPGA_result_c_i[28]
port 159 nsew signal input
rlabel metal2 s 71318 241210 71374 242010 6 eFPGA_result_c_i[29]
port 160 nsew signal input
rlabel metal2 s 32218 241210 32274 242010 6 eFPGA_result_c_i[2]
port 161 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 eFPGA_result_c_i[30]
port 162 nsew signal input
rlabel metal3 s 239066 78888 239866 79008 6 eFPGA_result_c_i[31]
port 163 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 eFPGA_result_c_i[3]
port 164 nsew signal input
rlabel metal2 s 51538 241210 51594 242010 6 eFPGA_result_c_i[4]
port 165 nsew signal input
rlabel metal3 s 0 201968 800 202088 6 eFPGA_result_c_i[5]
port 166 nsew signal input
rlabel metal3 s 239066 91128 239866 91248 6 eFPGA_result_c_i[6]
port 167 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 eFPGA_result_c_i[7]
port 168 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 eFPGA_result_c_i[8]
port 169 nsew signal input
rlabel metal2 s 74078 241210 74134 242010 6 eFPGA_result_c_i[9]
port 170 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 eFPGA_write_strobe_o
port 171 nsew signal output
rlabel metal2 s 76838 241210 76894 242010 6 ext_data_addr_i[0]
port 172 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 ext_data_addr_i[10]
port 173 nsew signal input
rlabel metal3 s 239066 688 239866 808 6 ext_data_addr_i[11]
port 174 nsew signal input
rlabel metal2 s 79598 241210 79654 242010 6 ext_data_addr_i[12]
port 175 nsew signal input
rlabel metal2 s 118238 241210 118294 242010 6 ext_data_addr_i[13]
port 176 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 ext_data_addr_i[14]
port 177 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 ext_data_addr_i[15]
port 178 nsew signal input
rlabel metal2 s 107198 241210 107254 242010 6 ext_data_addr_i[16]
port 179 nsew signal input
rlabel metal3 s 239066 74808 239866 74928 6 ext_data_addr_i[17]
port 180 nsew signal input
rlabel metal3 s 239066 157088 239866 157208 6 ext_data_addr_i[18]
port 181 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 ext_data_addr_i[19]
port 182 nsew signal input
rlabel metal3 s 0 189728 800 189848 6 ext_data_addr_i[1]
port 183 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 ext_data_addr_i[20]
port 184 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 ext_data_addr_i[21]
port 185 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 ext_data_addr_i[22]
port 186 nsew signal input
rlabel metal2 s 129738 241210 129794 242010 6 ext_data_addr_i[23]
port 187 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 ext_data_addr_i[24]
port 188 nsew signal input
rlabel metal3 s 239066 49648 239866 49768 6 ext_data_addr_i[25]
port 189 nsew signal input
rlabel metal2 s 224038 241210 224094 242010 6 ext_data_addr_i[26]
port 190 nsew signal input
rlabel metal2 s 200578 0 200634 800 6 ext_data_addr_i[27]
port 191 nsew signal input
rlabel metal2 s 48778 241210 48834 242010 6 ext_data_addr_i[28]
port 192 nsew signal input
rlabel metal2 s 236918 0 236974 800 6 ext_data_addr_i[29]
port 193 nsew signal input
rlabel metal2 s 135258 241210 135314 242010 6 ext_data_addr_i[2]
port 194 nsew signal input
rlabel metal3 s 0 234608 800 234728 6 ext_data_addr_i[30]
port 195 nsew signal input
rlabel metal2 s 82358 241210 82414 242010 6 ext_data_addr_i[31]
port 196 nsew signal input
rlabel metal2 s 478 0 534 800 6 ext_data_addr_i[3]
port 197 nsew signal input
rlabel metal2 s 59818 241210 59874 242010 6 ext_data_addr_i[4]
port 198 nsew signal input
rlabel metal3 s 0 218288 800 218408 6 ext_data_addr_i[5]
port 199 nsew signal input
rlabel metal2 s 185398 241210 185454 242010 6 ext_data_addr_i[6]
port 200 nsew signal input
rlabel metal2 s 43258 241210 43314 242010 6 ext_data_addr_i[7]
port 201 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 ext_data_addr_i[8]
port 202 nsew signal input
rlabel metal3 s 0 206048 800 206168 6 ext_data_addr_i[9]
port 203 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 ext_data_be_i[0]
port 204 nsew signal input
rlabel metal2 s 26698 241210 26754 242010 6 ext_data_be_i[1]
port 205 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 ext_data_be_i[2]
port 206 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 ext_data_be_i[3]
port 207 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 ext_data_gnt_o
port 208 nsew signal output
rlabel metal3 s 239066 226448 239866 226568 6 ext_data_rdata_o[0]
port 209 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 ext_data_rdata_o[10]
port 210 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 ext_data_rdata_o[11]
port 211 nsew signal output
rlabel metal2 s 178498 0 178554 800 6 ext_data_rdata_o[12]
port 212 nsew signal output
rlabel metal3 s 239066 57808 239866 57928 6 ext_data_rdata_o[13]
port 213 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 ext_data_rdata_o[14]
port 214 nsew signal output
rlabel metal2 s 104438 241210 104494 242010 6 ext_data_rdata_o[15]
port 215 nsew signal output
rlabel metal2 s 195058 0 195114 800 6 ext_data_rdata_o[16]
port 216 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 ext_data_rdata_o[17]
port 217 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 ext_data_rdata_o[18]
port 218 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 ext_data_rdata_o[19]
port 219 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 ext_data_rdata_o[1]
port 220 nsew signal output
rlabel metal2 s 197818 0 197874 800 6 ext_data_rdata_o[20]
port 221 nsew signal output
rlabel metal3 s 239066 127848 239866 127968 6 ext_data_rdata_o[21]
port 222 nsew signal output
rlabel metal2 s 151818 241210 151874 242010 6 ext_data_rdata_o[22]
port 223 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 ext_data_rdata_o[23]
port 224 nsew signal output
rlabel metal2 s 143538 241210 143594 242010 6 ext_data_rdata_o[24]
port 225 nsew signal output
rlabel metal2 s 193678 241210 193734 242010 6 ext_data_rdata_o[25]
port 226 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 ext_data_rdata_o[26]
port 227 nsew signal output
rlabel metal2 s 37738 241210 37794 242010 6 ext_data_rdata_o[27]
port 228 nsew signal output
rlabel metal2 s 218518 241210 218574 242010 6 ext_data_rdata_o[28]
port 229 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 ext_data_rdata_o[29]
port 230 nsew signal output
rlabel metal3 s 239066 82968 239866 83088 6 ext_data_rdata_o[2]
port 231 nsew signal output
rlabel metal2 s 138018 241210 138074 242010 6 ext_data_rdata_o[30]
port 232 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 ext_data_rdata_o[31]
port 233 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 ext_data_rdata_o[3]
port 234 nsew signal output
rlabel metal3 s 239066 131928 239866 132048 6 ext_data_rdata_o[4]
port 235 nsew signal output
rlabel metal2 s 12898 241210 12954 242010 6 ext_data_rdata_o[5]
port 236 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 ext_data_rdata_o[6]
port 237 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 ext_data_rdata_o[7]
port 238 nsew signal output
rlabel metal3 s 239066 53728 239866 53848 6 ext_data_rdata_o[8]
port 239 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 ext_data_rdata_o[9]
port 240 nsew signal output
rlabel metal2 s 173898 241210 173954 242010 6 ext_data_req_i
port 241 nsew signal input
rlabel metal2 s 207478 241210 207534 242010 6 ext_data_rvalid_i
port 242 nsew signal input
rlabel metal2 s 6918 241210 6974 242010 6 ext_data_wdata_i[0]
port 243 nsew signal input
rlabel metal2 s 123758 241210 123814 242010 6 ext_data_wdata_i[10]
port 244 nsew signal input
rlabel metal3 s 239066 152328 239866 152448 6 ext_data_wdata_i[11]
port 245 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 ext_data_wdata_i[12]
port 246 nsew signal input
rlabel metal2 s 212998 241210 213054 242010 6 ext_data_wdata_i[13]
port 247 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 ext_data_wdata_i[14]
port 248 nsew signal input
rlabel metal3 s 239066 99288 239866 99408 6 ext_data_wdata_i[15]
port 249 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 ext_data_wdata_i[16]
port 250 nsew signal input
rlabel metal2 s 149058 241210 149114 242010 6 ext_data_wdata_i[17]
port 251 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 ext_data_wdata_i[18]
port 252 nsew signal input
rlabel metal3 s 239066 144168 239866 144288 6 ext_data_wdata_i[19]
port 253 nsew signal input
rlabel metal3 s 239066 12928 239866 13048 6 ext_data_wdata_i[1]
port 254 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 ext_data_wdata_i[20]
port 255 nsew signal input
rlabel metal3 s 239066 210128 239866 210248 6 ext_data_wdata_i[21]
port 256 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 ext_data_wdata_i[22]
port 257 nsew signal input
rlabel metal3 s 239066 238688 239866 238808 6 ext_data_wdata_i[23]
port 258 nsew signal input
rlabel metal3 s 239066 45568 239866 45688 6 ext_data_wdata_i[24]
port 259 nsew signal input
rlabel metal2 s 235078 241210 235134 242010 6 ext_data_wdata_i[25]
port 260 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 ext_data_wdata_i[26]
port 261 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 ext_data_wdata_i[27]
port 262 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 ext_data_wdata_i[28]
port 263 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 ext_data_wdata_i[29]
port 264 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 ext_data_wdata_i[2]
port 265 nsew signal input
rlabel metal2 s 210238 241210 210294 242010 6 ext_data_wdata_i[30]
port 266 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 ext_data_wdata_i[31]
port 267 nsew signal input
rlabel metal2 s 120998 241210 121054 242010 6 ext_data_wdata_i[3]
port 268 nsew signal input
rlabel metal3 s 239066 41488 239866 41608 6 ext_data_wdata_i[4]
port 269 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 ext_data_wdata_i[5]
port 270 nsew signal input
rlabel metal3 s 239066 206048 239866 206168 6 ext_data_wdata_i[6]
port 271 nsew signal input
rlabel metal2 s 237838 241210 237894 242010 6 ext_data_wdata_i[7]
port 272 nsew signal input
rlabel metal3 s 239066 29248 239866 29368 6 ext_data_wdata_i[8]
port 273 nsew signal input
rlabel metal3 s 239066 197888 239866 198008 6 ext_data_wdata_i[9]
port 274 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 ext_data_we_i
port 275 nsew signal input
rlabel metal3 s 239066 4768 239866 4888 6 fetch_enable_i
port 276 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 irq_ack_o
port 277 nsew signal output
rlabel metal2 s 184018 0 184074 800 6 irq_i
port 278 nsew signal input
rlabel metal3 s 239066 189728 239866 189848 6 irq_id_i[0]
port 279 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 irq_id_i[1]
port 280 nsew signal input
rlabel metal2 s 112718 241210 112774 242010 6 irq_id_i[2]
port 281 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 irq_id_i[3]
port 282 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 irq_id_i[4]
port 283 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 irq_id_o[0]
port 284 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 irq_id_o[1]
port 285 nsew signal output
rlabel metal3 s 239066 95208 239866 95328 6 irq_id_o[2]
port 286 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 irq_id_o[3]
port 287 nsew signal output
rlabel metal3 s 0 185648 800 185768 6 irq_id_o[4]
port 288 nsew signal output
rlabel metal3 s 239066 214208 239866 214328 6 reset
port 289 nsew signal input
rlabel metal4 s 234208 2128 234528 239408 6 VPWR
port 290 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 239408 6 VPWR
port 291 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 239408 6 VPWR
port 292 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 239408 6 VPWR
port 293 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 239408 6 VPWR
port 294 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 239408 6 VPWR
port 295 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 239408 6 VPWR
port 296 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 239408 6 VPWR
port 297 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 239408 6 VPWR
port 298 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 239408 6 VPWR
port 299 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 239408 6 VPWR
port 300 nsew power bidirectional
rlabel metal4 s 124208 218452 124528 239408 6 VPWR
port 301 nsew power bidirectional
rlabel metal4 s 114208 218452 114528 239408 6 VPWR
port 302 nsew power bidirectional
rlabel metal4 s 104208 218452 104528 239408 6 VPWR
port 303 nsew power bidirectional
rlabel metal4 s 94208 218452 94528 239408 6 VPWR
port 304 nsew power bidirectional
rlabel metal4 s 84208 218452 84528 239408 6 VPWR
port 305 nsew power bidirectional
rlabel metal4 s 74208 218452 74528 239408 6 VPWR
port 306 nsew power bidirectional
rlabel metal4 s 64208 218452 64528 239408 6 VPWR
port 307 nsew power bidirectional
rlabel metal4 s 54208 218452 54528 239408 6 VPWR
port 308 nsew power bidirectional
rlabel metal4 s 44208 218452 44528 239408 6 VPWR
port 309 nsew power bidirectional
rlabel metal4 s 34208 218452 34528 239408 6 VPWR
port 310 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 239408 6 VPWR
port 311 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 239408 6 VPWR
port 312 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 239408 6 VPWR
port 313 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 137048 6 VPWR
port 314 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 137048 6 VPWR
port 315 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 137048 6 VPWR
port 316 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 137048 6 VPWR
port 317 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 137048 6 VPWR
port 318 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 137048 6 VPWR
port 319 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 137048 6 VPWR
port 320 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 137048 6 VPWR
port 321 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 137048 6 VPWR
port 322 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 137048 6 VPWR
port 323 nsew power bidirectional
rlabel metal5 s 1104 219750 238740 220070 6 VPWR
port 324 nsew power bidirectional
rlabel metal5 s 1104 189114 238740 189434 6 VPWR
port 325 nsew power bidirectional
rlabel metal5 s 1104 158478 238740 158798 6 VPWR
port 326 nsew power bidirectional
rlabel metal5 s 1104 127842 238740 128162 6 VPWR
port 327 nsew power bidirectional
rlabel metal5 s 1104 97206 238740 97526 6 VPWR
port 328 nsew power bidirectional
rlabel metal5 s 1104 66570 238740 66890 6 VPWR
port 329 nsew power bidirectional
rlabel metal5 s 1104 35934 238740 36254 6 VPWR
port 330 nsew power bidirectional
rlabel metal5 s 1104 5298 238740 5618 6 VPWR
port 331 nsew power bidirectional
rlabel metal4 s 229208 2128 229528 239408 6 VGND
port 332 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 239408 6 VGND
port 333 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 239408 6 VGND
port 334 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 239408 6 VGND
port 335 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 239408 6 VGND
port 336 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 239408 6 VGND
port 337 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 239408 6 VGND
port 338 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 239408 6 VGND
port 339 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 239408 6 VGND
port 340 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 239408 6 VGND
port 341 nsew ground bidirectional
rlabel metal4 s 129208 218452 129528 239408 6 VGND
port 342 nsew ground bidirectional
rlabel metal4 s 119208 218452 119528 239408 6 VGND
port 343 nsew ground bidirectional
rlabel metal4 s 109208 218452 109528 239408 6 VGND
port 344 nsew ground bidirectional
rlabel metal4 s 99208 218452 99528 239408 6 VGND
port 345 nsew ground bidirectional
rlabel metal4 s 89208 218452 89528 239408 6 VGND
port 346 nsew ground bidirectional
rlabel metal4 s 79208 218452 79528 239408 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 69208 218452 69528 239408 6 VGND
port 348 nsew ground bidirectional
rlabel metal4 s 59208 218452 59528 239408 6 VGND
port 349 nsew ground bidirectional
rlabel metal4 s 49208 218452 49528 239408 6 VGND
port 350 nsew ground bidirectional
rlabel metal4 s 39208 218452 39528 239408 6 VGND
port 351 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 239408 6 VGND
port 352 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 239408 6 VGND
port 353 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 239408 6 VGND
port 354 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 137048 6 VGND
port 355 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 137048 6 VGND
port 356 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 137048 6 VGND
port 357 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 137048 6 VGND
port 358 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 137048 6 VGND
port 359 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 137048 6 VGND
port 360 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 137048 6 VGND
port 361 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 137048 6 VGND
port 362 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 137048 6 VGND
port 363 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 137048 6 VGND
port 364 nsew ground bidirectional
rlabel metal5 s 1104 235068 238740 235388 6 VGND
port 365 nsew ground bidirectional
rlabel metal5 s 1104 204432 238740 204752 6 VGND
port 366 nsew ground bidirectional
rlabel metal5 s 1104 173796 238740 174116 6 VGND
port 367 nsew ground bidirectional
rlabel metal5 s 1104 143160 238740 143480 6 VGND
port 368 nsew ground bidirectional
rlabel metal5 s 1104 112524 238740 112844 6 VGND
port 369 nsew ground bidirectional
rlabel metal5 s 1104 81888 238740 82208 6 VGND
port 370 nsew ground bidirectional
rlabel metal5 s 1104 51252 238740 51572 6 VGND
port 371 nsew ground bidirectional
rlabel metal5 s 1104 20616 238740 20936 6 VGND
port 372 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 239866 242010
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 77608254
string GDS_START 10580018
<< end >>

