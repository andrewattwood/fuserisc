VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1197.990 BY 1208.710 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 1204.710 145.270 1208.710 ;
    END
  END clk_i
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 928.240 1197.990 928.840 ;
    END
  END debug_req_i
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 1204.710 1159.570 1208.710 ;
    END
  END eFPGA_delay_o[0]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 1204.710 853.670 1208.710 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 1204.710 437.370 1208.710 ;
    END
  END eFPGA_en_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 887.440 1197.990 888.040 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 333.240 1197.990 333.840 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1152.640 4.000 1153.240 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 1204.710 729.470 1208.710 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 1204.710 506.370 1208.710 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 537.240 1197.990 537.840 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 965.640 4.000 966.240 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 618.840 1197.990 619.440 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 1204.710 7.270 1208.710 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 1204.710 76.270 1208.710 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 805.840 1197.990 806.440 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 187.040 1197.990 187.640 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 700.440 1197.990 701.040 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 85.040 1197.990 85.640 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 1204.710 826.070 1208.710 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 1204.710 90.070 1208.710 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 1204.710 897.370 1208.710 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 1204.710 202.770 1208.710 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 1204.710 1104.370 1208.710 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 1204.710 464.970 1208.710 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 1204.710 784.670 1208.710 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 1204.710 550.070 1208.710 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 435.240 1197.990 435.840 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 1204.710 21.070 1208.710 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 802.440 4.000 803.040 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 0.000 711.070 4.000 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 0.000 1168.770 4.000 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 1204.710 980.170 1208.710 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 1204.710 423.570 1208.710 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 1204.710 478.770 1208.710 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 1204.710 1145.770 1208.710 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1173.040 1197.990 1173.640 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 1204.710 632.870 1208.710 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 907.840 1197.990 908.440 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 0.000 807.670 4.000 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 826.240 1197.990 826.840 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 1204.710 285.570 1208.710 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 0.000 515.570 4.000 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 353.640 1197.990 354.240 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 904.440 4.000 905.040 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 557.640 1197.990 558.240 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 1204.710 770.870 1208.710 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 1204.710 1021.570 1208.710 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 1204.710 103.870 1208.710 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 1204.710 172.870 1208.710 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1071.040 4.000 1071.640 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1091.440 1197.990 1092.040 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 312.840 1197.990 313.440 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 1204.710 911.170 1208.710 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 1204.710 271.770 1208.710 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 867.040 1197.990 867.640 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 1204.710 1007.770 1208.710 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 0.000 333.870 4.000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 105.440 1197.990 106.040 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 1204.710 326.970 1208.710 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 986.040 4.000 986.640 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 0.000 1154.970 4.000 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.390 1204.710 577.670 1208.710 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 1204.710 938.770 1208.710 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 0.000 931.870 4.000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1050.640 4.000 1051.240 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 680.040 1197.990 680.640 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 1204.710 1076.770 1208.710 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 1204.710 230.370 1208.710 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 166.640 1197.990 167.240 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.690 1204.710 993.970 1208.710 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 516.840 1197.990 517.440 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 1204.710 492.570 1208.710 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1152.640 1197.990 1153.240 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 1204.710 313.170 1208.710 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 125.840 1197.990 126.440 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 1204.710 451.170 1208.710 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1193.440 4.000 1194.040 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1111.840 1197.990 1112.440 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 0.000 1141.170 4.000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 0.000 1127.370 4.000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 1204.710 952.570 1208.710 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 578.040 1197.990 578.640 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 969.040 1197.990 969.640 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1009.840 1197.990 1010.440 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 1204.710 48.670 1208.710 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 44.240 1197.990 44.840 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 0.000 904.270 4.000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1132.240 4.000 1132.840 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 1204.710 660.470 1208.710 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 1204.710 883.570 1208.710 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 1204.710 340.770 1208.710 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 1204.710 812.270 1208.710 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 1204.710 839.870 1208.710 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 1204.710 701.870 1208.710 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 1204.710 117.670 1208.710 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.040 4.000 782.640 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 598.440 1197.990 599.040 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 744.640 1197.990 745.240 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 1204.710 1131.970 1208.710 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 0.000 612.170 4.000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 846.640 1197.990 847.240 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 1204.710 798.470 1208.710 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 1204.710 354.570 1208.710 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 1204.710 159.070 1208.710 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 394.440 1197.990 395.040 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 1204.710 257.970 1208.710 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.840 4.000 1010.440 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 455.640 1197.990 456.240 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 1204.710 368.370 1208.710 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END eFPGA_write_strobe_o
  PIN ext_data_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 1204.710 382.170 1208.710 ;
    END
  END ext_data_addr_i[0]
  PIN ext_data_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END ext_data_addr_i[10]
  PIN ext_data_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 3.440 1197.990 4.040 ;
    END
  END ext_data_addr_i[11]
  PIN ext_data_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 1204.710 395.970 1208.710 ;
    END
  END ext_data_addr_i[12]
  PIN ext_data_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 1204.710 591.470 1208.710 ;
    END
  END ext_data_addr_i[13]
  PIN ext_data_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.690 0.000 487.970 4.000 ;
    END
  END ext_data_addr_i[14]
  PIN ext_data_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END ext_data_addr_i[15]
  PIN ext_data_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 1204.710 536.270 1208.710 ;
    END
  END ext_data_addr_i[16]
  PIN ext_data_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 374.040 1197.990 374.640 ;
    END
  END ext_data_addr_i[17]
  PIN ext_data_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 785.440 1197.990 786.040 ;
    END
  END ext_data_addr_i[18]
  PIN ext_data_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END ext_data_addr_i[19]
  PIN ext_data_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 945.240 4.000 945.840 ;
    END
  END ext_data_addr_i[1]
  PIN ext_data_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END ext_data_addr_i[20]
  PIN ext_data_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END ext_data_addr_i[21]
  PIN ext_data_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END ext_data_addr_i[22]
  PIN ext_data_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 1204.710 646.670 1208.710 ;
    END
  END ext_data_addr_i[23]
  PIN ext_data_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 0.000 1113.570 4.000 ;
    END
  END ext_data_addr_i[24]
  PIN ext_data_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 251.640 1197.990 252.240 ;
    END
  END ext_data_addr_i[25]
  PIN ext_data_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 1204.710 1118.170 1208.710 ;
    END
  END ext_data_addr_i[26]
  PIN ext_data_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 0.000 1000.870 4.000 ;
    END
  END ext_data_addr_i[27]
  PIN ext_data_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 1204.710 244.170 1208.710 ;
    END
  END ext_data_addr_i[28]
  PIN ext_data_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 0.000 1182.570 4.000 ;
    END
  END ext_data_addr_i[29]
  PIN ext_data_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 1204.710 674.270 1208.710 ;
    END
  END ext_data_addr_i[2]
  PIN ext_data_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END ext_data_addr_i[30]
  PIN ext_data_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 1204.710 409.770 1208.710 ;
    END
  END ext_data_addr_i[31]
  PIN ext_data_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END ext_data_addr_i[3]
  PIN ext_data_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 1204.710 299.370 1208.710 ;
    END
  END ext_data_addr_i[4]
  PIN ext_data_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1091.440 4.000 1092.040 ;
    END
  END ext_data_addr_i[5]
  PIN ext_data_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 1204.710 924.970 1208.710 ;
    END
  END ext_data_addr_i[6]
  PIN ext_data_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 1204.710 216.570 1208.710 ;
    END
  END ext_data_addr_i[7]
  PIN ext_data_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END ext_data_addr_i[8]
  PIN ext_data_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1030.240 4.000 1030.840 ;
    END
  END ext_data_addr_i[9]
  PIN ext_data_be_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END ext_data_be_i[0]
  PIN ext_data_be_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 1204.710 131.470 1208.710 ;
    END
  END ext_data_be_i[1]
  PIN ext_data_be_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 0.000 1085.970 4.000 ;
    END
  END ext_data_be_i[2]
  PIN ext_data_be_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END ext_data_be_i[3]
  PIN ext_data_gnt_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 822.840 4.000 823.440 ;
    END
  END ext_data_gnt_o
  PIN ext_data_rdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1132.240 1197.990 1132.840 ;
    END
  END ext_data_rdata_o[0]
  PIN ext_data_rdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 0.000 959.470 4.000 ;
    END
  END ext_data_rdata_o[10]
  PIN ext_data_rdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END ext_data_rdata_o[11]
  PIN ext_data_rdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END ext_data_rdata_o[12]
  PIN ext_data_rdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 292.440 1197.990 293.040 ;
    END
  END ext_data_rdata_o[13]
  PIN ext_data_rdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 0.000 876.670 4.000 ;
    END
  END ext_data_rdata_o[14]
  PIN ext_data_rdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 1204.710 520.170 1208.710 ;
    END
  END ext_data_rdata_o[15]
  PIN ext_data_rdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 0.000 973.270 4.000 ;
    END
  END ext_data_rdata_o[16]
  PIN ext_data_rdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END ext_data_rdata_o[17]
  PIN ext_data_rdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END ext_data_rdata_o[18]
  PIN ext_data_rdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END ext_data_rdata_o[19]
  PIN ext_data_rdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END ext_data_rdata_o[1]
  PIN ext_data_rdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 0.000 987.070 4.000 ;
    END
  END ext_data_rdata_o[20]
  PIN ext_data_rdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 639.240 1197.990 639.840 ;
    END
  END ext_data_rdata_o[21]
  PIN ext_data_rdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 1204.710 757.070 1208.710 ;
    END
  END ext_data_rdata_o[22]
  PIN ext_data_rdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END ext_data_rdata_o[23]
  PIN ext_data_rdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 1204.710 715.670 1208.710 ;
    END
  END ext_data_rdata_o[24]
  PIN ext_data_rdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 1204.710 966.370 1208.710 ;
    END
  END ext_data_rdata_o[25]
  PIN ext_data_rdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.840 4.000 1112.440 ;
    END
  END ext_data_rdata_o[26]
  PIN ext_data_rdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 1204.710 186.670 1208.710 ;
    END
  END ext_data_rdata_o[27]
  PIN ext_data_rdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 1204.710 1090.570 1208.710 ;
    END
  END ext_data_rdata_o[28]
  PIN ext_data_rdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END ext_data_rdata_o[29]
  PIN ext_data_rdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 414.840 1197.990 415.440 ;
    END
  END ext_data_rdata_o[2]
  PIN ext_data_rdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 1204.710 688.070 1208.710 ;
    END
  END ext_data_rdata_o[30]
  PIN ext_data_rdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END ext_data_rdata_o[31]
  PIN ext_data_rdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END ext_data_rdata_o[3]
  PIN ext_data_rdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 659.640 1197.990 660.240 ;
    END
  END ext_data_rdata_o[4]
  PIN ext_data_rdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 1204.710 62.470 1208.710 ;
    END
  END ext_data_rdata_o[5]
  PIN ext_data_rdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END ext_data_rdata_o[6]
  PIN ext_data_rdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END ext_data_rdata_o[7]
  PIN ext_data_rdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 272.040 1197.990 272.640 ;
    END
  END ext_data_rdata_o[8]
  PIN ext_data_rdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END ext_data_rdata_o[9]
  PIN ext_data_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 1204.710 869.770 1208.710 ;
    END
  END ext_data_req_i
  PIN ext_data_rvalid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 1204.710 1035.370 1208.710 ;
    END
  END ext_data_rvalid_o
  PIN ext_data_wdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 1204.710 34.870 1208.710 ;
    END
  END ext_data_wdata_i[0]
  PIN ext_data_wdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 1204.710 619.070 1208.710 ;
    END
  END ext_data_wdata_i[10]
  PIN ext_data_wdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 765.040 1197.990 765.640 ;
    END
  END ext_data_wdata_i[11]
  PIN ext_data_wdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.490 0.000 501.770 4.000 ;
    END
  END ext_data_wdata_i[12]
  PIN ext_data_wdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 1204.710 1062.970 1208.710 ;
    END
  END ext_data_wdata_i[13]
  PIN ext_data_wdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 700.440 4.000 701.040 ;
    END
  END ext_data_wdata_i[14]
  PIN ext_data_wdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 496.440 1197.990 497.040 ;
    END
  END ext_data_wdata_i[15]
  PIN ext_data_wdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END ext_data_wdata_i[16]
  PIN ext_data_wdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 1204.710 743.270 1208.710 ;
    END
  END ext_data_wdata_i[17]
  PIN ext_data_wdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END ext_data_wdata_i[18]
  PIN ext_data_wdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 724.240 1197.990 724.840 ;
    END
  END ext_data_wdata_i[19]
  PIN ext_data_wdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 64.640 1197.990 65.240 ;
    END
  END ext_data_wdata_i[1]
  PIN ext_data_wdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.490 0.000 1099.770 4.000 ;
    END
  END ext_data_wdata_i[20]
  PIN ext_data_wdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1050.640 1197.990 1051.240 ;
    END
  END ext_data_wdata_i[21]
  PIN ext_data_wdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END ext_data_wdata_i[22]
  PIN ext_data_wdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1193.440 1197.990 1194.040 ;
    END
  END ext_data_wdata_i[23]
  PIN ext_data_wdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 231.240 1197.990 231.840 ;
    END
  END ext_data_wdata_i[24]
  PIN ext_data_wdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 1204.710 1173.370 1208.710 ;
    END
  END ext_data_wdata_i[25]
  PIN ext_data_wdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END ext_data_wdata_i[26]
  PIN ext_data_wdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END ext_data_wdata_i[27]
  PIN ext_data_wdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END ext_data_wdata_i[28]
  PIN ext_data_wdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END ext_data_wdata_i[29]
  PIN ext_data_wdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END ext_data_wdata_i[2]
  PIN ext_data_wdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 1204.710 1049.170 1208.710 ;
    END
  END ext_data_wdata_i[30]
  PIN ext_data_wdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END ext_data_wdata_i[31]
  PIN ext_data_wdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 1204.710 605.270 1208.710 ;
    END
  END ext_data_wdata_i[3]
  PIN ext_data_wdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 207.440 1197.990 208.040 ;
    END
  END ext_data_wdata_i[4]
  PIN ext_data_wdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END ext_data_wdata_i[5]
  PIN ext_data_wdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1030.240 1197.990 1030.840 ;
    END
  END ext_data_wdata_i[6]
  PIN ext_data_wdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 1204.710 1187.170 1208.710 ;
    END
  END ext_data_wdata_i[7]
  PIN ext_data_wdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 146.240 1197.990 146.840 ;
    END
  END ext_data_wdata_i[8]
  PIN ext_data_wdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 989.440 1197.990 990.040 ;
    END
  END ext_data_wdata_i[9]
  PIN ext_data_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END ext_data_we_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 23.840 1197.990 24.440 ;
    END
  END fetch_enable_i
  PIN irq_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END irq_ack_o
  PIN irq_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 0.000 918.070 4.000 ;
    END
  END irq_i
  PIN irq_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 948.640 1197.990 949.240 ;
    END
  END irq_id_i[0]
  PIN irq_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END irq_id_i[1]
  PIN irq_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 1204.710 563.870 1208.710 ;
    END
  END irq_id_i[2]
  PIN irq_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END irq_id_i[3]
  PIN irq_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END irq_id_i[4]
  PIN irq_id_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END irq_id_o[0]
  PIN irq_id_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END irq_id_o[1]
  PIN irq_id_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 476.040 1197.990 476.640 ;
    END
  END irq_id_o[2]
  PIN irq_id_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END irq_id_o[3]
  PIN irq_id_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 924.840 4.000 925.440 ;
    END
  END irq_id_o[4]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1193.990 1071.040 1197.990 1071.640 ;
    END
  END reset
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 1092.260 622.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 1092.260 572.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 1092.260 522.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 1092.260 472.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 1092.260 422.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 1092.260 372.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 1092.260 322.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 1092.260 272.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 1092.260 222.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 1092.260 172.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1197.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 685.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1098.750 1192.320 1100.350 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 945.570 1192.320 947.170 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 792.390 1192.320 793.990 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 1192.320 640.810 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 1192.320 487.630 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 1192.320 334.450 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 1192.320 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 1192.320 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 1092.260 647.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 1092.260 597.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 1092.260 547.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 1092.260 497.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 1092.260 447.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 1092.260 397.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 1092.260 347.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 1092.260 297.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 1092.260 247.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 1092.260 197.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 1197.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 685.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1175.340 1192.320 1176.940 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1022.160 1192.320 1023.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 868.980 1192.320 870.580 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 715.800 1192.320 717.400 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 1192.320 564.220 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 1192.320 411.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 1192.320 257.860 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 1192.320 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1192.320 1196.885 ;
      LAYER met1 ;
        RECT 2.370 7.860 1192.320 1197.440 ;
      LAYER met2 ;
        RECT 2.400 1204.430 6.710 1204.710 ;
        RECT 7.550 1204.430 20.510 1204.710 ;
        RECT 21.350 1204.430 34.310 1204.710 ;
        RECT 35.150 1204.430 48.110 1204.710 ;
        RECT 48.950 1204.430 61.910 1204.710 ;
        RECT 62.750 1204.430 75.710 1204.710 ;
        RECT 76.550 1204.430 89.510 1204.710 ;
        RECT 90.350 1204.430 103.310 1204.710 ;
        RECT 104.150 1204.430 117.110 1204.710 ;
        RECT 117.950 1204.430 130.910 1204.710 ;
        RECT 131.750 1204.430 144.710 1204.710 ;
        RECT 145.550 1204.430 158.510 1204.710 ;
        RECT 159.350 1204.430 172.310 1204.710 ;
        RECT 173.150 1204.430 186.110 1204.710 ;
        RECT 186.950 1204.430 202.210 1204.710 ;
        RECT 203.050 1204.430 216.010 1204.710 ;
        RECT 216.850 1204.430 229.810 1204.710 ;
        RECT 230.650 1204.430 243.610 1204.710 ;
        RECT 244.450 1204.430 257.410 1204.710 ;
        RECT 258.250 1204.430 271.210 1204.710 ;
        RECT 272.050 1204.430 285.010 1204.710 ;
        RECT 285.850 1204.430 298.810 1204.710 ;
        RECT 299.650 1204.430 312.610 1204.710 ;
        RECT 313.450 1204.430 326.410 1204.710 ;
        RECT 327.250 1204.430 340.210 1204.710 ;
        RECT 341.050 1204.430 354.010 1204.710 ;
        RECT 354.850 1204.430 367.810 1204.710 ;
        RECT 368.650 1204.430 381.610 1204.710 ;
        RECT 382.450 1204.430 395.410 1204.710 ;
        RECT 396.250 1204.430 409.210 1204.710 ;
        RECT 410.050 1204.430 423.010 1204.710 ;
        RECT 423.850 1204.430 436.810 1204.710 ;
        RECT 437.650 1204.430 450.610 1204.710 ;
        RECT 451.450 1204.430 464.410 1204.710 ;
        RECT 465.250 1204.430 478.210 1204.710 ;
        RECT 479.050 1204.430 492.010 1204.710 ;
        RECT 492.850 1204.430 505.810 1204.710 ;
        RECT 506.650 1204.430 519.610 1204.710 ;
        RECT 520.450 1204.430 535.710 1204.710 ;
        RECT 536.550 1204.430 549.510 1204.710 ;
        RECT 550.350 1204.430 563.310 1204.710 ;
        RECT 564.150 1204.430 577.110 1204.710 ;
        RECT 577.950 1204.430 590.910 1204.710 ;
        RECT 591.750 1204.430 604.710 1204.710 ;
        RECT 605.550 1204.430 618.510 1204.710 ;
        RECT 619.350 1204.430 632.310 1204.710 ;
        RECT 633.150 1204.430 646.110 1204.710 ;
        RECT 646.950 1204.430 659.910 1204.710 ;
        RECT 660.750 1204.430 673.710 1204.710 ;
        RECT 674.550 1204.430 687.510 1204.710 ;
        RECT 688.350 1204.430 701.310 1204.710 ;
        RECT 702.150 1204.430 715.110 1204.710 ;
        RECT 715.950 1204.430 728.910 1204.710 ;
        RECT 729.750 1204.430 742.710 1204.710 ;
        RECT 743.550 1204.430 756.510 1204.710 ;
        RECT 757.350 1204.430 770.310 1204.710 ;
        RECT 771.150 1204.430 784.110 1204.710 ;
        RECT 784.950 1204.430 797.910 1204.710 ;
        RECT 798.750 1204.430 811.710 1204.710 ;
        RECT 812.550 1204.430 825.510 1204.710 ;
        RECT 826.350 1204.430 839.310 1204.710 ;
        RECT 840.150 1204.430 853.110 1204.710 ;
        RECT 853.950 1204.430 869.210 1204.710 ;
        RECT 870.050 1204.430 883.010 1204.710 ;
        RECT 883.850 1204.430 896.810 1204.710 ;
        RECT 897.650 1204.430 910.610 1204.710 ;
        RECT 911.450 1204.430 924.410 1204.710 ;
        RECT 925.250 1204.430 938.210 1204.710 ;
        RECT 939.050 1204.430 952.010 1204.710 ;
        RECT 952.850 1204.430 965.810 1204.710 ;
        RECT 966.650 1204.430 979.610 1204.710 ;
        RECT 980.450 1204.430 993.410 1204.710 ;
        RECT 994.250 1204.430 1007.210 1204.710 ;
        RECT 1008.050 1204.430 1021.010 1204.710 ;
        RECT 1021.850 1204.430 1034.810 1204.710 ;
        RECT 1035.650 1204.430 1048.610 1204.710 ;
        RECT 1049.450 1204.430 1062.410 1204.710 ;
        RECT 1063.250 1204.430 1076.210 1204.710 ;
        RECT 1077.050 1204.430 1090.010 1204.710 ;
        RECT 1090.850 1204.430 1103.810 1204.710 ;
        RECT 1104.650 1204.430 1117.610 1204.710 ;
        RECT 1118.450 1204.430 1131.410 1204.710 ;
        RECT 1132.250 1204.430 1145.210 1204.710 ;
        RECT 1146.050 1204.430 1159.010 1204.710 ;
        RECT 1159.850 1204.430 1172.810 1204.710 ;
        RECT 1173.650 1204.430 1186.610 1204.710 ;
        RECT 1187.450 1204.430 1190.390 1204.710 ;
        RECT 2.400 4.280 1190.390 1204.430 ;
        RECT 2.950 3.555 15.910 4.280 ;
        RECT 16.750 3.555 29.710 4.280 ;
        RECT 30.550 3.555 43.510 4.280 ;
        RECT 44.350 3.555 57.310 4.280 ;
        RECT 58.150 3.555 71.110 4.280 ;
        RECT 71.950 3.555 84.910 4.280 ;
        RECT 85.750 3.555 98.710 4.280 ;
        RECT 99.550 3.555 112.510 4.280 ;
        RECT 113.350 3.555 126.310 4.280 ;
        RECT 127.150 3.555 140.110 4.280 ;
        RECT 140.950 3.555 153.910 4.280 ;
        RECT 154.750 3.555 167.710 4.280 ;
        RECT 168.550 3.555 181.510 4.280 ;
        RECT 182.350 3.555 195.310 4.280 ;
        RECT 196.150 3.555 209.110 4.280 ;
        RECT 209.950 3.555 222.910 4.280 ;
        RECT 223.750 3.555 236.710 4.280 ;
        RECT 237.550 3.555 250.510 4.280 ;
        RECT 251.350 3.555 264.310 4.280 ;
        RECT 265.150 3.555 278.110 4.280 ;
        RECT 278.950 3.555 291.910 4.280 ;
        RECT 292.750 3.555 305.710 4.280 ;
        RECT 306.550 3.555 319.510 4.280 ;
        RECT 320.350 3.555 333.310 4.280 ;
        RECT 334.150 3.555 349.410 4.280 ;
        RECT 350.250 3.555 363.210 4.280 ;
        RECT 364.050 3.555 377.010 4.280 ;
        RECT 377.850 3.555 390.810 4.280 ;
        RECT 391.650 3.555 404.610 4.280 ;
        RECT 405.450 3.555 418.410 4.280 ;
        RECT 419.250 3.555 432.210 4.280 ;
        RECT 433.050 3.555 446.010 4.280 ;
        RECT 446.850 3.555 459.810 4.280 ;
        RECT 460.650 3.555 473.610 4.280 ;
        RECT 474.450 3.555 487.410 4.280 ;
        RECT 488.250 3.555 501.210 4.280 ;
        RECT 502.050 3.555 515.010 4.280 ;
        RECT 515.850 3.555 528.810 4.280 ;
        RECT 529.650 3.555 542.610 4.280 ;
        RECT 543.450 3.555 556.410 4.280 ;
        RECT 557.250 3.555 570.210 4.280 ;
        RECT 571.050 3.555 584.010 4.280 ;
        RECT 584.850 3.555 597.810 4.280 ;
        RECT 598.650 3.555 611.610 4.280 ;
        RECT 612.450 3.555 625.410 4.280 ;
        RECT 626.250 3.555 639.210 4.280 ;
        RECT 640.050 3.555 653.010 4.280 ;
        RECT 653.850 3.555 666.810 4.280 ;
        RECT 667.650 3.555 682.910 4.280 ;
        RECT 683.750 3.555 696.710 4.280 ;
        RECT 697.550 3.555 710.510 4.280 ;
        RECT 711.350 3.555 724.310 4.280 ;
        RECT 725.150 3.555 738.110 4.280 ;
        RECT 738.950 3.555 751.910 4.280 ;
        RECT 752.750 3.555 765.710 4.280 ;
        RECT 766.550 3.555 779.510 4.280 ;
        RECT 780.350 3.555 793.310 4.280 ;
        RECT 794.150 3.555 807.110 4.280 ;
        RECT 807.950 3.555 820.910 4.280 ;
        RECT 821.750 3.555 834.710 4.280 ;
        RECT 835.550 3.555 848.510 4.280 ;
        RECT 849.350 3.555 862.310 4.280 ;
        RECT 863.150 3.555 876.110 4.280 ;
        RECT 876.950 3.555 889.910 4.280 ;
        RECT 890.750 3.555 903.710 4.280 ;
        RECT 904.550 3.555 917.510 4.280 ;
        RECT 918.350 3.555 931.310 4.280 ;
        RECT 932.150 3.555 945.110 4.280 ;
        RECT 945.950 3.555 958.910 4.280 ;
        RECT 959.750 3.555 972.710 4.280 ;
        RECT 973.550 3.555 986.510 4.280 ;
        RECT 987.350 3.555 1000.310 4.280 ;
        RECT 1001.150 3.555 1016.410 4.280 ;
        RECT 1017.250 3.555 1030.210 4.280 ;
        RECT 1031.050 3.555 1044.010 4.280 ;
        RECT 1044.850 3.555 1057.810 4.280 ;
        RECT 1058.650 3.555 1071.610 4.280 ;
        RECT 1072.450 3.555 1085.410 4.280 ;
        RECT 1086.250 3.555 1099.210 4.280 ;
        RECT 1100.050 3.555 1113.010 4.280 ;
        RECT 1113.850 3.555 1126.810 4.280 ;
        RECT 1127.650 3.555 1140.610 4.280 ;
        RECT 1141.450 3.555 1154.410 4.280 ;
        RECT 1155.250 3.555 1168.210 4.280 ;
        RECT 1169.050 3.555 1182.010 4.280 ;
        RECT 1182.850 3.555 1190.390 4.280 ;
      LAYER met3 ;
        RECT 4.000 1194.440 1193.990 1197.985 ;
        RECT 4.400 1193.040 1193.590 1194.440 ;
        RECT 4.000 1174.040 1193.990 1193.040 ;
        RECT 4.400 1172.640 1193.590 1174.040 ;
        RECT 4.000 1153.640 1193.990 1172.640 ;
        RECT 4.400 1152.240 1193.590 1153.640 ;
        RECT 4.000 1133.240 1193.990 1152.240 ;
        RECT 4.400 1131.840 1193.590 1133.240 ;
        RECT 4.000 1112.840 1193.990 1131.840 ;
        RECT 4.400 1111.440 1193.590 1112.840 ;
        RECT 4.000 1092.440 1193.990 1111.440 ;
        RECT 4.400 1091.040 1193.590 1092.440 ;
        RECT 4.000 1072.040 1193.990 1091.040 ;
        RECT 4.400 1070.640 1193.590 1072.040 ;
        RECT 4.000 1051.640 1193.990 1070.640 ;
        RECT 4.400 1050.240 1193.590 1051.640 ;
        RECT 4.000 1031.240 1193.990 1050.240 ;
        RECT 4.400 1029.840 1193.590 1031.240 ;
        RECT 4.000 1010.840 1193.990 1029.840 ;
        RECT 4.400 1009.440 1193.590 1010.840 ;
        RECT 4.000 990.440 1193.990 1009.440 ;
        RECT 4.000 989.040 1193.590 990.440 ;
        RECT 4.000 987.040 1193.990 989.040 ;
        RECT 4.400 985.640 1193.990 987.040 ;
        RECT 4.000 970.040 1193.990 985.640 ;
        RECT 4.000 968.640 1193.590 970.040 ;
        RECT 4.000 966.640 1193.990 968.640 ;
        RECT 4.400 965.240 1193.990 966.640 ;
        RECT 4.000 949.640 1193.990 965.240 ;
        RECT 4.000 948.240 1193.590 949.640 ;
        RECT 4.000 946.240 1193.990 948.240 ;
        RECT 4.400 944.840 1193.990 946.240 ;
        RECT 4.000 929.240 1193.990 944.840 ;
        RECT 4.000 927.840 1193.590 929.240 ;
        RECT 4.000 925.840 1193.990 927.840 ;
        RECT 4.400 924.440 1193.990 925.840 ;
        RECT 4.000 908.840 1193.990 924.440 ;
        RECT 4.000 907.440 1193.590 908.840 ;
        RECT 4.000 905.440 1193.990 907.440 ;
        RECT 4.400 904.040 1193.990 905.440 ;
        RECT 4.000 888.440 1193.990 904.040 ;
        RECT 4.000 887.040 1193.590 888.440 ;
        RECT 4.000 885.040 1193.990 887.040 ;
        RECT 4.400 883.640 1193.990 885.040 ;
        RECT 4.000 868.040 1193.990 883.640 ;
        RECT 4.000 866.640 1193.590 868.040 ;
        RECT 4.000 864.640 1193.990 866.640 ;
        RECT 4.400 863.240 1193.990 864.640 ;
        RECT 4.000 847.640 1193.990 863.240 ;
        RECT 4.000 846.240 1193.590 847.640 ;
        RECT 4.000 844.240 1193.990 846.240 ;
        RECT 4.400 842.840 1193.990 844.240 ;
        RECT 4.000 827.240 1193.990 842.840 ;
        RECT 4.000 825.840 1193.590 827.240 ;
        RECT 4.000 823.840 1193.990 825.840 ;
        RECT 4.400 822.440 1193.990 823.840 ;
        RECT 4.000 806.840 1193.990 822.440 ;
        RECT 4.000 805.440 1193.590 806.840 ;
        RECT 4.000 803.440 1193.990 805.440 ;
        RECT 4.400 802.040 1193.990 803.440 ;
        RECT 4.000 786.440 1193.990 802.040 ;
        RECT 4.000 785.040 1193.590 786.440 ;
        RECT 4.000 783.040 1193.990 785.040 ;
        RECT 4.400 781.640 1193.990 783.040 ;
        RECT 4.000 766.040 1193.990 781.640 ;
        RECT 4.000 764.640 1193.590 766.040 ;
        RECT 4.000 762.640 1193.990 764.640 ;
        RECT 4.400 761.240 1193.990 762.640 ;
        RECT 4.000 745.640 1193.990 761.240 ;
        RECT 4.000 744.240 1193.590 745.640 ;
        RECT 4.000 742.240 1193.990 744.240 ;
        RECT 4.400 740.840 1193.990 742.240 ;
        RECT 4.000 725.240 1193.990 740.840 ;
        RECT 4.000 723.840 1193.590 725.240 ;
        RECT 4.000 721.840 1193.990 723.840 ;
        RECT 4.400 720.440 1193.990 721.840 ;
        RECT 4.000 701.440 1193.990 720.440 ;
        RECT 4.400 700.040 1193.590 701.440 ;
        RECT 4.000 681.040 1193.990 700.040 ;
        RECT 4.400 679.640 1193.590 681.040 ;
        RECT 4.000 660.640 1193.990 679.640 ;
        RECT 4.400 659.240 1193.590 660.640 ;
        RECT 4.000 640.240 1193.990 659.240 ;
        RECT 4.400 638.840 1193.590 640.240 ;
        RECT 4.000 619.840 1193.990 638.840 ;
        RECT 4.400 618.440 1193.590 619.840 ;
        RECT 4.000 599.440 1193.990 618.440 ;
        RECT 4.400 598.040 1193.590 599.440 ;
        RECT 4.000 579.040 1193.990 598.040 ;
        RECT 4.400 577.640 1193.590 579.040 ;
        RECT 4.000 558.640 1193.990 577.640 ;
        RECT 4.400 557.240 1193.590 558.640 ;
        RECT 4.000 538.240 1193.990 557.240 ;
        RECT 4.400 536.840 1193.590 538.240 ;
        RECT 4.000 517.840 1193.990 536.840 ;
        RECT 4.400 516.440 1193.590 517.840 ;
        RECT 4.000 497.440 1193.990 516.440 ;
        RECT 4.000 496.040 1193.590 497.440 ;
        RECT 4.000 494.040 1193.990 496.040 ;
        RECT 4.400 492.640 1193.990 494.040 ;
        RECT 4.000 477.040 1193.990 492.640 ;
        RECT 4.000 475.640 1193.590 477.040 ;
        RECT 4.000 473.640 1193.990 475.640 ;
        RECT 4.400 472.240 1193.990 473.640 ;
        RECT 4.000 456.640 1193.990 472.240 ;
        RECT 4.000 455.240 1193.590 456.640 ;
        RECT 4.000 453.240 1193.990 455.240 ;
        RECT 4.400 451.840 1193.990 453.240 ;
        RECT 4.000 436.240 1193.990 451.840 ;
        RECT 4.000 434.840 1193.590 436.240 ;
        RECT 4.000 432.840 1193.990 434.840 ;
        RECT 4.400 431.440 1193.990 432.840 ;
        RECT 4.000 415.840 1193.990 431.440 ;
        RECT 4.000 414.440 1193.590 415.840 ;
        RECT 4.000 412.440 1193.990 414.440 ;
        RECT 4.400 411.040 1193.990 412.440 ;
        RECT 4.000 395.440 1193.990 411.040 ;
        RECT 4.000 394.040 1193.590 395.440 ;
        RECT 4.000 392.040 1193.990 394.040 ;
        RECT 4.400 390.640 1193.990 392.040 ;
        RECT 4.000 375.040 1193.990 390.640 ;
        RECT 4.000 373.640 1193.590 375.040 ;
        RECT 4.000 371.640 1193.990 373.640 ;
        RECT 4.400 370.240 1193.990 371.640 ;
        RECT 4.000 354.640 1193.990 370.240 ;
        RECT 4.000 353.240 1193.590 354.640 ;
        RECT 4.000 351.240 1193.990 353.240 ;
        RECT 4.400 349.840 1193.990 351.240 ;
        RECT 4.000 334.240 1193.990 349.840 ;
        RECT 4.000 332.840 1193.590 334.240 ;
        RECT 4.000 330.840 1193.990 332.840 ;
        RECT 4.400 329.440 1193.990 330.840 ;
        RECT 4.000 313.840 1193.990 329.440 ;
        RECT 4.000 312.440 1193.590 313.840 ;
        RECT 4.000 310.440 1193.990 312.440 ;
        RECT 4.400 309.040 1193.990 310.440 ;
        RECT 4.000 293.440 1193.990 309.040 ;
        RECT 4.000 292.040 1193.590 293.440 ;
        RECT 4.000 290.040 1193.990 292.040 ;
        RECT 4.400 288.640 1193.990 290.040 ;
        RECT 4.000 273.040 1193.990 288.640 ;
        RECT 4.000 271.640 1193.590 273.040 ;
        RECT 4.000 269.640 1193.990 271.640 ;
        RECT 4.400 268.240 1193.990 269.640 ;
        RECT 4.000 252.640 1193.990 268.240 ;
        RECT 4.000 251.240 1193.590 252.640 ;
        RECT 4.000 249.240 1193.990 251.240 ;
        RECT 4.400 247.840 1193.990 249.240 ;
        RECT 4.000 232.240 1193.990 247.840 ;
        RECT 4.000 230.840 1193.590 232.240 ;
        RECT 4.000 228.840 1193.990 230.840 ;
        RECT 4.400 227.440 1193.990 228.840 ;
        RECT 4.000 208.440 1193.990 227.440 ;
        RECT 4.400 207.040 1193.590 208.440 ;
        RECT 4.000 188.040 1193.990 207.040 ;
        RECT 4.400 186.640 1193.590 188.040 ;
        RECT 4.000 167.640 1193.990 186.640 ;
        RECT 4.400 166.240 1193.590 167.640 ;
        RECT 4.000 147.240 1193.990 166.240 ;
        RECT 4.400 145.840 1193.590 147.240 ;
        RECT 4.000 126.840 1193.990 145.840 ;
        RECT 4.400 125.440 1193.590 126.840 ;
        RECT 4.000 106.440 1193.990 125.440 ;
        RECT 4.400 105.040 1193.590 106.440 ;
        RECT 4.000 86.040 1193.990 105.040 ;
        RECT 4.400 84.640 1193.590 86.040 ;
        RECT 4.000 65.640 1193.990 84.640 ;
        RECT 4.400 64.240 1193.590 65.640 ;
        RECT 4.000 45.240 1193.990 64.240 ;
        RECT 4.400 43.840 1193.590 45.240 ;
        RECT 4.000 24.840 1193.990 43.840 ;
        RECT 4.400 23.440 1193.590 24.840 ;
        RECT 4.000 4.440 1193.990 23.440 ;
        RECT 4.000 3.575 1193.590 4.440 ;
      LAYER met4 ;
        RECT 159.455 1197.440 869.105 1197.985 ;
        RECT 159.455 1091.860 170.640 1197.440 ;
        RECT 173.040 1091.860 195.640 1197.440 ;
        RECT 198.040 1091.860 220.640 1197.440 ;
        RECT 223.040 1091.860 245.640 1197.440 ;
        RECT 248.040 1091.860 270.640 1197.440 ;
        RECT 273.040 1091.860 295.640 1197.440 ;
        RECT 298.040 1091.860 320.640 1197.440 ;
        RECT 323.040 1091.860 345.640 1197.440 ;
        RECT 348.040 1091.860 370.640 1197.440 ;
        RECT 373.040 1091.860 395.640 1197.440 ;
        RECT 398.040 1091.860 420.640 1197.440 ;
        RECT 423.040 1091.860 445.640 1197.440 ;
        RECT 448.040 1091.860 470.640 1197.440 ;
        RECT 473.040 1091.860 495.640 1197.440 ;
        RECT 498.040 1091.860 520.640 1197.440 ;
        RECT 523.040 1091.860 545.640 1197.440 ;
        RECT 548.040 1091.860 570.640 1197.440 ;
        RECT 573.040 1091.860 595.640 1197.440 ;
        RECT 598.040 1091.860 620.640 1197.440 ;
        RECT 623.040 1091.860 645.640 1197.440 ;
        RECT 648.040 1091.860 670.640 1197.440 ;
        RECT 159.455 685.640 670.640 1091.860 ;
        RECT 159.455 10.240 170.640 685.640 ;
        RECT 173.040 10.240 195.640 685.640 ;
        RECT 198.040 10.240 220.640 685.640 ;
        RECT 223.040 10.240 245.640 685.640 ;
        RECT 248.040 10.240 270.640 685.640 ;
        RECT 273.040 10.240 295.640 685.640 ;
        RECT 298.040 10.240 320.640 685.640 ;
        RECT 323.040 10.240 345.640 685.640 ;
        RECT 348.040 10.240 370.640 685.640 ;
        RECT 373.040 10.240 395.640 685.640 ;
        RECT 398.040 10.240 420.640 685.640 ;
        RECT 423.040 10.240 445.640 685.640 ;
        RECT 448.040 10.240 470.640 685.640 ;
        RECT 473.040 10.240 495.640 685.640 ;
        RECT 498.040 10.240 520.640 685.640 ;
        RECT 523.040 10.240 545.640 685.640 ;
        RECT 548.040 10.240 570.640 685.640 ;
        RECT 573.040 10.240 595.640 685.640 ;
        RECT 598.040 10.240 620.640 685.640 ;
        RECT 623.040 10.240 645.640 685.640 ;
        RECT 648.040 10.240 670.640 685.640 ;
        RECT 673.040 10.240 695.640 1197.440 ;
        RECT 698.040 10.240 720.640 1197.440 ;
        RECT 723.040 10.240 745.640 1197.440 ;
        RECT 748.040 10.240 770.640 1197.440 ;
        RECT 773.040 10.240 795.640 1197.440 ;
        RECT 798.040 10.240 820.640 1197.440 ;
        RECT 823.040 10.240 845.640 1197.440 ;
        RECT 848.040 10.240 869.105 1197.440 ;
        RECT 159.455 9.015 869.105 10.240 ;
  END
END user_proj_example
END LIBRARY

