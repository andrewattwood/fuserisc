magic
tech sky130A
magscale 1 2
timestamp 1624298571
<< obsli1 >>
rect 1104 2159 238464 239377
<< obsm1 >>
rect 474 1572 238464 239488
<< metal2 >>
rect 1398 240942 1454 241742
rect 4158 240942 4214 241742
rect 6918 240942 6974 241742
rect 9678 240942 9734 241742
rect 12438 240942 12494 241742
rect 15198 240942 15254 241742
rect 17958 240942 18014 241742
rect 20718 240942 20774 241742
rect 23478 240942 23534 241742
rect 26238 240942 26294 241742
rect 28998 240942 29054 241742
rect 31758 240942 31814 241742
rect 34518 240942 34574 241742
rect 37278 240942 37334 241742
rect 40498 240942 40554 241742
rect 43258 240942 43314 241742
rect 46018 240942 46074 241742
rect 48778 240942 48834 241742
rect 51538 240942 51594 241742
rect 54298 240942 54354 241742
rect 57058 240942 57114 241742
rect 59818 240942 59874 241742
rect 62578 240942 62634 241742
rect 65338 240942 65394 241742
rect 68098 240942 68154 241742
rect 70858 240942 70914 241742
rect 73618 240942 73674 241742
rect 76378 240942 76434 241742
rect 79138 240942 79194 241742
rect 81898 240942 81954 241742
rect 84658 240942 84714 241742
rect 87418 240942 87474 241742
rect 90178 240942 90234 241742
rect 92938 240942 92994 241742
rect 95698 240942 95754 241742
rect 98458 240942 98514 241742
rect 101218 240942 101274 241742
rect 103978 240942 104034 241742
rect 107198 240942 107254 241742
rect 109958 240942 110014 241742
rect 112718 240942 112774 241742
rect 115478 240942 115534 241742
rect 118238 240942 118294 241742
rect 120998 240942 121054 241742
rect 123758 240942 123814 241742
rect 126518 240942 126574 241742
rect 129278 240942 129334 241742
rect 132038 240942 132094 241742
rect 134798 240942 134854 241742
rect 137558 240942 137614 241742
rect 140318 240942 140374 241742
rect 143078 240942 143134 241742
rect 145838 240942 145894 241742
rect 148598 240942 148654 241742
rect 151358 240942 151414 241742
rect 154118 240942 154174 241742
rect 156878 240942 156934 241742
rect 159638 240942 159694 241742
rect 162398 240942 162454 241742
rect 165158 240942 165214 241742
rect 167918 240942 167974 241742
rect 170678 240942 170734 241742
rect 173898 240942 173954 241742
rect 176658 240942 176714 241742
rect 179418 240942 179474 241742
rect 182178 240942 182234 241742
rect 184938 240942 184994 241742
rect 187698 240942 187754 241742
rect 190458 240942 190514 241742
rect 193218 240942 193274 241742
rect 195978 240942 196034 241742
rect 198738 240942 198794 241742
rect 201498 240942 201554 241742
rect 204258 240942 204314 241742
rect 207018 240942 207074 241742
rect 209778 240942 209834 241742
rect 212538 240942 212594 241742
rect 215298 240942 215354 241742
rect 218058 240942 218114 241742
rect 220818 240942 220874 241742
rect 223578 240942 223634 241742
rect 226338 240942 226394 241742
rect 229098 240942 229154 241742
rect 231858 240942 231914 241742
rect 234618 240942 234674 241742
rect 237378 240942 237434 241742
rect 478 0 534 800
rect 3238 0 3294 800
rect 5998 0 6054 800
rect 8758 0 8814 800
rect 11518 0 11574 800
rect 14278 0 14334 800
rect 17038 0 17094 800
rect 19798 0 19854 800
rect 22558 0 22614 800
rect 25318 0 25374 800
rect 28078 0 28134 800
rect 30838 0 30894 800
rect 33598 0 33654 800
rect 36358 0 36414 800
rect 39118 0 39174 800
rect 41878 0 41934 800
rect 44638 0 44694 800
rect 47398 0 47454 800
rect 50158 0 50214 800
rect 52918 0 52974 800
rect 55678 0 55734 800
rect 58438 0 58494 800
rect 61198 0 61254 800
rect 63958 0 64014 800
rect 66718 0 66774 800
rect 69938 0 69994 800
rect 72698 0 72754 800
rect 75458 0 75514 800
rect 78218 0 78274 800
rect 80978 0 81034 800
rect 83738 0 83794 800
rect 86498 0 86554 800
rect 89258 0 89314 800
rect 92018 0 92074 800
rect 94778 0 94834 800
rect 97538 0 97594 800
rect 100298 0 100354 800
rect 103058 0 103114 800
rect 105818 0 105874 800
rect 108578 0 108634 800
rect 111338 0 111394 800
rect 114098 0 114154 800
rect 116858 0 116914 800
rect 119618 0 119674 800
rect 122378 0 122434 800
rect 125138 0 125194 800
rect 127898 0 127954 800
rect 130658 0 130714 800
rect 133418 0 133474 800
rect 136638 0 136694 800
rect 139398 0 139454 800
rect 142158 0 142214 800
rect 144918 0 144974 800
rect 147678 0 147734 800
rect 150438 0 150494 800
rect 153198 0 153254 800
rect 155958 0 156014 800
rect 158718 0 158774 800
rect 161478 0 161534 800
rect 164238 0 164294 800
rect 166998 0 167054 800
rect 169758 0 169814 800
rect 172518 0 172574 800
rect 175278 0 175334 800
rect 178038 0 178094 800
rect 180798 0 180854 800
rect 183558 0 183614 800
rect 186318 0 186374 800
rect 189078 0 189134 800
rect 191838 0 191894 800
rect 194598 0 194654 800
rect 197358 0 197414 800
rect 200118 0 200174 800
rect 203338 0 203394 800
rect 206098 0 206154 800
rect 208858 0 208914 800
rect 211618 0 211674 800
rect 214378 0 214434 800
rect 217138 0 217194 800
rect 219898 0 219954 800
rect 222658 0 222714 800
rect 225418 0 225474 800
rect 228178 0 228234 800
rect 230938 0 230994 800
rect 233698 0 233754 800
rect 236458 0 236514 800
<< obsm2 >>
rect 480 240886 1342 240942
rect 1510 240886 4102 240942
rect 4270 240886 6862 240942
rect 7030 240886 9622 240942
rect 9790 240886 12382 240942
rect 12550 240886 15142 240942
rect 15310 240886 17902 240942
rect 18070 240886 20662 240942
rect 20830 240886 23422 240942
rect 23590 240886 26182 240942
rect 26350 240886 28942 240942
rect 29110 240886 31702 240942
rect 31870 240886 34462 240942
rect 34630 240886 37222 240942
rect 37390 240886 40442 240942
rect 40610 240886 43202 240942
rect 43370 240886 45962 240942
rect 46130 240886 48722 240942
rect 48890 240886 51482 240942
rect 51650 240886 54242 240942
rect 54410 240886 57002 240942
rect 57170 240886 59762 240942
rect 59930 240886 62522 240942
rect 62690 240886 65282 240942
rect 65450 240886 68042 240942
rect 68210 240886 70802 240942
rect 70970 240886 73562 240942
rect 73730 240886 76322 240942
rect 76490 240886 79082 240942
rect 79250 240886 81842 240942
rect 82010 240886 84602 240942
rect 84770 240886 87362 240942
rect 87530 240886 90122 240942
rect 90290 240886 92882 240942
rect 93050 240886 95642 240942
rect 95810 240886 98402 240942
rect 98570 240886 101162 240942
rect 101330 240886 103922 240942
rect 104090 240886 107142 240942
rect 107310 240886 109902 240942
rect 110070 240886 112662 240942
rect 112830 240886 115422 240942
rect 115590 240886 118182 240942
rect 118350 240886 120942 240942
rect 121110 240886 123702 240942
rect 123870 240886 126462 240942
rect 126630 240886 129222 240942
rect 129390 240886 131982 240942
rect 132150 240886 134742 240942
rect 134910 240886 137502 240942
rect 137670 240886 140262 240942
rect 140430 240886 143022 240942
rect 143190 240886 145782 240942
rect 145950 240886 148542 240942
rect 148710 240886 151302 240942
rect 151470 240886 154062 240942
rect 154230 240886 156822 240942
rect 156990 240886 159582 240942
rect 159750 240886 162342 240942
rect 162510 240886 165102 240942
rect 165270 240886 167862 240942
rect 168030 240886 170622 240942
rect 170790 240886 173842 240942
rect 174010 240886 176602 240942
rect 176770 240886 179362 240942
rect 179530 240886 182122 240942
rect 182290 240886 184882 240942
rect 185050 240886 187642 240942
rect 187810 240886 190402 240942
rect 190570 240886 193162 240942
rect 193330 240886 195922 240942
rect 196090 240886 198682 240942
rect 198850 240886 201442 240942
rect 201610 240886 204202 240942
rect 204370 240886 206962 240942
rect 207130 240886 209722 240942
rect 209890 240886 212482 240942
rect 212650 240886 215242 240942
rect 215410 240886 218002 240942
rect 218170 240886 220762 240942
rect 220930 240886 223522 240942
rect 223690 240886 226282 240942
rect 226450 240886 229042 240942
rect 229210 240886 231802 240942
rect 231970 240886 234562 240942
rect 234730 240886 237322 240942
rect 237490 240886 238078 240942
rect 480 856 238078 240886
rect 590 711 3182 856
rect 3350 711 5942 856
rect 6110 711 8702 856
rect 8870 711 11462 856
rect 11630 711 14222 856
rect 14390 711 16982 856
rect 17150 711 19742 856
rect 19910 711 22502 856
rect 22670 711 25262 856
rect 25430 711 28022 856
rect 28190 711 30782 856
rect 30950 711 33542 856
rect 33710 711 36302 856
rect 36470 711 39062 856
rect 39230 711 41822 856
rect 41990 711 44582 856
rect 44750 711 47342 856
rect 47510 711 50102 856
rect 50270 711 52862 856
rect 53030 711 55622 856
rect 55790 711 58382 856
rect 58550 711 61142 856
rect 61310 711 63902 856
rect 64070 711 66662 856
rect 66830 711 69882 856
rect 70050 711 72642 856
rect 72810 711 75402 856
rect 75570 711 78162 856
rect 78330 711 80922 856
rect 81090 711 83682 856
rect 83850 711 86442 856
rect 86610 711 89202 856
rect 89370 711 91962 856
rect 92130 711 94722 856
rect 94890 711 97482 856
rect 97650 711 100242 856
rect 100410 711 103002 856
rect 103170 711 105762 856
rect 105930 711 108522 856
rect 108690 711 111282 856
rect 111450 711 114042 856
rect 114210 711 116802 856
rect 116970 711 119562 856
rect 119730 711 122322 856
rect 122490 711 125082 856
rect 125250 711 127842 856
rect 128010 711 130602 856
rect 130770 711 133362 856
rect 133530 711 136582 856
rect 136750 711 139342 856
rect 139510 711 142102 856
rect 142270 711 144862 856
rect 145030 711 147622 856
rect 147790 711 150382 856
rect 150550 711 153142 856
rect 153310 711 155902 856
rect 156070 711 158662 856
rect 158830 711 161422 856
rect 161590 711 164182 856
rect 164350 711 166942 856
rect 167110 711 169702 856
rect 169870 711 172462 856
rect 172630 711 175222 856
rect 175390 711 177982 856
rect 178150 711 180742 856
rect 180910 711 183502 856
rect 183670 711 186262 856
rect 186430 711 189022 856
rect 189190 711 191782 856
rect 191950 711 194542 856
rect 194710 711 197302 856
rect 197470 711 200062 856
rect 200230 711 203282 856
rect 203450 711 206042 856
rect 206210 711 208802 856
rect 208970 711 211562 856
rect 211730 711 214322 856
rect 214490 711 217082 856
rect 217250 711 219842 856
rect 220010 711 222602 856
rect 222770 711 225362 856
rect 225530 711 228122 856
rect 228290 711 230882 856
rect 231050 711 233642 856
rect 233810 711 236402 856
rect 236570 711 238078 856
<< metal3 >>
rect 0 238688 800 238808
rect 238798 238688 239598 238808
rect 0 234608 800 234728
rect 238798 234608 239598 234728
rect 0 230528 800 230648
rect 238798 230528 239598 230648
rect 0 226448 800 226568
rect 238798 226448 239598 226568
rect 0 222368 800 222488
rect 238798 222368 239598 222488
rect 0 218288 800 218408
rect 238798 218288 239598 218408
rect 0 214208 800 214328
rect 238798 214208 239598 214328
rect 0 210128 800 210248
rect 238798 210128 239598 210248
rect 0 206048 800 206168
rect 238798 206048 239598 206168
rect 0 201968 800 202088
rect 238798 201968 239598 202088
rect 238798 197888 239598 198008
rect 0 197208 800 197328
rect 238798 193808 239598 193928
rect 0 193128 800 193248
rect 238798 189728 239598 189848
rect 0 189048 800 189168
rect 238798 185648 239598 185768
rect 0 184968 800 185088
rect 238798 181568 239598 181688
rect 0 180888 800 181008
rect 238798 177488 239598 177608
rect 0 176808 800 176928
rect 238798 173408 239598 173528
rect 0 172728 800 172848
rect 238798 169328 239598 169448
rect 0 168648 800 168768
rect 238798 165248 239598 165368
rect 0 164568 800 164688
rect 238798 161168 239598 161288
rect 0 160488 800 160608
rect 238798 157088 239598 157208
rect 0 156408 800 156528
rect 238798 153008 239598 153128
rect 0 152328 800 152448
rect 238798 148928 239598 149048
rect 0 148248 800 148368
rect 238798 144848 239598 144968
rect 0 144168 800 144288
rect 0 140088 800 140208
rect 238798 140088 239598 140208
rect 0 136008 800 136128
rect 238798 136008 239598 136128
rect 0 131928 800 132048
rect 238798 131928 239598 132048
rect 0 127848 800 127968
rect 238798 127848 239598 127968
rect 0 123768 800 123888
rect 238798 123768 239598 123888
rect 0 119688 800 119808
rect 238798 119688 239598 119808
rect 0 115608 800 115728
rect 238798 115608 239598 115728
rect 0 111528 800 111648
rect 238798 111528 239598 111648
rect 0 107448 800 107568
rect 238798 107448 239598 107568
rect 0 103368 800 103488
rect 238798 103368 239598 103488
rect 238798 99288 239598 99408
rect 0 98608 800 98728
rect 238798 95208 239598 95328
rect 0 94528 800 94648
rect 238798 91128 239598 91248
rect 0 90448 800 90568
rect 238798 87048 239598 87168
rect 0 86368 800 86488
rect 238798 82968 239598 83088
rect 0 82288 800 82408
rect 238798 78888 239598 79008
rect 0 78208 800 78328
rect 238798 74808 239598 74928
rect 0 74128 800 74248
rect 238798 70728 239598 70848
rect 0 70048 800 70168
rect 238798 66648 239598 66768
rect 0 65968 800 66088
rect 238798 62568 239598 62688
rect 0 61888 800 62008
rect 238798 58488 239598 58608
rect 0 57808 800 57928
rect 238798 54408 239598 54528
rect 0 53728 800 53848
rect 238798 50328 239598 50448
rect 0 49648 800 49768
rect 238798 46248 239598 46368
rect 0 45568 800 45688
rect 0 41488 800 41608
rect 238798 41488 239598 41608
rect 0 37408 800 37528
rect 238798 37408 239598 37528
rect 0 33328 800 33448
rect 238798 33328 239598 33448
rect 0 29248 800 29368
rect 238798 29248 239598 29368
rect 0 25168 800 25288
rect 238798 25168 239598 25288
rect 0 21088 800 21208
rect 238798 21088 239598 21208
rect 0 17008 800 17128
rect 238798 17008 239598 17128
rect 0 12928 800 13048
rect 238798 12928 239598 13048
rect 0 8848 800 8968
rect 238798 8848 239598 8968
rect 0 4768 800 4888
rect 238798 4768 239598 4888
rect 238798 688 239598 808
<< obsm3 >>
rect 800 238888 238798 239597
rect 880 238608 238718 238888
rect 800 234808 238798 238608
rect 880 234528 238718 234808
rect 800 230728 238798 234528
rect 880 230448 238718 230728
rect 800 226648 238798 230448
rect 880 226368 238718 226648
rect 800 222568 238798 226368
rect 880 222288 238718 222568
rect 800 218488 238798 222288
rect 880 218208 238718 218488
rect 800 214408 238798 218208
rect 880 214128 238718 214408
rect 800 210328 238798 214128
rect 880 210048 238718 210328
rect 800 206248 238798 210048
rect 880 205968 238718 206248
rect 800 202168 238798 205968
rect 880 201888 238718 202168
rect 800 198088 238798 201888
rect 800 197808 238718 198088
rect 800 197408 238798 197808
rect 880 197128 238798 197408
rect 800 194008 238798 197128
rect 800 193728 238718 194008
rect 800 193328 238798 193728
rect 880 193048 238798 193328
rect 800 189928 238798 193048
rect 800 189648 238718 189928
rect 800 189248 238798 189648
rect 880 188968 238798 189248
rect 800 185848 238798 188968
rect 800 185568 238718 185848
rect 800 185168 238798 185568
rect 880 184888 238798 185168
rect 800 181768 238798 184888
rect 800 181488 238718 181768
rect 800 181088 238798 181488
rect 880 180808 238798 181088
rect 800 177688 238798 180808
rect 800 177408 238718 177688
rect 800 177008 238798 177408
rect 880 176728 238798 177008
rect 800 173608 238798 176728
rect 800 173328 238718 173608
rect 800 172928 238798 173328
rect 880 172648 238798 172928
rect 800 169528 238798 172648
rect 800 169248 238718 169528
rect 800 168848 238798 169248
rect 880 168568 238798 168848
rect 800 165448 238798 168568
rect 800 165168 238718 165448
rect 800 164768 238798 165168
rect 880 164488 238798 164768
rect 800 161368 238798 164488
rect 800 161088 238718 161368
rect 800 160688 238798 161088
rect 880 160408 238798 160688
rect 800 157288 238798 160408
rect 800 157008 238718 157288
rect 800 156608 238798 157008
rect 880 156328 238798 156608
rect 800 153208 238798 156328
rect 800 152928 238718 153208
rect 800 152528 238798 152928
rect 880 152248 238798 152528
rect 800 149128 238798 152248
rect 800 148848 238718 149128
rect 800 148448 238798 148848
rect 880 148168 238798 148448
rect 800 145048 238798 148168
rect 800 144768 238718 145048
rect 800 144368 238798 144768
rect 880 144088 238798 144368
rect 800 140288 238798 144088
rect 880 140008 238718 140288
rect 800 136208 238798 140008
rect 880 135928 238718 136208
rect 800 132128 238798 135928
rect 880 131848 238718 132128
rect 800 128048 238798 131848
rect 880 127768 238718 128048
rect 800 123968 238798 127768
rect 880 123688 238718 123968
rect 800 119888 238798 123688
rect 880 119608 238718 119888
rect 800 115808 238798 119608
rect 880 115528 238718 115808
rect 800 111728 238798 115528
rect 880 111448 238718 111728
rect 800 107648 238798 111448
rect 880 107368 238718 107648
rect 800 103568 238798 107368
rect 880 103288 238718 103568
rect 800 99488 238798 103288
rect 800 99208 238718 99488
rect 800 98808 238798 99208
rect 880 98528 238798 98808
rect 800 95408 238798 98528
rect 800 95128 238718 95408
rect 800 94728 238798 95128
rect 880 94448 238798 94728
rect 800 91328 238798 94448
rect 800 91048 238718 91328
rect 800 90648 238798 91048
rect 880 90368 238798 90648
rect 800 87248 238798 90368
rect 800 86968 238718 87248
rect 800 86568 238798 86968
rect 880 86288 238798 86568
rect 800 83168 238798 86288
rect 800 82888 238718 83168
rect 800 82488 238798 82888
rect 880 82208 238798 82488
rect 800 79088 238798 82208
rect 800 78808 238718 79088
rect 800 78408 238798 78808
rect 880 78128 238798 78408
rect 800 75008 238798 78128
rect 800 74728 238718 75008
rect 800 74328 238798 74728
rect 880 74048 238798 74328
rect 800 70928 238798 74048
rect 800 70648 238718 70928
rect 800 70248 238798 70648
rect 880 69968 238798 70248
rect 800 66848 238798 69968
rect 800 66568 238718 66848
rect 800 66168 238798 66568
rect 880 65888 238798 66168
rect 800 62768 238798 65888
rect 800 62488 238718 62768
rect 800 62088 238798 62488
rect 880 61808 238798 62088
rect 800 58688 238798 61808
rect 800 58408 238718 58688
rect 800 58008 238798 58408
rect 880 57728 238798 58008
rect 800 54608 238798 57728
rect 800 54328 238718 54608
rect 800 53928 238798 54328
rect 880 53648 238798 53928
rect 800 50528 238798 53648
rect 800 50248 238718 50528
rect 800 49848 238798 50248
rect 880 49568 238798 49848
rect 800 46448 238798 49568
rect 800 46168 238718 46448
rect 800 45768 238798 46168
rect 880 45488 238798 45768
rect 800 41688 238798 45488
rect 880 41408 238718 41688
rect 800 37608 238798 41408
rect 880 37328 238718 37608
rect 800 33528 238798 37328
rect 880 33248 238718 33528
rect 800 29448 238798 33248
rect 880 29168 238718 29448
rect 800 25368 238798 29168
rect 880 25088 238718 25368
rect 800 21288 238798 25088
rect 880 21008 238718 21288
rect 800 17208 238798 21008
rect 880 16928 238718 17208
rect 800 13128 238798 16928
rect 880 12848 238718 13128
rect 800 9048 238798 12848
rect 880 8768 238718 9048
rect 800 4968 238798 8768
rect 880 4688 238718 4968
rect 800 888 238798 4688
rect 800 715 238718 888
<< metal4 >>
rect 4208 2128 4528 239408
rect 9208 2128 9528 239408
rect 14208 2128 14528 239408
rect 19208 2128 19528 239408
rect 24208 2128 24528 239408
rect 29208 2128 29528 239408
rect 34208 218452 34528 239408
rect 39208 218452 39528 239408
rect 44208 218452 44528 239408
rect 49208 218452 49528 239408
rect 54208 218452 54528 239408
rect 59208 218452 59528 239408
rect 64208 218452 64528 239408
rect 69208 218452 69528 239408
rect 74208 218452 74528 239408
rect 79208 218452 79528 239408
rect 84208 218452 84528 239408
rect 89208 218452 89528 239408
rect 94208 218452 94528 239408
rect 99208 218452 99528 239408
rect 104208 218452 104528 239408
rect 109208 218452 109528 239408
rect 114208 218452 114528 239408
rect 119208 218452 119528 239408
rect 124208 218452 124528 239408
rect 129208 218452 129528 239408
rect 34208 2128 34528 137048
rect 39208 2128 39528 137048
rect 44208 2128 44528 137048
rect 49208 2128 49528 137048
rect 54208 2128 54528 137048
rect 59208 2128 59528 137048
rect 64208 2128 64528 137048
rect 69208 2128 69528 137048
rect 74208 2128 74528 137048
rect 79208 2128 79528 137048
rect 84208 2128 84528 137048
rect 89208 2128 89528 137048
rect 94208 2128 94528 137048
rect 99208 2128 99528 137048
rect 104208 2128 104528 137048
rect 109208 2128 109528 137048
rect 114208 2128 114528 137048
rect 119208 2128 119528 137048
rect 124208 2128 124528 137048
rect 129208 2128 129528 137048
rect 134208 2128 134528 239408
rect 139208 2128 139528 239408
rect 144208 2128 144528 239408
rect 149208 2128 149528 239408
rect 154208 2128 154528 239408
rect 159208 2128 159528 239408
rect 164208 2128 164528 239408
rect 169208 2128 169528 239408
rect 174208 2128 174528 239408
rect 179208 2128 179528 239408
rect 184208 2128 184528 239408
rect 189208 2128 189528 239408
rect 194208 2128 194528 239408
rect 199208 2128 199528 239408
rect 204208 2128 204528 239408
rect 209208 2128 209528 239408
rect 214208 2128 214528 239408
rect 219208 2128 219528 239408
rect 224208 2128 224528 239408
rect 229208 2128 229528 239408
rect 234208 2128 234528 239408
<< obsm4 >>
rect 31891 239488 173821 239597
rect 31891 218372 34128 239488
rect 34608 218372 39128 239488
rect 39608 218372 44128 239488
rect 44608 218372 49128 239488
rect 49608 218372 54128 239488
rect 54608 218372 59128 239488
rect 59608 218372 64128 239488
rect 64608 218372 69128 239488
rect 69608 218372 74128 239488
rect 74608 218372 79128 239488
rect 79608 218372 84128 239488
rect 84608 218372 89128 239488
rect 89608 218372 94128 239488
rect 94608 218372 99128 239488
rect 99608 218372 104128 239488
rect 104608 218372 109128 239488
rect 109608 218372 114128 239488
rect 114608 218372 119128 239488
rect 119608 218372 124128 239488
rect 124608 218372 129128 239488
rect 129608 218372 134128 239488
rect 31891 137128 134128 218372
rect 31891 2048 34128 137128
rect 34608 2048 39128 137128
rect 39608 2048 44128 137128
rect 44608 2048 49128 137128
rect 49608 2048 54128 137128
rect 54608 2048 59128 137128
rect 59608 2048 64128 137128
rect 64608 2048 69128 137128
rect 69608 2048 74128 137128
rect 74608 2048 79128 137128
rect 79608 2048 84128 137128
rect 84608 2048 89128 137128
rect 89608 2048 94128 137128
rect 94608 2048 99128 137128
rect 99608 2048 104128 137128
rect 104608 2048 109128 137128
rect 109608 2048 114128 137128
rect 114608 2048 119128 137128
rect 119608 2048 124128 137128
rect 124608 2048 129128 137128
rect 129608 2048 134128 137128
rect 134608 2048 139128 239488
rect 139608 2048 144128 239488
rect 144608 2048 149128 239488
rect 149608 2048 154128 239488
rect 154608 2048 159128 239488
rect 159608 2048 164128 239488
rect 164608 2048 169128 239488
rect 169608 2048 173821 239488
rect 31891 1803 173821 2048
<< metal5 >>
rect 1104 235068 238464 235388
rect 1104 219750 238464 220070
rect 1104 204432 238464 204752
rect 1104 189114 238464 189434
rect 1104 173796 238464 174116
rect 1104 158478 238464 158798
rect 1104 143160 238464 143480
rect 1104 127842 238464 128162
rect 1104 112524 238464 112844
rect 1104 97206 238464 97526
rect 1104 81888 238464 82208
rect 1104 66570 238464 66890
rect 1104 51252 238464 51572
rect 1104 35934 238464 36254
rect 1104 20616 238464 20936
rect 1104 5298 238464 5618
<< labels >>
rlabel metal2 s 28998 240942 29054 241742 6 clk_i
port 1 nsew signal input
rlabel metal3 s 238798 185648 239598 185768 6 debug_req_i
port 2 nsew signal input
rlabel metal2 s 231858 240942 231914 241742 6 eFPGA_delay_o[0]
port 3 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 eFPGA_delay_o[1]
port 4 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 eFPGA_delay_o[2]
port 5 nsew signal output
rlabel metal2 s 170678 240942 170734 241742 6 eFPGA_delay_o[3]
port 6 nsew signal output
rlabel metal2 s 87418 240942 87474 241742 6 eFPGA_en_o
port 7 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 eFPGA_fpga_done_i
port 8 nsew signal input
rlabel metal3 s 238798 177488 239598 177608 6 eFPGA_operand_a_o[0]
port 9 nsew signal output
rlabel metal3 s 238798 66648 239598 66768 6 eFPGA_operand_a_o[10]
port 10 nsew signal output
rlabel metal3 s 0 230528 800 230648 6 eFPGA_operand_a_o[11]
port 11 nsew signal output
rlabel metal2 s 145838 240942 145894 241742 6 eFPGA_operand_a_o[12]
port 12 nsew signal output
rlabel metal2 s 101218 240942 101274 241742 6 eFPGA_operand_a_o[13]
port 13 nsew signal output
rlabel metal3 s 238798 107448 239598 107568 6 eFPGA_operand_a_o[14]
port 14 nsew signal output
rlabel metal3 s 0 193128 800 193248 6 eFPGA_operand_a_o[15]
port 15 nsew signal output
rlabel metal2 s 94778 0 94834 800 6 eFPGA_operand_a_o[16]
port 16 nsew signal output
rlabel metal3 s 238798 123768 239598 123888 6 eFPGA_operand_a_o[17]
port 17 nsew signal output
rlabel metal2 s 1398 240942 1454 241742 6 eFPGA_operand_a_o[18]
port 18 nsew signal output
rlabel metal2 s 30838 0 30894 800 6 eFPGA_operand_a_o[19]
port 19 nsew signal output
rlabel metal2 s 15198 240942 15254 241742 6 eFPGA_operand_a_o[1]
port 20 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 eFPGA_operand_a_o[20]
port 21 nsew signal output
rlabel metal3 s 238798 161168 239598 161288 6 eFPGA_operand_a_o[21]
port 22 nsew signal output
rlabel metal3 s 238798 37408 239598 37528 6 eFPGA_operand_a_o[22]
port 23 nsew signal output
rlabel metal3 s 238798 140088 239598 140208 6 eFPGA_operand_a_o[23]
port 24 nsew signal output
rlabel metal2 s 78218 0 78274 800 6 eFPGA_operand_a_o[24]
port 25 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 eFPGA_operand_a_o[25]
port 26 nsew signal output
rlabel metal3 s 238798 17008 239598 17128 6 eFPGA_operand_a_o[26]
port 27 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 eFPGA_operand_a_o[27]
port 28 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 eFPGA_operand_a_o[28]
port 29 nsew signal output
rlabel metal2 s 165158 240942 165214 241742 6 eFPGA_operand_a_o[29]
port 30 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 eFPGA_operand_a_o[2]
port 31 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 eFPGA_operand_a_o[30]
port 32 nsew signal output
rlabel metal2 s 17958 240942 18014 241742 6 eFPGA_operand_a_o[31]
port 33 nsew signal output
rlabel metal2 s 179418 240942 179474 241742 6 eFPGA_operand_a_o[3]
port 34 nsew signal output
rlabel metal2 s 40498 240942 40554 241742 6 eFPGA_operand_a_o[4]
port 35 nsew signal output
rlabel metal2 s 220818 240942 220874 241742 6 eFPGA_operand_a_o[5]
port 36 nsew signal output
rlabel metal2 s 92938 240942 92994 241742 6 eFPGA_operand_a_o[6]
port 37 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 eFPGA_operand_a_o[7]
port 38 nsew signal output
rlabel metal2 s 156878 240942 156934 241742 6 eFPGA_operand_a_o[8]
port 39 nsew signal output
rlabel metal2 s 109958 240942 110014 241742 6 eFPGA_operand_a_o[9]
port 40 nsew signal output
rlabel metal2 s 189078 0 189134 800 6 eFPGA_operand_b_o[0]
port 41 nsew signal output
rlabel metal3 s 238798 87048 239598 87168 6 eFPGA_operand_b_o[10]
port 42 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 eFPGA_operand_b_o[11]
port 43 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 eFPGA_operand_b_o[12]
port 44 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 eFPGA_operand_b_o[13]
port 45 nsew signal output
rlabel metal2 s 4158 240942 4214 241742 6 eFPGA_operand_b_o[14]
port 46 nsew signal output
rlabel metal3 s 0 160488 800 160608 6 eFPGA_operand_b_o[15]
port 47 nsew signal output
rlabel metal2 s 50158 0 50214 800 6 eFPGA_operand_b_o[16]
port 48 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 eFPGA_operand_b_o[17]
port 49 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 eFPGA_operand_b_o[18]
port 50 nsew signal output
rlabel metal2 s 233698 0 233754 800 6 eFPGA_operand_b_o[19]
port 51 nsew signal output
rlabel metal2 s 195978 240942 196034 241742 6 eFPGA_operand_b_o[1]
port 52 nsew signal output
rlabel metal2 s 84658 240942 84714 241742 6 eFPGA_operand_b_o[20]
port 53 nsew signal output
rlabel metal2 s 95698 240942 95754 241742 6 eFPGA_operand_b_o[21]
port 54 nsew signal output
rlabel metal2 s 229098 240942 229154 241742 6 eFPGA_operand_b_o[22]
port 55 nsew signal output
rlabel metal3 s 238798 234608 239598 234728 6 eFPGA_operand_b_o[23]
port 56 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 eFPGA_operand_b_o[24]
port 57 nsew signal output
rlabel metal2 s 126518 240942 126574 241742 6 eFPGA_operand_b_o[25]
port 58 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 eFPGA_operand_b_o[26]
port 59 nsew signal output
rlabel metal3 s 238798 181568 239598 181688 6 eFPGA_operand_b_o[27]
port 60 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 eFPGA_operand_b_o[28]
port 61 nsew signal output
rlabel metal3 s 238798 165248 239598 165368 6 eFPGA_operand_b_o[29]
port 62 nsew signal output
rlabel metal2 s 57058 240942 57114 241742 6 eFPGA_operand_b_o[2]
port 63 nsew signal output
rlabel metal2 s 103058 0 103114 800 6 eFPGA_operand_b_o[30]
port 64 nsew signal output
rlabel metal3 s 238798 70728 239598 70848 6 eFPGA_operand_b_o[31]
port 65 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 eFPGA_operand_b_o[3]
port 66 nsew signal output
rlabel metal3 s 0 180888 800 181008 6 eFPGA_operand_b_o[4]
port 67 nsew signal output
rlabel metal3 s 238798 111528 239598 111648 6 eFPGA_operand_b_o[5]
port 68 nsew signal output
rlabel metal2 s 154118 240942 154174 241742 6 eFPGA_operand_b_o[6]
port 69 nsew signal output
rlabel metal2 s 204258 240942 204314 241742 6 eFPGA_operand_b_o[7]
port 70 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 eFPGA_operand_b_o[8]
port 71 nsew signal output
rlabel metal2 s 153198 0 153254 800 6 eFPGA_operand_b_o[9]
port 72 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 eFPGA_operator_o[0]
port 73 nsew signal output
rlabel metal2 s 20718 240942 20774 241742 6 eFPGA_operator_o[1]
port 74 nsew signal output
rlabel metal2 s 34518 240942 34574 241742 6 eFPGA_result_a_i[0]
port 75 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 eFPGA_result_a_i[10]
port 76 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 eFPGA_result_a_i[11]
port 77 nsew signal input
rlabel metal3 s 0 214208 800 214328 6 eFPGA_result_a_i[12]
port 78 nsew signal input
rlabel metal3 s 238798 218288 239598 218408 6 eFPGA_result_a_i[13]
port 79 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 eFPGA_result_a_i[14]
port 80 nsew signal input
rlabel metal3 s 238798 62568 239598 62688 6 eFPGA_result_a_i[15]
port 81 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 eFPGA_result_a_i[16]
port 82 nsew signal input
rlabel metal2 s 182178 240942 182234 241742 6 eFPGA_result_a_i[17]
port 83 nsew signal input
rlabel metal2 s 54298 240942 54354 241742 6 eFPGA_result_a_i[18]
port 84 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 eFPGA_result_a_i[19]
port 85 nsew signal input
rlabel metal3 s 238798 173408 239598 173528 6 eFPGA_result_a_i[1]
port 86 nsew signal input
rlabel metal2 s 201498 240942 201554 241742 6 eFPGA_result_a_i[20]
port 87 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 eFPGA_result_a_i[21]
port 88 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 eFPGA_result_a_i[22]
port 89 nsew signal input
rlabel metal3 s 238798 21088 239598 21208 6 eFPGA_result_a_i[23]
port 90 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 eFPGA_result_a_i[24]
port 91 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 eFPGA_result_a_i[25]
port 92 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 eFPGA_result_a_i[26]
port 93 nsew signal input
rlabel metal2 s 65338 240942 65394 241742 6 eFPGA_result_a_i[27]
port 94 nsew signal input
rlabel metal3 s 0 197208 800 197328 6 eFPGA_result_a_i[28]
port 95 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 eFPGA_result_a_i[29]
port 96 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 eFPGA_result_a_i[2]
port 97 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 eFPGA_result_a_i[30]
port 98 nsew signal input
rlabel metal2 s 115478 240942 115534 241742 6 eFPGA_result_a_i[31]
port 99 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 eFPGA_result_a_i[3]
port 100 nsew signal input
rlabel metal2 s 187698 240942 187754 241742 6 eFPGA_result_a_i[4]
port 101 nsew signal input
rlabel metal2 s 186318 0 186374 800 6 eFPGA_result_a_i[5]
port 102 nsew signal input
rlabel metal3 s 0 210128 800 210248 6 eFPGA_result_a_i[6]
port 103 nsew signal input
rlabel metal3 s 238798 136008 239598 136128 6 eFPGA_result_a_i[7]
port 104 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 eFPGA_result_a_i[8]
port 105 nsew signal input
rlabel metal2 s 215298 240942 215354 241742 6 eFPGA_result_a_i[9]
port 106 nsew signal input
rlabel metal2 s 46018 240942 46074 241742 6 eFPGA_result_b_i[0]
port 107 nsew signal input
rlabel metal3 s 238798 33328 239598 33448 6 eFPGA_result_b_i[10]
port 108 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 eFPGA_result_b_i[11]
port 109 nsew signal input
rlabel metal2 s 198738 240942 198794 241742 6 eFPGA_result_b_i[12]
port 110 nsew signal input
rlabel metal3 s 238798 103368 239598 103488 6 eFPGA_result_b_i[13]
port 111 nsew signal input
rlabel metal2 s 98458 240942 98514 241742 6 eFPGA_result_b_i[14]
port 112 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 eFPGA_result_b_i[15]
port 113 nsew signal input
rlabel metal3 s 238798 230528 239598 230648 6 eFPGA_result_b_i[16]
port 114 nsew signal input
rlabel metal2 s 62578 240942 62634 241742 6 eFPGA_result_b_i[17]
port 115 nsew signal input
rlabel metal3 s 238798 25168 239598 25288 6 eFPGA_result_b_i[18]
port 116 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 eFPGA_result_b_i[19]
port 117 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 eFPGA_result_b_i[1]
port 118 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 eFPGA_result_b_i[20]
port 119 nsew signal input
rlabel metal2 s 90178 240942 90234 241742 6 eFPGA_result_b_i[21]
port 120 nsew signal input
rlabel metal3 s 0 238688 800 238808 6 eFPGA_result_b_i[22]
port 121 nsew signal input
rlabel metal3 s 238798 222368 239598 222488 6 eFPGA_result_b_i[23]
port 122 nsew signal input
rlabel metal2 s 228178 0 228234 800 6 eFPGA_result_b_i[24]
port 123 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 eFPGA_result_b_i[25]
port 124 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 eFPGA_result_b_i[26]
port 125 nsew signal input
rlabel metal2 s 190458 240942 190514 241742 6 eFPGA_result_b_i[27]
port 126 nsew signal input
rlabel metal3 s 238798 115608 239598 115728 6 eFPGA_result_b_i[28]
port 127 nsew signal input
rlabel metal3 s 238798 193808 239598 193928 6 eFPGA_result_b_i[29]
port 128 nsew signal input
rlabel metal3 s 238798 201968 239598 202088 6 eFPGA_result_b_i[2]
port 129 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 eFPGA_result_b_i[30]
port 130 nsew signal input
rlabel metal2 s 9678 240942 9734 241742 6 eFPGA_result_b_i[31]
port 131 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 eFPGA_result_b_i[3]
port 132 nsew signal input
rlabel metal3 s 238798 8848 239598 8968 6 eFPGA_result_b_i[4]
port 133 nsew signal input
rlabel metal3 s 0 172728 800 172848 6 eFPGA_result_b_i[5]
port 134 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 eFPGA_result_b_i[6]
port 135 nsew signal input
rlabel metal2 s 169758 0 169814 800 6 eFPGA_result_b_i[7]
port 136 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 eFPGA_result_b_i[8]
port 137 nsew signal input
rlabel metal3 s 0 226448 800 226568 6 eFPGA_result_b_i[9]
port 138 nsew signal input
rlabel metal2 s 132038 240942 132094 241742 6 eFPGA_result_c_i[0]
port 139 nsew signal input
rlabel metal2 s 176658 240942 176714 241742 6 eFPGA_result_c_i[10]
port 140 nsew signal input
rlabel metal2 s 68098 240942 68154 241742 6 eFPGA_result_c_i[11]
port 141 nsew signal input
rlabel metal2 s 162398 240942 162454 241742 6 eFPGA_result_c_i[12]
port 142 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 eFPGA_result_c_i[13]
port 143 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 eFPGA_result_c_i[14]
port 144 nsew signal input
rlabel metal2 s 167918 240942 167974 241742 6 eFPGA_result_c_i[15]
port 145 nsew signal input
rlabel metal2 s 140318 240942 140374 241742 6 eFPGA_result_c_i[16]
port 146 nsew signal input
rlabel metal2 s 23478 240942 23534 241742 6 eFPGA_result_c_i[17]
port 147 nsew signal input
rlabel metal3 s 0 156408 800 156528 6 eFPGA_result_c_i[18]
port 148 nsew signal input
rlabel metal3 s 238798 119688 239598 119808 6 eFPGA_result_c_i[19]
port 149 nsew signal input
rlabel metal3 s 238798 148928 239598 149048 6 eFPGA_result_c_i[1]
port 150 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 eFPGA_result_c_i[20]
port 151 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 eFPGA_result_c_i[21]
port 152 nsew signal input
rlabel metal2 s 226338 240942 226394 241742 6 eFPGA_result_c_i[22]
port 153 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 eFPGA_result_c_i[23]
port 154 nsew signal input
rlabel metal3 s 238798 169328 239598 169448 6 eFPGA_result_c_i[24]
port 155 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 eFPGA_result_c_i[25]
port 156 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 eFPGA_result_c_i[26]
port 157 nsew signal input
rlabel metal3 s 0 123768 800 123888 6 eFPGA_result_c_i[27]
port 158 nsew signal input
rlabel metal2 s 159638 240942 159694 241742 6 eFPGA_result_c_i[28]
port 159 nsew signal input
rlabel metal2 s 70858 240942 70914 241742 6 eFPGA_result_c_i[29]
port 160 nsew signal input
rlabel metal2 s 31758 240942 31814 241742 6 eFPGA_result_c_i[2]
port 161 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 eFPGA_result_c_i[30]
port 162 nsew signal input
rlabel metal3 s 238798 78888 239598 79008 6 eFPGA_result_c_i[31]
port 163 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 eFPGA_result_c_i[3]
port 164 nsew signal input
rlabel metal2 s 51538 240942 51594 241742 6 eFPGA_result_c_i[4]
port 165 nsew signal input
rlabel metal3 s 0 201968 800 202088 6 eFPGA_result_c_i[5]
port 166 nsew signal input
rlabel metal3 s 238798 91128 239598 91248 6 eFPGA_result_c_i[6]
port 167 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 eFPGA_result_c_i[7]
port 168 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 eFPGA_result_c_i[8]
port 169 nsew signal input
rlabel metal2 s 73618 240942 73674 241742 6 eFPGA_result_c_i[9]
port 170 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 eFPGA_write_strobe_o
port 171 nsew signal output
rlabel metal2 s 76378 240942 76434 241742 6 ext_data_addr_i[0]
port 172 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 ext_data_addr_i[10]
port 173 nsew signal input
rlabel metal3 s 238798 688 239598 808 6 ext_data_addr_i[11]
port 174 nsew signal input
rlabel metal2 s 79138 240942 79194 241742 6 ext_data_addr_i[12]
port 175 nsew signal input
rlabel metal2 s 118238 240942 118294 241742 6 ext_data_addr_i[13]
port 176 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 ext_data_addr_i[14]
port 177 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 ext_data_addr_i[15]
port 178 nsew signal input
rlabel metal2 s 107198 240942 107254 241742 6 ext_data_addr_i[16]
port 179 nsew signal input
rlabel metal3 s 238798 74808 239598 74928 6 ext_data_addr_i[17]
port 180 nsew signal input
rlabel metal3 s 238798 157088 239598 157208 6 ext_data_addr_i[18]
port 181 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 ext_data_addr_i[19]
port 182 nsew signal input
rlabel metal3 s 0 189048 800 189168 6 ext_data_addr_i[1]
port 183 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 ext_data_addr_i[20]
port 184 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 ext_data_addr_i[21]
port 185 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 ext_data_addr_i[22]
port 186 nsew signal input
rlabel metal2 s 129278 240942 129334 241742 6 ext_data_addr_i[23]
port 187 nsew signal input
rlabel metal2 s 222658 0 222714 800 6 ext_data_addr_i[24]
port 188 nsew signal input
rlabel metal3 s 238798 50328 239598 50448 6 ext_data_addr_i[25]
port 189 nsew signal input
rlabel metal2 s 223578 240942 223634 241742 6 ext_data_addr_i[26]
port 190 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 ext_data_addr_i[27]
port 191 nsew signal input
rlabel metal2 s 48778 240942 48834 241742 6 ext_data_addr_i[28]
port 192 nsew signal input
rlabel metal2 s 236458 0 236514 800 6 ext_data_addr_i[29]
port 193 nsew signal input
rlabel metal2 s 134798 240942 134854 241742 6 ext_data_addr_i[2]
port 194 nsew signal input
rlabel metal3 s 0 234608 800 234728 6 ext_data_addr_i[30]
port 195 nsew signal input
rlabel metal2 s 81898 240942 81954 241742 6 ext_data_addr_i[31]
port 196 nsew signal input
rlabel metal2 s 478 0 534 800 6 ext_data_addr_i[3]
port 197 nsew signal input
rlabel metal2 s 59818 240942 59874 241742 6 ext_data_addr_i[4]
port 198 nsew signal input
rlabel metal3 s 0 218288 800 218408 6 ext_data_addr_i[5]
port 199 nsew signal input
rlabel metal2 s 184938 240942 184994 241742 6 ext_data_addr_i[6]
port 200 nsew signal input
rlabel metal2 s 43258 240942 43314 241742 6 ext_data_addr_i[7]
port 201 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 ext_data_addr_i[8]
port 202 nsew signal input
rlabel metal3 s 0 206048 800 206168 6 ext_data_addr_i[9]
port 203 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 ext_data_be_i[0]
port 204 nsew signal input
rlabel metal2 s 26238 240942 26294 241742 6 ext_data_be_i[1]
port 205 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 ext_data_be_i[2]
port 206 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 ext_data_be_i[3]
port 207 nsew signal input
rlabel metal3 s 0 164568 800 164688 6 ext_data_gnt_o
port 208 nsew signal output
rlabel metal3 s 238798 226448 239598 226568 6 ext_data_rdata_o[0]
port 209 nsew signal output
rlabel metal2 s 191838 0 191894 800 6 ext_data_rdata_o[10]
port 210 nsew signal output
rlabel metal3 s 0 168648 800 168768 6 ext_data_rdata_o[11]
port 211 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 ext_data_rdata_o[12]
port 212 nsew signal output
rlabel metal3 s 238798 58488 239598 58608 6 ext_data_rdata_o[13]
port 213 nsew signal output
rlabel metal2 s 175278 0 175334 800 6 ext_data_rdata_o[14]
port 214 nsew signal output
rlabel metal2 s 103978 240942 104034 241742 6 ext_data_rdata_o[15]
port 215 nsew signal output
rlabel metal2 s 194598 0 194654 800 6 ext_data_rdata_o[16]
port 216 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 ext_data_rdata_o[17]
port 217 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 ext_data_rdata_o[18]
port 218 nsew signal output
rlabel metal3 s 0 152328 800 152448 6 ext_data_rdata_o[19]
port 219 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 ext_data_rdata_o[1]
port 220 nsew signal output
rlabel metal2 s 197358 0 197414 800 6 ext_data_rdata_o[20]
port 221 nsew signal output
rlabel metal3 s 238798 127848 239598 127968 6 ext_data_rdata_o[21]
port 222 nsew signal output
rlabel metal2 s 151358 240942 151414 241742 6 ext_data_rdata_o[22]
port 223 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 ext_data_rdata_o[23]
port 224 nsew signal output
rlabel metal2 s 143078 240942 143134 241742 6 ext_data_rdata_o[24]
port 225 nsew signal output
rlabel metal2 s 193218 240942 193274 241742 6 ext_data_rdata_o[25]
port 226 nsew signal output
rlabel metal3 s 0 222368 800 222488 6 ext_data_rdata_o[26]
port 227 nsew signal output
rlabel metal2 s 37278 240942 37334 241742 6 ext_data_rdata_o[27]
port 228 nsew signal output
rlabel metal2 s 218058 240942 218114 241742 6 ext_data_rdata_o[28]
port 229 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 ext_data_rdata_o[29]
port 230 nsew signal output
rlabel metal3 s 238798 82968 239598 83088 6 ext_data_rdata_o[2]
port 231 nsew signal output
rlabel metal2 s 137558 240942 137614 241742 6 ext_data_rdata_o[30]
port 232 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 ext_data_rdata_o[31]
port 233 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 ext_data_rdata_o[3]
port 234 nsew signal output
rlabel metal3 s 238798 131928 239598 132048 6 ext_data_rdata_o[4]
port 235 nsew signal output
rlabel metal2 s 12438 240942 12494 241742 6 ext_data_rdata_o[5]
port 236 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 ext_data_rdata_o[6]
port 237 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 ext_data_rdata_o[7]
port 238 nsew signal output
rlabel metal3 s 238798 54408 239598 54528 6 ext_data_rdata_o[8]
port 239 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 ext_data_rdata_o[9]
port 240 nsew signal output
rlabel metal2 s 173898 240942 173954 241742 6 ext_data_req_i
port 241 nsew signal input
rlabel metal2 s 207018 240942 207074 241742 6 ext_data_rvalid_o
port 242 nsew signal output
rlabel metal2 s 6918 240942 6974 241742 6 ext_data_wdata_i[0]
port 243 nsew signal input
rlabel metal2 s 123758 240942 123814 241742 6 ext_data_wdata_i[10]
port 244 nsew signal input
rlabel metal3 s 238798 153008 239598 153128 6 ext_data_wdata_i[11]
port 245 nsew signal input
rlabel metal2 s 100298 0 100354 800 6 ext_data_wdata_i[12]
port 246 nsew signal input
rlabel metal2 s 212538 240942 212594 241742 6 ext_data_wdata_i[13]
port 247 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 ext_data_wdata_i[14]
port 248 nsew signal input
rlabel metal3 s 238798 99288 239598 99408 6 ext_data_wdata_i[15]
port 249 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 ext_data_wdata_i[16]
port 250 nsew signal input
rlabel metal2 s 148598 240942 148654 241742 6 ext_data_wdata_i[17]
port 251 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 ext_data_wdata_i[18]
port 252 nsew signal input
rlabel metal3 s 238798 144848 239598 144968 6 ext_data_wdata_i[19]
port 253 nsew signal input
rlabel metal3 s 238798 12928 239598 13048 6 ext_data_wdata_i[1]
port 254 nsew signal input
rlabel metal2 s 219898 0 219954 800 6 ext_data_wdata_i[20]
port 255 nsew signal input
rlabel metal3 s 238798 210128 239598 210248 6 ext_data_wdata_i[21]
port 256 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 ext_data_wdata_i[22]
port 257 nsew signal input
rlabel metal3 s 238798 238688 239598 238808 6 ext_data_wdata_i[23]
port 258 nsew signal input
rlabel metal3 s 238798 46248 239598 46368 6 ext_data_wdata_i[24]
port 259 nsew signal input
rlabel metal2 s 234618 240942 234674 241742 6 ext_data_wdata_i[25]
port 260 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 ext_data_wdata_i[26]
port 261 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 ext_data_wdata_i[27]
port 262 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 ext_data_wdata_i[28]
port 263 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 ext_data_wdata_i[29]
port 264 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 ext_data_wdata_i[2]
port 265 nsew signal input
rlabel metal2 s 209778 240942 209834 241742 6 ext_data_wdata_i[30]
port 266 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 ext_data_wdata_i[31]
port 267 nsew signal input
rlabel metal2 s 120998 240942 121054 241742 6 ext_data_wdata_i[3]
port 268 nsew signal input
rlabel metal3 s 238798 41488 239598 41608 6 ext_data_wdata_i[4]
port 269 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 ext_data_wdata_i[5]
port 270 nsew signal input
rlabel metal3 s 238798 206048 239598 206168 6 ext_data_wdata_i[6]
port 271 nsew signal input
rlabel metal2 s 237378 240942 237434 241742 6 ext_data_wdata_i[7]
port 272 nsew signal input
rlabel metal3 s 238798 29248 239598 29368 6 ext_data_wdata_i[8]
port 273 nsew signal input
rlabel metal3 s 238798 197888 239598 198008 6 ext_data_wdata_i[9]
port 274 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 ext_data_we_i
port 275 nsew signal input
rlabel metal3 s 238798 4768 239598 4888 6 fetch_enable_i
port 276 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 irq_ack_o
port 277 nsew signal output
rlabel metal2 s 183558 0 183614 800 6 irq_i
port 278 nsew signal input
rlabel metal3 s 238798 189728 239598 189848 6 irq_id_i[0]
port 279 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 irq_id_i[1]
port 280 nsew signal input
rlabel metal2 s 112718 240942 112774 241742 6 irq_id_i[2]
port 281 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 irq_id_i[3]
port 282 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 irq_id_i[4]
port 283 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 irq_id_o[0]
port 284 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 irq_id_o[1]
port 285 nsew signal output
rlabel metal3 s 238798 95208 239598 95328 6 irq_id_o[2]
port 286 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 irq_id_o[3]
port 287 nsew signal output
rlabel metal3 s 0 184968 800 185088 6 irq_id_o[4]
port 288 nsew signal output
rlabel metal3 s 238798 214208 239598 214328 6 reset
port 289 nsew signal input
rlabel metal4 s 234208 2128 234528 239408 6 VPWR
port 290 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 239408 6 VPWR
port 291 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 239408 6 VPWR
port 292 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 239408 6 VPWR
port 293 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 239408 6 VPWR
port 294 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 239408 6 VPWR
port 295 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 239408 6 VPWR
port 296 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 239408 6 VPWR
port 297 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 239408 6 VPWR
port 298 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 239408 6 VPWR
port 299 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 239408 6 VPWR
port 300 nsew power bidirectional
rlabel metal4 s 124208 218452 124528 239408 6 VPWR
port 301 nsew power bidirectional
rlabel metal4 s 114208 218452 114528 239408 6 VPWR
port 302 nsew power bidirectional
rlabel metal4 s 104208 218452 104528 239408 6 VPWR
port 303 nsew power bidirectional
rlabel metal4 s 94208 218452 94528 239408 6 VPWR
port 304 nsew power bidirectional
rlabel metal4 s 84208 218452 84528 239408 6 VPWR
port 305 nsew power bidirectional
rlabel metal4 s 74208 218452 74528 239408 6 VPWR
port 306 nsew power bidirectional
rlabel metal4 s 64208 218452 64528 239408 6 VPWR
port 307 nsew power bidirectional
rlabel metal4 s 54208 218452 54528 239408 6 VPWR
port 308 nsew power bidirectional
rlabel metal4 s 44208 218452 44528 239408 6 VPWR
port 309 nsew power bidirectional
rlabel metal4 s 34208 218452 34528 239408 6 VPWR
port 310 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 239408 6 VPWR
port 311 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 239408 6 VPWR
port 312 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 239408 6 VPWR
port 313 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 137048 6 VPWR
port 314 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 137048 6 VPWR
port 315 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 137048 6 VPWR
port 316 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 137048 6 VPWR
port 317 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 137048 6 VPWR
port 318 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 137048 6 VPWR
port 319 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 137048 6 VPWR
port 320 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 137048 6 VPWR
port 321 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 137048 6 VPWR
port 322 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 137048 6 VPWR
port 323 nsew power bidirectional
rlabel metal5 s 1104 219750 238464 220070 6 VPWR
port 324 nsew power bidirectional
rlabel metal5 s 1104 189114 238464 189434 6 VPWR
port 325 nsew power bidirectional
rlabel metal5 s 1104 158478 238464 158798 6 VPWR
port 326 nsew power bidirectional
rlabel metal5 s 1104 127842 238464 128162 6 VPWR
port 327 nsew power bidirectional
rlabel metal5 s 1104 97206 238464 97526 6 VPWR
port 328 nsew power bidirectional
rlabel metal5 s 1104 66570 238464 66890 6 VPWR
port 329 nsew power bidirectional
rlabel metal5 s 1104 35934 238464 36254 6 VPWR
port 330 nsew power bidirectional
rlabel metal5 s 1104 5298 238464 5618 6 VPWR
port 331 nsew power bidirectional
rlabel metal4 s 229208 2128 229528 239408 6 VGND
port 332 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 239408 6 VGND
port 333 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 239408 6 VGND
port 334 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 239408 6 VGND
port 335 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 239408 6 VGND
port 336 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 239408 6 VGND
port 337 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 239408 6 VGND
port 338 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 239408 6 VGND
port 339 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 239408 6 VGND
port 340 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 239408 6 VGND
port 341 nsew ground bidirectional
rlabel metal4 s 129208 218452 129528 239408 6 VGND
port 342 nsew ground bidirectional
rlabel metal4 s 119208 218452 119528 239408 6 VGND
port 343 nsew ground bidirectional
rlabel metal4 s 109208 218452 109528 239408 6 VGND
port 344 nsew ground bidirectional
rlabel metal4 s 99208 218452 99528 239408 6 VGND
port 345 nsew ground bidirectional
rlabel metal4 s 89208 218452 89528 239408 6 VGND
port 346 nsew ground bidirectional
rlabel metal4 s 79208 218452 79528 239408 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 69208 218452 69528 239408 6 VGND
port 348 nsew ground bidirectional
rlabel metal4 s 59208 218452 59528 239408 6 VGND
port 349 nsew ground bidirectional
rlabel metal4 s 49208 218452 49528 239408 6 VGND
port 350 nsew ground bidirectional
rlabel metal4 s 39208 218452 39528 239408 6 VGND
port 351 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 239408 6 VGND
port 352 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 239408 6 VGND
port 353 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 239408 6 VGND
port 354 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 137048 6 VGND
port 355 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 137048 6 VGND
port 356 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 137048 6 VGND
port 357 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 137048 6 VGND
port 358 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 137048 6 VGND
port 359 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 137048 6 VGND
port 360 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 137048 6 VGND
port 361 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 137048 6 VGND
port 362 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 137048 6 VGND
port 363 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 137048 6 VGND
port 364 nsew ground bidirectional
rlabel metal5 s 1104 235068 238464 235388 6 VGND
port 365 nsew ground bidirectional
rlabel metal5 s 1104 204432 238464 204752 6 VGND
port 366 nsew ground bidirectional
rlabel metal5 s 1104 173796 238464 174116 6 VGND
port 367 nsew ground bidirectional
rlabel metal5 s 1104 143160 238464 143480 6 VGND
port 368 nsew ground bidirectional
rlabel metal5 s 1104 112524 238464 112844 6 VGND
port 369 nsew ground bidirectional
rlabel metal5 s 1104 81888 238464 82208 6 VGND
port 370 nsew ground bidirectional
rlabel metal5 s 1104 51252 238464 51572 6 VGND
port 371 nsew ground bidirectional
rlabel metal5 s 1104 20616 238464 20936 6 VGND
port 372 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 239598 241742
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 76839396
string GDS_START 10542526
<< end >>

