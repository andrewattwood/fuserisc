* NGSPICE file created from wb_mem_split.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

.subckt wb_mem_split core_a_data_addr_o[0] core_a_data_addr_o[1] core_a_data_addr_o[2]
+ core_a_data_addr_o[3] core_a_data_addr_o[4] core_a_data_addr_o[5] core_a_data_addr_o[6]
+ core_a_data_addr_o[7] core_a_data_addr_o[8] core_a_data_addr_o[9] core_a_data_be_o[0]
+ core_a_data_be_o[1] core_a_data_be_o[2] core_a_data_be_o[3] core_a_data_rdata_i[0]
+ core_a_data_rdata_i[10] core_a_data_rdata_i[11] core_a_data_rdata_i[12] core_a_data_rdata_i[13]
+ core_a_data_rdata_i[14] core_a_data_rdata_i[15] core_a_data_rdata_i[16] core_a_data_rdata_i[17]
+ core_a_data_rdata_i[18] core_a_data_rdata_i[19] core_a_data_rdata_i[1] core_a_data_rdata_i[20]
+ core_a_data_rdata_i[21] core_a_data_rdata_i[22] core_a_data_rdata_i[23] core_a_data_rdata_i[24]
+ core_a_data_rdata_i[25] core_a_data_rdata_i[26] core_a_data_rdata_i[27] core_a_data_rdata_i[28]
+ core_a_data_rdata_i[29] core_a_data_rdata_i[2] core_a_data_rdata_i[30] core_a_data_rdata_i[31]
+ core_a_data_rdata_i[3] core_a_data_rdata_i[4] core_a_data_rdata_i[5] core_a_data_rdata_i[6]
+ core_a_data_rdata_i[7] core_a_data_rdata_i[8] core_a_data_rdata_i[9] core_a_data_req_o
+ core_a_data_rvalid_i core_a_data_wdata_o[0] core_a_data_wdata_o[10] core_a_data_wdata_o[11]
+ core_a_data_wdata_o[12] core_a_data_wdata_o[13] core_a_data_wdata_o[14] core_a_data_wdata_o[15]
+ core_a_data_wdata_o[16] core_a_data_wdata_o[17] core_a_data_wdata_o[18] core_a_data_wdata_o[19]
+ core_a_data_wdata_o[1] core_a_data_wdata_o[20] core_a_data_wdata_o[21] core_a_data_wdata_o[22]
+ core_a_data_wdata_o[23] core_a_data_wdata_o[24] core_a_data_wdata_o[25] core_a_data_wdata_o[26]
+ core_a_data_wdata_o[27] core_a_data_wdata_o[28] core_a_data_wdata_o[29] core_a_data_wdata_o[2]
+ core_a_data_wdata_o[30] core_a_data_wdata_o[31] core_a_data_wdata_o[3] core_a_data_wdata_o[4]
+ core_a_data_wdata_o[5] core_a_data_wdata_o[6] core_a_data_wdata_o[7] core_a_data_wdata_o[8]
+ core_a_data_wdata_o[9] core_a_data_we_o core_b_data_addr_o[0] core_b_data_addr_o[1]
+ core_b_data_addr_o[2] core_b_data_addr_o[3] core_b_data_addr_o[4] core_b_data_addr_o[5]
+ core_b_data_addr_o[6] core_b_data_addr_o[7] core_b_data_addr_o[8] core_b_data_addr_o[9]
+ core_b_data_be_o[0] core_b_data_be_o[1] core_b_data_be_o[2] core_b_data_be_o[3]
+ core_b_data_rdata_i[0] core_b_data_rdata_i[10] core_b_data_rdata_i[11] core_b_data_rdata_i[12]
+ core_b_data_rdata_i[13] core_b_data_rdata_i[14] core_b_data_rdata_i[15] core_b_data_rdata_i[16]
+ core_b_data_rdata_i[17] core_b_data_rdata_i[18] core_b_data_rdata_i[19] core_b_data_rdata_i[1]
+ core_b_data_rdata_i[20] core_b_data_rdata_i[21] core_b_data_rdata_i[22] core_b_data_rdata_i[23]
+ core_b_data_rdata_i[24] core_b_data_rdata_i[25] core_b_data_rdata_i[26] core_b_data_rdata_i[27]
+ core_b_data_rdata_i[28] core_b_data_rdata_i[29] core_b_data_rdata_i[2] core_b_data_rdata_i[30]
+ core_b_data_rdata_i[31] core_b_data_rdata_i[3] core_b_data_rdata_i[4] core_b_data_rdata_i[5]
+ core_b_data_rdata_i[6] core_b_data_rdata_i[7] core_b_data_rdata_i[8] core_b_data_rdata_i[9]
+ core_b_data_req_o core_b_data_rvalid_i core_b_data_wdata_o[0] core_b_data_wdata_o[10]
+ core_b_data_wdata_o[11] core_b_data_wdata_o[12] core_b_data_wdata_o[13] core_b_data_wdata_o[14]
+ core_b_data_wdata_o[15] core_b_data_wdata_o[16] core_b_data_wdata_o[17] core_b_data_wdata_o[18]
+ core_b_data_wdata_o[19] core_b_data_wdata_o[1] core_b_data_wdata_o[20] core_b_data_wdata_o[21]
+ core_b_data_wdata_o[22] core_b_data_wdata_o[23] core_b_data_wdata_o[24] core_b_data_wdata_o[25]
+ core_b_data_wdata_o[26] core_b_data_wdata_o[27] core_b_data_wdata_o[28] core_b_data_wdata_o[29]
+ core_b_data_wdata_o[2] core_b_data_wdata_o[30] core_b_data_wdata_o[31] core_b_data_wdata_o[3]
+ core_b_data_wdata_o[4] core_b_data_wdata_o[5] core_b_data_wdata_o[6] core_b_data_wdata_o[7]
+ core_b_data_wdata_o[8] core_b_data_wdata_o[9] core_b_data_we_o wb_data_addr_i[0]
+ wb_data_addr_i[10] wb_data_addr_i[1] wb_data_addr_i[2] wb_data_addr_i[3] wb_data_addr_i[4]
+ wb_data_addr_i[5] wb_data_addr_i[6] wb_data_addr_i[7] wb_data_addr_i[8] wb_data_addr_i[9]
+ wb_data_be_i[0] wb_data_be_i[1] wb_data_be_i[2] wb_data_be_i[3] wb_data_rdata_o[0]
+ wb_data_rdata_o[10] wb_data_rdata_o[11] wb_data_rdata_o[12] wb_data_rdata_o[13]
+ wb_data_rdata_o[14] wb_data_rdata_o[15] wb_data_rdata_o[16] wb_data_rdata_o[17]
+ wb_data_rdata_o[18] wb_data_rdata_o[19] wb_data_rdata_o[1] wb_data_rdata_o[20] wb_data_rdata_o[21]
+ wb_data_rdata_o[22] wb_data_rdata_o[23] wb_data_rdata_o[24] wb_data_rdata_o[25]
+ wb_data_rdata_o[26] wb_data_rdata_o[27] wb_data_rdata_o[28] wb_data_rdata_o[29]
+ wb_data_rdata_o[2] wb_data_rdata_o[30] wb_data_rdata_o[31] wb_data_rdata_o[3] wb_data_rdata_o[4]
+ wb_data_rdata_o[5] wb_data_rdata_o[6] wb_data_rdata_o[7] wb_data_rdata_o[8] wb_data_rdata_o[9]
+ wb_data_rvalid_o wb_data_wdata_i[0] wb_data_wdata_i[10] wb_data_wdata_i[11] wb_data_wdata_i[12]
+ wb_data_wdata_i[13] wb_data_wdata_i[14] wb_data_wdata_i[15] wb_data_wdata_i[16]
+ wb_data_wdata_i[17] wb_data_wdata_i[18] wb_data_wdata_i[19] wb_data_wdata_i[1] wb_data_wdata_i[20]
+ wb_data_wdata_i[21] wb_data_wdata_i[22] wb_data_wdata_i[23] wb_data_wdata_i[24]
+ wb_data_wdata_i[25] wb_data_wdata_i[26] wb_data_wdata_i[27] wb_data_wdata_i[28]
+ wb_data_wdata_i[29] wb_data_wdata_i[2] wb_data_wdata_i[30] wb_data_wdata_i[31] wb_data_wdata_i[3]
+ wb_data_wdata_i[4] wb_data_wdata_i[5] wb_data_wdata_i[6] wb_data_wdata_i[7] wb_data_wdata_i[8]
+ wb_data_wdata_i[9] wb_data_we_i wbs_cyc_i wbs_stb_i VPWR VGND
XFILLER_39_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__274__A0 _274_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input92_A wb_data_wdata_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__113__B _206_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__265__A0 input5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__275__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_277_ _277_/A0 _277_/A1 _281_/S VGND VGND VPWR VPWR _277_/X sky130_fd_sc_hd__mux2_2
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput231 _278_/X VGND VGND VPWR VPWR wb_data_rdata_o[26] sky130_fd_sc_hd__clkbuf_2
Xoutput242 _259_/X VGND VGND VPWR VPWR wb_data_rdata_o[7] sky130_fd_sc_hd__clkbuf_2
Xoutput220 _268_/X VGND VGND VPWR VPWR wb_data_rdata_o[16] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_200_ _201_/A _200_/B VGND VGND VPWR VPWR _200_/Y sky130_fd_sc_hd__nor2_2
XFILLER_11_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_131_ _131_/A VGND VGND VPWR VPWR _217_/B sky130_fd_sc_hd__inv_2
XFILLER_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input55_A core_b_data_rdata_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output211_A _134_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__119__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_114_ _114_/A VGND VGND VPWR VPWR _207_/B sky130_fd_sc_hd__inv_2
XANTENNA_output161_A _216_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__283__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__206__B _206_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__222__A _223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input18_A core_a_data_rdata_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__278__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__217__A _218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__127__A _127_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input85_A wb_data_wdata_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__265__A1 _265_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__256__A1 _256_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_276_ _276_/A0 _276_/A1 _283_/S VGND VGND VPWR VPWR _276_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput221 _269_/X VGND VGND VPWR VPWR wb_data_rdata_o[17] sky130_fd_sc_hd__clkbuf_2
Xoutput210 _132_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput232 _279_/X VGND VGND VPWR VPWR wb_data_rdata_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput243 _260_/X VGND VGND VPWR VPWR wb_data_rdata_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_130_ _134_/A _216_/B VGND VGND VPWR VPWR _130_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input48_A core_b_data_rdata_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output204_A _185_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_259_ _259_/A0 _259_/A1 _281_/S VGND VGND VPWR VPWR _259_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input102_A wb_data_wdata_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_113_ _115_/A _206_/B VGND VGND VPWR VPWR _113_/Y sky130_fd_sc_hd__nor2_2
XFILLER_11_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 wb_data_wdata_i[6] VGND VGND VPWR VPWR _127_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output117_A _188_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input30_A core_a_data_rdata_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__143__A _143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input78_A wb_data_be_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_275_ _275_/A0 _275_/A1 _284_/S VGND VGND VPWR VPWR _275_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput200 _178_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput244 _261_/X VGND VGND VPWR VPWR wb_data_rdata_o[9] sky130_fd_sc_hd__clkbuf_2
Xoutput222 _270_/X VGND VGND VPWR VPWR wb_data_rdata_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput233 _280_/X VGND VGND VPWR VPWR wb_data_rdata_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput211 _134_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_189_ _191_/A _189_/B VGND VGND VPWR VPWR _189_/Y sky130_fd_sc_hd__nor2_4
X_258_ _258_/A0 _258_/A1 _284_/S VGND VGND VPWR VPWR _258_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__151__A _151_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_112_ _112_/A VGND VGND VPWR VPWR _206_/B sky130_fd_sc_hd__inv_2
XANTENNA_input60_A core_b_data_rdata_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output147_A _237_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput100 wb_data_wdata_i[26] VGND VGND VPWR VPWR _173_/A sky130_fd_sc_hd__buf_1
XANTENNA__277__A0 _277_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput111 wb_data_wdata_i[7] VGND VGND VPWR VPWR _129_/A sky130_fd_sc_hd__buf_1
XANTENNA_input23_A core_a_data_rdata_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__268__A0 input8/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output227_A _274_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_274_ _274_/A0 _274_/A1 _283_/S VGND VGND VPWR VPWR _274_/X sky130_fd_sc_hd__mux2_2
XANTENNA_input90_A wb_data_wdata_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput212 _251_/Y VGND VGND VPWR VPWR core_b_data_we_o sky130_fd_sc_hd__clkbuf_2
Xoutput223 _271_/X VGND VGND VPWR VPWR wb_data_rdata_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput201 _180_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_9_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput234 _281_/X VGND VGND VPWR VPWR wb_data_rdata_o[29] sky130_fd_sc_hd__clkbuf_2
Xoutput245 _284_/X VGND VGND VPWR VPWR wb_data_rvalid_o sky130_fd_sc_hd__clkbuf_2
XFILLER_23_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_257_ _257_/A0 _257_/A1 _284_/S VGND VGND VPWR VPWR _257_/X sky130_fd_sc_hd__mux2_4
X_188_ _191_/A _188_/B VGND VGND VPWR VPWR _188_/Y sky130_fd_sc_hd__nor2_2
XFILLER_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_111_ _115_/A _204_/B VGND VGND VPWR VPWR _111_/Y sky130_fd_sc_hd__nor2_4
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input53_A core_b_data_rdata_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__157__A _157_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput112 wb_data_wdata_i[8] VGND VGND VPWR VPWR _131_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput101 wb_data_wdata_i[27] VGND VGND VPWR VPWR _175_/A sky130_fd_sc_hd__buf_2
XANTENNA_input16_A core_a_data_rdata_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input8_A core_a_data_rdata_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__259__A1 _259_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__170__A _170_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_273_ _273_/A0 _273_/A1 _284_/S VGND VGND VPWR VPWR _273_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input83_A wb_data_wdata_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput202 _119_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput235 _254_/X VGND VGND VPWR VPWR wb_data_rdata_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput213 _252_/X VGND VGND VPWR VPWR wb_data_rdata_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput224 _253_/X VGND VGND VPWR VPWR wb_data_rdata_o[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_187_ _202_/A VGND VGND VPWR VPWR _191_/A sky130_fd_sc_hd__buf_4
X_256_ _256_/A0 _256_/A1 _284_/S VGND VGND VPWR VPWR _256_/X sky130_fd_sc_hd__mux2_2
XFILLER_6_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_110_ _110_/A VGND VGND VPWR VPWR _204_/B sky130_fd_sc_hd__inv_2
XANTENNA_input46_A core_b_data_rdata_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output202_A _119_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_239_ _239_/A _239_/B VGND VGND VPWR VPWR _239_/Y sky130_fd_sc_hd__nor2_2
XFILLER_30_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input100_A wb_data_wdata_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output152_A _243_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput113 wb_data_wdata_i[9] VGND VGND VPWR VPWR _133_/A sky130_fd_sc_hd__buf_1
Xinput102 wb_data_wdata_i[28] VGND VGND VPWR VPWR _177_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__168__A _168_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__078__A _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_272_ _272_/A0 _272_/A1 _284_/S VGND VGND VPWR VPWR _272_/X sky130_fd_sc_hd__mux2_2
XANTENNA_input76_A wb_data_addr_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output232_A _279_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput203 _183_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[30] sky130_fd_sc_hd__clkbuf_2
Xoutput214 _262_/X VGND VGND VPWR VPWR wb_data_rdata_o[10] sky130_fd_sc_hd__clkbuf_2
Xoutput225 _272_/X VGND VGND VPWR VPWR wb_data_rdata_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput236 _282_/X VGND VGND VPWR VPWR wb_data_rdata_o[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_23_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__091__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_255_ _255_/A0 _255_/A1 _281_/S VGND VGND VPWR VPWR _255_/X sky130_fd_sc_hd__mux2_1
XFILLER_43_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_186_ _283_/S VGND VGND VPWR VPWR _202_/A sky130_fd_sc_hd__buf_1
XFILLER_6_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__086__A _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input39_A core_b_data_rdata_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_169_ _171_/A _238_/B VGND VGND VPWR VPWR _169_/Y sky130_fd_sc_hd__nor2_1
X_238_ _239_/A _238_/B VGND VGND VPWR VPWR _238_/Y sky130_fd_sc_hd__nor2_4
XFILLER_30_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output145_A _234_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput103 wb_data_wdata_i[29] VGND VGND VPWR VPWR _179_/A sky130_fd_sc_hd__buf_1
XFILLER_44_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput114 wb_data_we_i VGND VGND VPWR VPWR _248_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__184__A _184_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input21_A core_a_data_rdata_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__179__A _179_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_271_ _271_/A0 _271_/A1 _284_/S VGND VGND VPWR VPWR _271_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input69_A wb_data_addr_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output225_A _272_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput215 _263_/X VGND VGND VPWR VPWR wb_data_rdata_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput226 _273_/X VGND VGND VPWR VPWR wb_data_rdata_o[21] sky130_fd_sc_hd__clkbuf_2
Xoutput237 _283_/X VGND VGND VPWR VPWR wb_data_rdata_o[31] sky130_fd_sc_hd__clkbuf_2
Xoutput204 _185_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_254_ _254_/A0 _254_/A1 _283_/S VGND VGND VPWR VPWR _254_/X sky130_fd_sc_hd__mux2_1
X_185_ _251_/A _247_/B VGND VGND VPWR VPWR _185_/Y sky130_fd_sc_hd__nor2_4
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_237_ _239_/A _237_/B VGND VGND VPWR VPWR _237_/Y sky130_fd_sc_hd__nor2_4
X_168_ _168_/A VGND VGND VPWR VPWR _238_/B sky130_fd_sc_hd__inv_2
XFILLER_30_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ _099_/A VGND VGND VPWR VPWR _198_/B sky130_fd_sc_hd__inv_2
XFILLER_41_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input51_A core_b_data_rdata_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput115 wbs_cyc_i VGND VGND VPWR VPWR _250_/A sky130_fd_sc_hd__buf_1
XFILLER_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput104 wb_data_wdata_i[2] VGND VGND VPWR VPWR _118_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input99_A wb_data_wdata_i[25] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input14_A core_a_data_rdata_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__195__A _196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input6_A core_a_data_rdata_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_270_ _270_/A0 _270_/A1 _283_/S VGND VGND VPWR VPWR _270_/X sky130_fd_sc_hd__mux2_2
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput205 _121_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_43_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput216 _264_/X VGND VGND VPWR VPWR wb_data_rdata_o[12] sky130_fd_sc_hd__clkbuf_2
XFILLER_13_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput227 _274_/X VGND VGND VPWR VPWR wb_data_rdata_o[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput238 _255_/X VGND VGND VPWR VPWR wb_data_rdata_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_2_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input116_A wbs_stb_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_184_ _184_/A VGND VGND VPWR VPWR _247_/B sky130_fd_sc_hd__inv_2
XANTENNA_input81_A wb_data_be_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_253_ _253_/A0 _253_/A1 _284_/S VGND VGND VPWR VPWR _253_/X sky130_fd_sc_hd__mux2_2
XFILLER_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output168_A _088_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_167_ _171_/A _237_/B VGND VGND VPWR VPWR _167_/Y sky130_fd_sc_hd__nor2_1
X_236_ _239_/A _236_/B VGND VGND VPWR VPWR _236_/Y sky130_fd_sc_hd__nor2_2
X_098_ _107_/A VGND VGND VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input44_A core_b_data_rdata_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output200_A _178_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_219_ _224_/A VGND VGND VPWR VPWR _223_/A sky130_fd_sc_hd__buf_4
XFILLER_7_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__198__A _201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput116 wbs_stb_i VGND VGND VPWR VPWR _250_/B sky130_fd_sc_hd__buf_1
XFILLER_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput105 wb_data_wdata_i[30] VGND VGND VPWR VPWR _182_/A sky130_fd_sc_hd__buf_1
XFILLER_44_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output150_A _241_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__270__A0 _270_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__261__A0 _261_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput206 _123_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput228 _275_/X VGND VGND VPWR VPWR wb_data_rdata_o[23] sky130_fd_sc_hd__clkbuf_2
Xoutput217 _265_/X VGND VGND VPWR VPWR wb_data_rdata_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput239 _256_/X VGND VGND VPWR VPWR wb_data_rdata_o[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input109_A wb_data_wdata_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_252_ input1/X _252_/A1 _281_/S VGND VGND VPWR VPWR _252_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input74_A wb_data_addr_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_183_ _251_/A _246_/B VGND VGND VPWR VPWR _183_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output230_A _277_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_235_ _245_/A VGND VGND VPWR VPWR _239_/A sky130_fd_sc_hd__clkbuf_4
X_166_ _166_/A VGND VGND VPWR VPWR _237_/B sky130_fd_sc_hd__inv_2
X_097_ _097_/A _196_/B VGND VGND VPWR VPWR _097_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_output180_A _113_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input37_A core_b_data_rdata_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_218_ _218_/A _218_/B VGND VGND VPWR VPWR _218_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_149_ _149_/A VGND VGND VPWR VPWR _227_/B sky130_fd_sc_hd__inv_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput106 wb_data_wdata_i[31] VGND VGND VPWR VPWR _184_/A sky130_fd_sc_hd__buf_1
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output143_A _207_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__270__A1 _270_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput229 _276_/X VGND VGND VPWR VPWR wb_data_rdata_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput218 _266_/X VGND VGND VPWR VPWR wb_data_rdata_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput207 _125_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__252__A1 _252_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_251_ _251_/A _251_/B VGND VGND VPWR VPWR _251_/Y sky130_fd_sc_hd__nor2_2
X_182_ _182_/A VGND VGND VPWR VPWR _246_/B sky130_fd_sc_hd__inv_2
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input67_A wb_data_addr_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__100__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_165_ _171_/A _236_/B VGND VGND VPWR VPWR _165_/Y sky130_fd_sc_hd__nor2_2
X_234_ _234_/A _234_/B VGND VGND VPWR VPWR _234_/Y sky130_fd_sc_hd__nor2_4
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_096_ _096_/A VGND VGND VPWR VPWR _196_/B sky130_fd_sc_hd__inv_2
XANTENNA_output173_A _100_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_217_ _218_/A _217_/B VGND VGND VPWR VPWR _217_/Y sky130_fd_sc_hd__nor2_2
X_148_ _152_/A _226_/B VGND VGND VPWR VPWR _148_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_079_ _153_/A VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__buf_1
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput107 wb_data_wdata_i[3] VGND VGND VPWR VPWR _120_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output136_A _223_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__254__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input97_A wb_data_wdata_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input12_A core_a_data_rdata_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput208 _128_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput219 _267_/X VGND VGND VPWR VPWR wb_data_rdata_o[15] sky130_fd_sc_hd__clkbuf_2
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input4_A core_a_data_rdata_i[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_250_ _250_/A _250_/B _250_/C VGND VGND VPWR VPWR _250_/X sky130_fd_sc_hd__and3_1
X_181_ _181_/A VGND VGND VPWR VPWR _251_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output216_A _264_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__262__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__201__A _201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input114_A wb_data_we_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_164_ _164_/A VGND VGND VPWR VPWR _236_/B sky130_fd_sc_hd__inv_2
X_233_ _234_/A _233_/B VGND VGND VPWR VPWR _233_/Y sky130_fd_sc_hd__nor2_4
X_095_ _097_/A _195_/B VGND VGND VPWR VPWR _095_/Y sky130_fd_sc_hd__nor2_2
XFILLER_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__257__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_078_ _283_/S VGND VGND VPWR VPWR _153_/A sky130_fd_sc_hd__inv_2
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_147_ _147_/A VGND VGND VPWR VPWR _226_/B sky130_fd_sc_hd__inv_2
X_216_ _218_/A _216_/B VGND VGND VPWR VPWR _216_/Y sky130_fd_sc_hd__nor2_2
XFILLER_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput108 wb_data_wdata_i[4] VGND VGND VPWR VPWR _122_/A sky130_fd_sc_hd__buf_1
XFILLER_29_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input42_A core_b_data_rdata_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__270__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput90 wb_data_wdata_i[17] VGND VGND VPWR VPWR _151_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__273__A0 _273_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__264__A0 input4/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__265__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__255__A0 _255_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__204__A _207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput209 _130_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[7] sky130_fd_sc_hd__clkbuf_2
XANTENNA__114__A _114_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_180_ _180_/A _244_/B VGND VGND VPWR VPWR _180_/Y sky130_fd_sc_hd__nor2_4
XFILLER_22_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_232_ _234_/A _232_/B VGND VGND VPWR VPWR _232_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_input107_A wb_data_wdata_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_163_ _181_/A VGND VGND VPWR VPWR _171_/A sky130_fd_sc_hd__clkbuf_2
X_094_ _094_/A VGND VGND VPWR VPWR _195_/B sky130_fd_sc_hd__inv_2
XANTENNA_input72_A wb_data_addr_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__273__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__212__A _213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_215_ _218_/A _215_/B VGND VGND VPWR VPWR _215_/Y sky130_fd_sc_hd__nor2_2
XFILLER_11_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_146_ _152_/A _225_/B VGND VGND VPWR VPWR _146_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__268__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput109 wb_data_wdata_i[5] VGND VGND VPWR VPWR _124_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__207__A _207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input35_A core_b_data_rdata_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_129_ _129_/A VGND VGND VPWR VPWR _216_/B sky130_fd_sc_hd__inv_2
XANTENNA__282__A1 _282_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput80 wb_data_be_i[2] VGND VGND VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
Xinput91 wb_data_wdata_i[18] VGND VGND VPWR VPWR _155_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output239_A _256_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__281__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__220__A _223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__276__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__215__A _218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__125__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_231_ _234_/A _231_/B VGND VGND VPWR VPWR _231_/Y sky130_fd_sc_hd__nor2_1
X_162_ _162_/A _234_/B VGND VGND VPWR VPWR _162_/Y sky130_fd_sc_hd__nor2_2
XFILLER_24_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input65_A core_b_data_rdata_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_093_ _097_/A _194_/B VGND VGND VPWR VPWR _093_/Y sky130_fd_sc_hd__nor2_2
XFILLER_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 core_a_data_rdata_i[0] VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__buf_1
XFILLER_24_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_214_ _224_/A VGND VGND VPWR VPWR _218_/A sky130_fd_sc_hd__buf_2
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_145_ _145_/A VGND VGND VPWR VPWR _225_/B sky130_fd_sc_hd__inv_2
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__284__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__207__B _207_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__223__A _223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput190 _158_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[19] sky130_fd_sc_hd__clkbuf_2
XANTENNA_input28_A core_a_data_rdata_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ _134_/A _215_/B VGND VGND VPWR VPWR _128_/Y sky130_fd_sc_hd__nor2_4
XFILLER_30_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__279__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput81 wb_data_be_i[3] VGND VGND VPWR VPWR _110_/A sky130_fd_sc_hd__buf_1
Xinput92 wb_data_wdata_i[19] VGND VGND VPWR VPWR _157_/A sky130_fd_sc_hd__clkbuf_2
Xinput70 wb_data_addr_i[2] VGND VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__218__A _218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input95_A wb_data_wdata_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input10_A core_a_data_rdata_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_repeater247_A _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__141__A _143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input2_A core_a_data_rdata_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_230_ _245_/A VGND VGND VPWR VPWR _234_/A sky130_fd_sc_hd__clkbuf_4
X_161_ _161_/A VGND VGND VPWR VPWR _234_/B sky130_fd_sc_hd__inv_2
XFILLER_24_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input58_A core_b_data_rdata_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_092_ _092_/A VGND VGND VPWR VPWR _194_/B sky130_fd_sc_hd__inv_2
XFILLER_6_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output214_A _262_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput2 core_a_data_rdata_i[10] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input112_A wb_data_wdata_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_144_ _144_/A VGND VGND VPWR VPWR _152_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_213_ _213_/A _213_/B VGND VGND VPWR VPWR _213_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_output164_A _249_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput191 _115_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[1] sky130_fd_sc_hd__clkbuf_2
XANTENNA__276__A0 _276_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput180 _113_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_127_ _127_/A VGND VGND VPWR VPWR _215_/B sky130_fd_sc_hd__inv_2
XFILLER_30_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__267__A0 input7/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput60 core_b_data_rdata_i[4] VGND VGND VPWR VPWR _256_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput93 wb_data_wdata_i[1] VGND VGND VPWR VPWR _114_/A sky130_fd_sc_hd__buf_1
Xinput82 wb_data_wdata_i[0] VGND VGND VPWR VPWR _112_/A sky130_fd_sc_hd__clkbuf_2
Xinput71 wb_data_addr_i[3] VGND VGND VPWR VPWR _087_/A sky130_fd_sc_hd__buf_2
XFILLER_40_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A core_b_data_rdata_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output127_A _200_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__229__A _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input88_A wb_data_wdata_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__139__A _143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output194_A _165_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_160_ _162_/A _233_/B VGND VGND VPWR VPWR _160_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_091_ _097_/A _193_/B VGND VGND VPWR VPWR _091_/Y sky130_fd_sc_hd__nor2_8
XFILLER_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output207_A _125_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput3 core_a_data_rdata_i[11] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__buf_1
XFILLER_24_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_212_ _213_/A _212_/B VGND VGND VPWR VPWR _212_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input105_A wb_data_wdata_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_143_ _143_/A _223_/B VGND VGND VPWR VPWR _143_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_input70_A wb_data_addr_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput170 _093_/Y VGND VGND VPWR VPWR core_b_data_addr_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput192 _160_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput181 _137_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[10] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_126_ _144_/A VGND VGND VPWR VPWR _134_/A sky130_fd_sc_hd__buf_2
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput50 core_b_data_rdata_i[24] VGND VGND VPWR VPWR _276_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput61 core_b_data_rdata_i[5] VGND VGND VPWR VPWR _257_/A1 sky130_fd_sc_hd__buf_1
Xinput72 wb_data_addr_i[4] VGND VGND VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_1
Xinput94 wb_data_wdata_i[20] VGND VGND VPWR VPWR _159_/A sky130_fd_sc_hd__buf_1
XFILLER_1_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput83 wb_data_wdata_i[10] VGND VGND VPWR VPWR _136_/A sky130_fd_sc_hd__buf_1
XFILLER_44_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__250__A _250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input33_A core_a_data_rvalid_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_109_ _115_/A _203_/B VGND VGND VPWR VPWR _109_/Y sky130_fd_sc_hd__nor2_2
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output237_A _283_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__155__A _155_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output187_A _150_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_090_ _090_/A VGND VGND VPWR VPWR _193_/B sky130_fd_sc_hd__inv_2
XFILLER_10_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput4 core_a_data_rdata_i[12] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_1
XFILLER_24_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_142_ _142_/A VGND VGND VPWR VPWR _223_/B sky130_fd_sc_hd__inv_2
XFILLER_42_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_211_ _213_/A _211_/B VGND VGND VPWR VPWR _211_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input63_A core_b_data_rdata_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput182 _139_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput193 _162_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[21] sky130_fd_sc_hd__clkbuf_2
Xoutput160 _215_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput171 _095_/Y VGND VGND VPWR VPWR core_b_data_addr_o[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__248__A _248_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_125_ _125_/A _213_/B VGND VGND VPWR VPWR _125_/Y sky130_fd_sc_hd__nor2_4
XFILLER_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput51 core_b_data_rdata_i[25] VGND VGND VPWR VPWR _277_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput62 core_b_data_rdata_i[6] VGND VGND VPWR VPWR _258_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput73 wb_data_addr_i[5] VGND VGND VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_2
Xinput95 wb_data_wdata_i[21] VGND VGND VPWR VPWR _161_/A sky130_fd_sc_hd__buf_1
Xinput40 core_b_data_rdata_i[15] VGND VGND VPWR VPWR _267_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput84 wb_data_wdata_i[11] VGND VGND VPWR VPWR _138_/A sky130_fd_sc_hd__buf_1
XFILLER_25_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__250__B _250_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input26_A core_a_data_rdata_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_108_ _108_/A VGND VGND VPWR VPWR _203_/B sky130_fd_sc_hd__inv_2
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__081__A _081_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input93_A wb_data_wdata_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput5 core_a_data_rdata_i[13] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_141_ _143_/A _222_/B VGND VGND VPWR VPWR _141_/Y sky130_fd_sc_hd__nor2_2
X_210_ _213_/A _210_/B VGND VGND VPWR VPWR _210_/Y sky130_fd_sc_hd__nor2_2
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__279__A0 _279_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input56_A core_b_data_rdata_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput150 _241_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[26] sky130_fd_sc_hd__clkbuf_2
Xoutput161 _216_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput183 _141_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput194 _165_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput172 _097_/Y VGND VGND VPWR VPWR core_b_data_addr_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input110_A wb_data_wdata_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_124_ _124_/A VGND VGND VPWR VPWR _213_/B sky130_fd_sc_hd__inv_2
XFILLER_7_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output162_A _217_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput52 core_b_data_rdata_i[26] VGND VGND VPWR VPWR _278_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput96 wb_data_wdata_i[22] VGND VGND VPWR VPWR _164_/A sky130_fd_sc_hd__clkbuf_1
Xinput74 wb_data_addr_i[6] VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__buf_1
Xinput30 core_a_data_rdata_i[7] VGND VGND VPWR VPWR _259_/A0 sky130_fd_sc_hd__buf_1
Xinput85 wb_data_wdata_i[12] VGND VGND VPWR VPWR _140_/A sky130_fd_sc_hd__clkbuf_1
Xinput63 core_b_data_rdata_i[7] VGND VGND VPWR VPWR _259_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput41 core_b_data_rdata_i[16] VGND VGND VPWR VPWR _268_/A1 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__084__A _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input19_A core_a_data_rdata_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_107_ _107_/A VGND VGND VPWR VPWR _115_/A sky130_fd_sc_hd__buf_2
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output125_A _198_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input86_A wb_data_wdata_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__092__A _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__177__A _177_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput6 core_a_data_rdata_i[14] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__087__A _087_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_140_ _140_/A VGND VGND VPWR VPWR _222_/B sky130_fd_sc_hd__inv_2
XANTENNA_input49_A core_b_data_rdata_i[23] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output205_A _121_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_269_ input9/X _269_/A1 _284_/S VGND VGND VPWR VPWR _269_/X sky130_fd_sc_hd__mux2_2
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput162 _217_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput184 _143_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput195 _167_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[23] sky130_fd_sc_hd__clkbuf_2
Xoutput151 _242_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput140 _228_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[17] sky130_fd_sc_hd__clkbuf_2
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput173 _100_/Y VGND VGND VPWR VPWR core_b_data_addr_o[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input103_A wb_data_wdata_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_123_ _125_/A _212_/B VGND VGND VPWR VPWR _123_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput31 core_a_data_rdata_i[8] VGND VGND VPWR VPWR _260_/A0 sky130_fd_sc_hd__buf_1
Xinput20 core_a_data_rdata_i[27] VGND VGND VPWR VPWR _279_/A0 sky130_fd_sc_hd__buf_1
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput86 wb_data_wdata_i[13] VGND VGND VPWR VPWR _142_/A sky130_fd_sc_hd__buf_1
Xinput53 core_b_data_rdata_i[27] VGND VGND VPWR VPWR _279_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput64 core_b_data_rdata_i[8] VGND VGND VPWR VPWR _260_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput97 wb_data_wdata_i[23] VGND VGND VPWR VPWR _166_/A sky130_fd_sc_hd__buf_1
XANTENNA__190__A _191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput42 core_b_data_rdata_i[17] VGND VGND VPWR VPWR _269_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput75 wb_data_addr_i[7] VGND VGND VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_106_ _106_/A _201_/B VGND VGND VPWR VPWR _106_/Y sky130_fd_sc_hd__nor2_2
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__095__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input31_A core_a_data_rdata_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output118_A _189_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input79_A wb_data_be_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput7 core_a_data_rdata_i[15] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__193__A _196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_268_ input8/X _268_/A1 _281_/S VGND VGND VPWR VPWR _268_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_199_ _201_/A _199_/B VGND VGND VPWR VPWR _199_/Y sky130_fd_sc_hd__nor2_2
XFILLER_37_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__188__A _191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput152 _243_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[28] sky130_fd_sc_hd__clkbuf_2
Xoutput141 _231_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput163 _218_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[9] sky130_fd_sc_hd__clkbuf_2
Xoutput196 _169_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput130 _204_/Y VGND VGND VPWR VPWR core_a_data_be_o[3] sky130_fd_sc_hd__clkbuf_2
Xoutput185 _146_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput174 _102_/Y VGND VGND VPWR VPWR core_b_data_addr_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_122_ _122_/A VGND VGND VPWR VPWR _212_/B sky130_fd_sc_hd__inv_2
XANTENNA_input61_A core_b_data_rdata_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output148_A _238_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput21 core_a_data_rdata_i[28] VGND VGND VPWR VPWR _280_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput10 core_a_data_rdata_i[18] VGND VGND VPWR VPWR _270_/A0 sky130_fd_sc_hd__buf_1
Xinput32 core_a_data_rdata_i[9] VGND VGND VPWR VPWR _261_/A0 sky130_fd_sc_hd__buf_2
Xinput54 core_b_data_rdata_i[28] VGND VGND VPWR VPWR _280_/A1 sky130_fd_sc_hd__clkbuf_4
Xinput43 core_b_data_rdata_i[18] VGND VGND VPWR VPWR _270_/A1 sky130_fd_sc_hd__buf_1
Xinput76 wb_data_addr_i[8] VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_2
Xinput65 core_b_data_rdata_i[9] VGND VGND VPWR VPWR _261_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput87 wb_data_wdata_i[14] VGND VGND VPWR VPWR _145_/A sky130_fd_sc_hd__clkbuf_1
Xinput98 wb_data_wdata_i[24] VGND VGND VPWR VPWR _168_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_37_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_105_ _105_/A VGND VGND VPWR VPWR _201_/B sky130_fd_sc_hd__inv_2
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input24_A core_a_data_rdata_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__196__A _196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output130_A _204_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input91_A wb_data_wdata_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_284_ _284_/A0 _284_/A1 _284_/S VGND VGND VPWR VPWR _284_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output178_A _111_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput8 core_a_data_rdata_i[16] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_267_ input7/X _267_/A1 _284_/S VGND VGND VPWR VPWR _267_/X sky130_fd_sc_hd__mux2_2
X_198_ _201_/A _198_/B VGND VGND VPWR VPWR _198_/Y sky130_fd_sc_hd__nor2_2
XFILLER_37_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput153 _244_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[29] sky130_fd_sc_hd__clkbuf_2
Xoutput131 _205_/X VGND VGND VPWR VPWR core_a_data_req_o sky130_fd_sc_hd__clkbuf_2
Xoutput197 _171_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[25] sky130_fd_sc_hd__clkbuf_2
Xoutput142 _232_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[19] sky130_fd_sc_hd__clkbuf_2
Xoutput175 _104_/Y VGND VGND VPWR VPWR core_b_data_be_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput120 _191_/Y VGND VGND VPWR VPWR core_a_data_addr_o[3] sky130_fd_sc_hd__clkbuf_2
Xoutput186 _148_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput164 _249_/Y VGND VGND VPWR VPWR core_a_data_we_o sky130_fd_sc_hd__clkbuf_2
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_121_ _125_/A _211_/B VGND VGND VPWR VPWR _121_/Y sky130_fd_sc_hd__nor2_8
XFILLER_23_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input54_A core_b_data_rdata_i[28] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output210_A _132_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput66 core_b_data_rvalid_i VGND VGND VPWR VPWR _284_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput22 core_a_data_rdata_i[29] VGND VGND VPWR VPWR _281_/A0 sky130_fd_sc_hd__buf_2
Xinput44 core_b_data_rdata_i[19] VGND VGND VPWR VPWR _271_/A1 sky130_fd_sc_hd__buf_1
Xinput11 core_a_data_rdata_i[19] VGND VGND VPWR VPWR _271_/A0 sky130_fd_sc_hd__buf_1
Xinput55 core_b_data_rdata_i[29] VGND VGND VPWR VPWR _281_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput33 core_a_data_rvalid_i VGND VGND VPWR VPWR _284_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput77 wb_data_addr_i[9] VGND VGND VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_1
Xinput88 wb_data_wdata_i[15] VGND VGND VPWR VPWR _147_/A sky130_fd_sc_hd__buf_1
Xinput99 wb_data_wdata_i[25] VGND VGND VPWR VPWR _170_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__199__A _201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_104_ _106_/A _200_/B VGND VGND VPWR VPWR _104_/Y sky130_fd_sc_hd__nor2_1
XFILLER_34_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input17_A core_a_data_rdata_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input9_A core_a_data_rdata_i[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_283_ _283_/A0 _283_/A1 _283_/S VGND VGND VPWR VPWR _283_/X sky130_fd_sc_hd__mux2_2
XFILLER_41_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input84_A wb_data_wdata_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output240_A _257_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 core_a_data_rdata_i[17] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__buf_1
XFILLER_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_266_ input6/X _266_/A1 _281_/S VGND VGND VPWR VPWR _266_/X sky130_fd_sc_hd__mux2_1
X_197_ _202_/A VGND VGND VPWR VPWR _201_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput143 _207_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput121 _193_/Y VGND VGND VPWR VPWR core_a_data_addr_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput132 _206_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput176 _106_/Y VGND VGND VPWR VPWR core_b_data_be_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput165 _082_/Y VGND VGND VPWR VPWR core_b_data_addr_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput154 _210_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput187 _150_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[16] sky130_fd_sc_hd__clkbuf_2
Xoutput198 _174_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[26] sky130_fd_sc_hd__clkbuf_2
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_120_ _120_/A VGND VGND VPWR VPWR _211_/B sky130_fd_sc_hd__inv_2
XFILLER_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input47_A core_b_data_rdata_i[21] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput45 core_b_data_rdata_i[1] VGND VGND VPWR VPWR _253_/A1 sky130_fd_sc_hd__buf_2
Xinput23 core_a_data_rdata_i[2] VGND VGND VPWR VPWR _254_/A0 sky130_fd_sc_hd__buf_1
X_249_ _250_/C _251_/B VGND VGND VPWR VPWR _249_/Y sky130_fd_sc_hd__nor2_4
Xinput67 wb_data_addr_i[0] VGND VGND VPWR VPWR _081_/A sky130_fd_sc_hd__buf_2
Xinput78 wb_data_be_i[0] VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_2
Xinput34 core_b_data_rdata_i[0] VGND VGND VPWR VPWR _252_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput56 core_b_data_rdata_i[2] VGND VGND VPWR VPWR _254_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput12 core_a_data_rdata_i[1] VGND VGND VPWR VPWR _253_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput89 wb_data_wdata_i[16] VGND VGND VPWR VPWR _149_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input101_A wb_data_wdata_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_103_ _103_/A VGND VGND VPWR VPWR _200_/B sky130_fd_sc_hd__inv_2
XFILLER_19_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__252__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_282_ _282_/A0 _282_/A1 _283_/S VGND VGND VPWR VPWR _282_/X sky130_fd_sc_hd__mux2_2
XFILLER_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input77_A wb_data_addr_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_196_ _196_/A _196_/B VGND VGND VPWR VPWR _196_/Y sky130_fd_sc_hd__nor2_1
X_265_ input5/X _265_/A1 _284_/S VGND VGND VPWR VPWR _265_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput166 _084_/Y VGND VGND VPWR VPWR core_b_data_addr_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput122 _194_/Y VGND VGND VPWR VPWR core_a_data_addr_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput177 _109_/Y VGND VGND VPWR VPWR core_b_data_be_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput144 _233_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[20] sky130_fd_sc_hd__clkbuf_2
Xoutput155 _246_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[30] sky130_fd_sc_hd__clkbuf_2
Xoutput133 _220_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[10] sky130_fd_sc_hd__clkbuf_2
Xoutput199 _176_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[27] sky130_fd_sc_hd__clkbuf_2
Xoutput188 _152_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[17] sky130_fd_sc_hd__clkbuf_2
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput13 core_a_data_rdata_i[20] VGND VGND VPWR VPWR _272_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput24 core_a_data_rdata_i[30] VGND VGND VPWR VPWR _282_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput79 wb_data_be_i[1] VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__buf_1
XANTENNA__260__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_179_ _179_/A VGND VGND VPWR VPWR _244_/B sky130_fd_sc_hd__inv_2
X_248_ _248_/A VGND VGND VPWR VPWR _251_/B sky130_fd_sc_hd__inv_2
Xinput46 core_b_data_rdata_i[20] VGND VGND VPWR VPWR _272_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput35 core_b_data_rdata_i[10] VGND VGND VPWR VPWR _262_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput57 core_b_data_rdata_i[30] VGND VGND VPWR VPWR _282_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput68 wb_data_addr_i[10] VGND VGND VPWR VPWR _281_/S sky130_fd_sc_hd__buf_6
XFILLER_6_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__281__A0 _281_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_102_ _106_/A _199_/B VGND VGND VPWR VPWR _102_/Y sky130_fd_sc_hd__nor2_2
XFILLER_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output146_A _236_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__255__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__254__A0 _254_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__104__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input22_A core_a_data_rdata_i[29] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_281_ _281_/A0 _281_/A1 _281_/S VGND VGND VPWR VPWR _281_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__263__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_264_ input4/X _264_/A1 _283_/S VGND VGND VPWR VPWR _264_/X sky130_fd_sc_hd__mux2_2
XFILLER_42_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_195_ _196_/A _195_/B VGND VGND VPWR VPWR _195_/Y sky130_fd_sc_hd__nor2_2
XFILLER_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__112__A _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__258__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput156 _247_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[31] sky130_fd_sc_hd__clkbuf_2
Xoutput189 _156_/Y VGND VGND VPWR VPWR core_b_data_wdata_o[18] sky130_fd_sc_hd__clkbuf_2
Xoutput123 _195_/Y VGND VGND VPWR VPWR core_a_data_addr_o[6] sky130_fd_sc_hd__clkbuf_2
Xoutput167 _086_/Y VGND VGND VPWR VPWR core_b_data_addr_o[2] sky130_fd_sc_hd__clkbuf_2
Xoutput145 _234_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[21] sky130_fd_sc_hd__clkbuf_2
Xoutput134 _221_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[11] sky130_fd_sc_hd__clkbuf_2
Xoutput178 _111_/Y VGND VGND VPWR VPWR core_b_data_be_o[3] sky130_fd_sc_hd__clkbuf_2
XFILLER_46_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput25 core_a_data_rdata_i[31] VGND VGND VPWR VPWR _283_/A0 sky130_fd_sc_hd__buf_1
X_247_ _250_/C _247_/B VGND VGND VPWR VPWR _247_/Y sky130_fd_sc_hd__nor2_1
XFILLER_30_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput36 core_b_data_rdata_i[11] VGND VGND VPWR VPWR _263_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput14 core_a_data_rdata_i[21] VGND VGND VPWR VPWR _273_/A0 sky130_fd_sc_hd__clkbuf_2
Xinput58 core_b_data_rdata_i[31] VGND VGND VPWR VPWR _283_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput69 wb_data_addr_i[1] VGND VGND VPWR VPWR _083_/A sky130_fd_sc_hd__buf_1
X_178_ _180_/A _243_/B VGND VGND VPWR VPWR _178_/Y sky130_fd_sc_hd__nor2_4
Xinput47 core_b_data_rdata_i[21] VGND VGND VPWR VPWR _273_/A1 sky130_fd_sc_hd__buf_1
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_101_ _101_/A VGND VGND VPWR VPWR _199_/B sky130_fd_sc_hd__inv_2
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input52_A core_b_data_rdata_i[26] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output139_A _227_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__263__A1 _263_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__271__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__254__A1 _254_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__210__A _213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__266__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__205__A _250_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input15_A core_a_data_rdata_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input7_A core_a_data_rdata_i[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_280_ _280_/A0 _280_/A1 _283_/S VGND VGND VPWR VPWR _280_/X sky130_fd_sc_hd__mux2_1
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output219_A _267_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output121_A _193_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A wb_data_wdata_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ input3/X _263_/A1 _284_/S VGND VGND VPWR VPWR _263_/X sky130_fd_sc_hd__mux2_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output169_A _091_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_194_ _196_/A _194_/B VGND VGND VPWR VPWR _194_/Y sky130_fd_sc_hd__nor2_2
XFILLER_6_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__274__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput179 _250_/X VGND VGND VPWR VPWR core_b_data_req_o sky130_fd_sc_hd__clkbuf_2
Xoutput135 _222_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[12] sky130_fd_sc_hd__clkbuf_2
Xoutput146 _236_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[22] sky130_fd_sc_hd__clkbuf_2
Xoutput157 _211_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[3] sky130_fd_sc_hd__clkbuf_2
Xoutput168 _088_/Y VGND VGND VPWR VPWR core_b_data_addr_o[3] sky130_fd_sc_hd__clkbuf_2
Xoutput124 _196_/Y VGND VGND VPWR VPWR core_a_data_addr_o[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_24_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__213__A _213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput37 core_b_data_rdata_i[12] VGND VGND VPWR VPWR _264_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput26 core_a_data_rdata_i[3] VGND VGND VPWR VPWR _255_/A0 sky130_fd_sc_hd__buf_1
Xinput48 core_b_data_rdata_i[22] VGND VGND VPWR VPWR _274_/A1 sky130_fd_sc_hd__clkbuf_1
X_177_ _177_/A VGND VGND VPWR VPWR _243_/B sky130_fd_sc_hd__inv_2
X_246_ _250_/C _246_/B VGND VGND VPWR VPWR _246_/Y sky130_fd_sc_hd__nor2_2
Xinput59 core_b_data_rdata_i[3] VGND VGND VPWR VPWR _255_/A1 sky130_fd_sc_hd__clkbuf_1
Xinput15 core_a_data_rdata_i[22] VGND VGND VPWR VPWR _274_/A0 sky130_fd_sc_hd__buf_1
XANTENNA__123__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__269__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__208__A _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_100_ _106_/A _198_/B VGND VGND VPWR VPWR _100_/Y sky130_fd_sc_hd__nor2_4
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input45_A core_b_data_rdata_i[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output201_A _180_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_229_ _283_/S VGND VGND VPWR VPWR _245_/A sky130_fd_sc_hd__buf_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output151_A _242_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__282__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__205__B _250_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__221__A _223_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output199_A _176_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__115__B _207_/B VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__277__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__216__A _218_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_193_ _196_/A _193_/B VGND VGND VPWR VPWR _193_/Y sky130_fd_sc_hd__nor2_4
X_262_ input2/X _262_/A1 _281_/S VGND VGND VPWR VPWR _262_/X sky130_fd_sc_hd__mux2_2
XPHY_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input75_A wb_data_addr_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput125 _198_/Y VGND VGND VPWR VPWR core_a_data_addr_o[8] sky130_fd_sc_hd__clkbuf_2
Xoutput136 _223_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[13] sky130_fd_sc_hd__clkbuf_2
Xoutput169 _091_/Y VGND VGND VPWR VPWR core_b_data_addr_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput158 _212_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[4] sky130_fd_sc_hd__clkbuf_2
Xoutput147 _237_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[23] sky130_fd_sc_hd__clkbuf_2
XANTENNA__284__A0 _284_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__275__A0 _275_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput38 core_b_data_rdata_i[13] VGND VGND VPWR VPWR _265_/A1 sky130_fd_sc_hd__clkbuf_2
Xinput16 core_a_data_rdata_i[23] VGND VGND VPWR VPWR _275_/A0 sky130_fd_sc_hd__clkbuf_2
X_245_ _245_/A VGND VGND VPWR VPWR _250_/C sky130_fd_sc_hd__buf_2
X_176_ _180_/A _242_/B VGND VGND VPWR VPWR _176_/Y sky130_fd_sc_hd__nor2_2
Xinput49 core_b_data_rdata_i[23] VGND VGND VPWR VPWR _275_/A1 sky130_fd_sc_hd__clkbuf_1
XANTENNA_output181_A _137_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput27 core_a_data_rdata_i[4] VGND VGND VPWR VPWR _256_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input38_A core_b_data_rdata_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_159_ _159_/A VGND VGND VPWR VPWR _233_/B sky130_fd_sc_hd__inv_2
X_228_ _228_/A _228_/B VGND VGND VPWR VPWR _228_/Y sky130_fd_sc_hd__nor2_2
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output144_A _233_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input20_A core_a_data_rdata_i[27] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__142__A _142_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_261_ _261_/A0 _261_/A1 _284_/S VGND VGND VPWR VPWR _261_/X sky130_fd_sc_hd__mux2_1
X_192_ _202_/A VGND VGND VPWR VPWR _196_/A sky130_fd_sc_hd__buf_4
XFILLER_22_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input68_A wb_data_addr_i[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output224_A _253_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__137__A _143_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput137 _225_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[14] sky130_fd_sc_hd__clkbuf_2
Xoutput159 _213_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[5] sky130_fd_sc_hd__clkbuf_2
Xoutput148 _238_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[24] sky130_fd_sc_hd__clkbuf_2
Xoutput126 _199_/Y VGND VGND VPWR VPWR core_a_data_addr_o[9] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__284__A1 _284_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_244_ _244_/A _244_/B VGND VGND VPWR VPWR _244_/Y sky130_fd_sc_hd__nor2_1
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput39 core_b_data_rdata_i[14] VGND VGND VPWR VPWR _266_/A1 sky130_fd_sc_hd__clkbuf_2
X_175_ _175_/A VGND VGND VPWR VPWR _242_/B sky130_fd_sc_hd__inv_2
Xinput28 core_a_data_rdata_i[5] VGND VGND VPWR VPWR _257_/A0 sky130_fd_sc_hd__clkbuf_1
Xinput17 core_a_data_rdata_i[24] VGND VGND VPWR VPWR _276_/A0 sky130_fd_sc_hd__buf_1
XANTENNA_output174_A _102_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__266__A1 _266_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_227_ _228_/A _227_/B VGND VGND VPWR VPWR _227_/Y sky130_fd_sc_hd__nor2_2
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_158_ _162_/A _232_/B VGND VGND VPWR VPWR _158_/Y sky130_fd_sc_hd__nor2_1
X_089_ _107_/A VGND VGND VPWR VPWR _097_/A sky130_fd_sc_hd__buf_4
XFILLER_10_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input50_A core_b_data_rdata_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output137_A _225_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input98_A wb_data_wdata_i[24] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input13_A core_a_data_rdata_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input5_A core_a_data_rdata_i[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_260_ _260_/A0 _260_/A1 _283_/S VGND VGND VPWR VPWR _260_/X sky130_fd_sc_hd__mux2_2
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_191_ _191_/A _191_/B VGND VGND VPWR VPWR _191_/Y sky130_fd_sc_hd__nor2_2
XFILLER_10_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput138 _226_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[15] sky130_fd_sc_hd__clkbuf_2
Xoutput127 _200_/Y VGND VGND VPWR VPWR core_a_data_be_o[0] sky130_fd_sc_hd__clkbuf_2
Xoutput149 _239_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input115_A wbs_cyc_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input80_A wb_data_be_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_243_ _244_/A _243_/B VGND VGND VPWR VPWR _243_/Y sky130_fd_sc_hd__nor2_2
Xinput18 core_a_data_rdata_i[25] VGND VGND VPWR VPWR _277_/A0 sky130_fd_sc_hd__clkbuf_2
XFILLER_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_174_ _180_/A _241_/B VGND VGND VPWR VPWR _174_/Y sky130_fd_sc_hd__nor2_2
Xinput29 core_a_data_rdata_i[6] VGND VGND VPWR VPWR _258_/A0 sky130_fd_sc_hd__buf_1
XFILLER_2_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_157_ _157_/A VGND VGND VPWR VPWR _232_/B sky130_fd_sc_hd__inv_2
X_226_ _228_/A _226_/B VGND VGND VPWR VPWR _226_/Y sky130_fd_sc_hd__nor2_2
X_088_ _088_/A _191_/B VGND VGND VPWR VPWR _088_/Y sky130_fd_sc_hd__nor2_2
XFILLER_21_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input43_A core_b_data_rdata_i[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_209_ _224_/A VGND VGND VPWR VPWR _213_/A sky130_fd_sc_hd__clkbuf_4
Xrepeater246 _283_/S VGND VGND VPWR VPWR _284_/S sky130_fd_sc_hd__buf_8
XFILLER_21_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output197_A _171_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_190_ _191_/A _190_/B VGND VGND VPWR VPWR _190_/Y sky130_fd_sc_hd__nor2_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput139 _227_/Y VGND VGND VPWR VPWR core_a_data_wdata_o[16] sky130_fd_sc_hd__clkbuf_2
Xoutput128 _201_/Y VGND VGND VPWR VPWR core_a_data_be_o[1] sky130_fd_sc_hd__clkbuf_2
XANTENNA__269__A0 input9/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput117 _188_/Y VGND VGND VPWR VPWR core_a_data_addr_o[0] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input108_A wb_data_wdata_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_173_ _173_/A VGND VGND VPWR VPWR _241_/B sky130_fd_sc_hd__inv_2
Xinput19 core_a_data_rdata_i[26] VGND VGND VPWR VPWR _278_/A0 sky130_fd_sc_hd__buf_1
X_242_ _244_/A _242_/B VGND VGND VPWR VPWR _242_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_input73_A wb_data_addr_i[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_156_ _162_/A _231_/B VGND VGND VPWR VPWR _156_/Y sky130_fd_sc_hd__nor2_1
X_225_ _228_/A _225_/B VGND VGND VPWR VPWR _225_/Y sky130_fd_sc_hd__nor2_4
X_087_ _087_/A VGND VGND VPWR VPWR _191_/B sky130_fd_sc_hd__inv_2
XFILLER_33_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input36_A core_b_data_rdata_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_208_ _283_/S VGND VGND VPWR VPWR _224_/A sky130_fd_sc_hd__buf_1
X_139_ _143_/A _221_/B VGND VGND VPWR VPWR _139_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xrepeater247 _281_/S VGND VGND VPWR VPWR _283_/S sky130_fd_sc_hd__buf_8
XFILLER_34_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__082__A _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__278__A1 _278_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput118 _189_/Y VGND VGND VPWR VPWR core_a_data_addr_o[1] sky130_fd_sc_hd__clkbuf_2
Xoutput129 _203_/Y VGND VGND VPWR VPWR core_a_data_be_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_172_ _181_/A VGND VGND VPWR VPWR _180_/A sky130_fd_sc_hd__buf_2
X_241_ _244_/A _241_/B VGND VGND VPWR VPWR _241_/Y sky130_fd_sc_hd__nor2_4
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input66_A core_b_data_rvalid_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_224_ _224_/A VGND VGND VPWR VPWR _228_/A sky130_fd_sc_hd__buf_2
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_086_ _088_/A _190_/B VGND VGND VPWR VPWR _086_/Y sky130_fd_sc_hd__nor2_1
X_155_ _155_/A VGND VGND VPWR VPWR _231_/B sky130_fd_sc_hd__inv_2
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__175__A _175_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__085__A _085_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input29_A core_a_data_rdata_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_207_ _207_/A _207_/B VGND VGND VPWR VPWR _207_/Y sky130_fd_sc_hd__nor2_2
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_138_ _138_/A VGND VGND VPWR VPWR _221_/B sky130_fd_sc_hd__inv_2
XFILLER_38_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output135_A _222_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input96_A wb_data_wdata_i[22] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__093__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input11_A core_a_data_rdata_i[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput119 _190_/Y VGND VGND VPWR VPWR core_a_data_addr_o[2] sky130_fd_sc_hd__clkbuf_2
XFILLER_5_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input3_A core_a_data_rdata_i[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__088__A _088_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_240_ _245_/A VGND VGND VPWR VPWR _244_/A sky130_fd_sc_hd__clkbuf_2
X_171_ _171_/A _239_/B VGND VGND VPWR VPWR _171_/Y sky130_fd_sc_hd__nor2_2
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input59_A core_b_data_rdata_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input113_A wb_data_wdata_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_223_ _223_/A _223_/B VGND VGND VPWR VPWR _223_/Y sky130_fd_sc_hd__nor2_4
XFILLER_15_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ _085_/A VGND VGND VPWR VPWR _190_/B sky130_fd_sc_hd__inv_2
X_154_ _181_/A VGND VGND VPWR VPWR _162_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_output165_A _082_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__191__A _191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_206_ _207_/A _206_/B VGND VGND VPWR VPWR _206_/Y sky130_fd_sc_hd__nor2_2
X_137_ _143_/A _220_/B VGND VGND VPWR VPWR _137_/Y sky130_fd_sc_hd__nor2_8
XFILLER_19_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__186__A _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input41_A core_b_data_rdata_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input89_A wb_data_wdata_i[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__194__A _196_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_170_ _170_/A VGND VGND VPWR VPWR _239_/B sky130_fd_sc_hd__inv_2
XFILLER_6_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output208_A _128_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__189__A _191_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input106_A wb_data_wdata_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_153_ _153_/A VGND VGND VPWR VPWR _181_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_222_ _223_/A _222_/B VGND VGND VPWR VPWR _222_/Y sky130_fd_sc_hd__nor2_4
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_084_ _088_/A _189_/B VGND VGND VPWR VPWR _084_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_input71_A wb_data_addr_i[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_205_ _250_/A _250_/B _251_/A VGND VGND VPWR VPWR _205_/X sky130_fd_sc_hd__and3_1
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_136_ _136_/A VGND VGND VPWR VPWR _220_/B sky130_fd_sc_hd__inv_2
XFILLER_7_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input34_A core_b_data_rdata_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_119_ _125_/A _210_/B VGND VGND VPWR VPWR _119_/Y sky130_fd_sc_hd__nor2_8
XFILLER_7_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output188_A _152_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ _083_/A VGND VGND VPWR VPWR _189_/B sky130_fd_sc_hd__inv_2
X_152_ _152_/A _228_/B VGND VGND VPWR VPWR _152_/Y sky130_fd_sc_hd__nor2_4
XFILLER_23_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_221_ _223_/A _221_/B VGND VGND VPWR VPWR _221_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input64_A core_b_data_rdata_i[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_204_ _207_/A _204_/B VGND VGND VPWR VPWR _204_/Y sky130_fd_sc_hd__nor2_4
X_135_ _144_/A VGND VGND VPWR VPWR _143_/A sky130_fd_sc_hd__buf_4
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input27_A core_a_data_rdata_i[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_118_ _118_/A VGND VGND VPWR VPWR _210_/B sky130_fd_sc_hd__inv_2
XFILLER_7_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output133_A _220_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input94_A wb_data_wdata_i[20] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_repeater246_A _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input1_A core_a_data_rdata_i[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__271__A0 _271_/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_220_ _223_/A _220_/B VGND VGND VPWR VPWR _220_/Y sky130_fd_sc_hd__nor2_4
X_151_ _151_/A VGND VGND VPWR VPWR _228_/B sky130_fd_sc_hd__inv_2
X_082_ _088_/A _188_/B VGND VGND VPWR VPWR _082_/Y sky130_fd_sc_hd__nor2_2
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_input57_A core_b_data_rdata_i[30] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input111_A wb_data_wdata_i[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_203_ _207_/A _203_/B VGND VGND VPWR VPWR _203_/Y sky130_fd_sc_hd__nor2_1
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_134_ _134_/A _218_/B VGND VGND VPWR VPWR _134_/Y sky130_fd_sc_hd__nor2_4
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_117_ _144_/A VGND VGND VPWR VPWR _125_/A sky130_fd_sc_hd__buf_6
XFILLER_7_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output126_A _199_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__253__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input87_A wb_data_wdata_i[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__102__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output243_A _260_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__280__A1 _280_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__271__A1 _271_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_150_ _152_/A _227_/B VGND VGND VPWR VPWR _150_/Y sky130_fd_sc_hd__nor2_4
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_081_ _081_/A VGND VGND VPWR VPWR _188_/B sky130_fd_sc_hd__inv_2
XFILLER_2_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__262__A1 _262_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_279_ _279_/A0 _279_/A1 _283_/S VGND VGND VPWR VPWR _279_/X sky130_fd_sc_hd__mux2_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__261__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__253__A1 _253_/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput240 _257_/X VGND VGND VPWR VPWR wb_data_rdata_o[5] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__200__A _201_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input104_A wb_data_wdata_i[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_133_ _133_/A VGND VGND VPWR VPWR _218_/B sky130_fd_sc_hd__inv_2
X_202_ _202_/A VGND VGND VPWR VPWR _207_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__256__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_116_ _153_/A VGND VGND VPWR VPWR _144_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA_output119_A _190_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input32_A core_a_data_rdata_i[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_output236_A _282_/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__264__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__203__A _207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__259__S _281_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_080_ _107_/A VGND VGND VPWR VPWR _088_/A sky130_fd_sc_hd__buf_2
XFILLER_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_278_ _278_/A0 _278_/A1 _283_/S VGND VGND VPWR VPWR _278_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput230 _277_/X VGND VGND VPWR VPWR wb_data_rdata_o[25] sky130_fd_sc_hd__clkbuf_2
Xoutput241 _258_/X VGND VGND VPWR VPWR wb_data_rdata_o[6] sky130_fd_sc_hd__clkbuf_2
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_132_ _134_/A _217_/B VGND VGND VPWR VPWR _132_/Y sky130_fd_sc_hd__nor2_2
X_201_ _201_/A _201_/B VGND VGND VPWR VPWR _201_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input62_A core_b_data_rdata_i[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output149_A _239_/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__272__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__211__A _213_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_115_ _115_/A _207_/B VGND VGND VPWR VPWR _115_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__121__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__267__S _284_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__206__A _207_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input25_A core_a_data_rdata_i[31] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XANTENNA__280__S _283_/S VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

