magic
tech sky130A
magscale 1 2
timestamp 1625057774
<< obsli1 >>
rect 1104 2159 238832 157777
<< obsm1 >>
rect 474 1844 239278 158500
<< metal2 >>
rect 938 159200 994 160000
rect 3238 159200 3294 160000
rect 5998 159200 6054 160000
rect 8298 159200 8354 160000
rect 10598 159200 10654 160000
rect 12898 159200 12954 160000
rect 15658 159200 15714 160000
rect 17958 159200 18014 160000
rect 20258 159200 20314 160000
rect 22558 159200 22614 160000
rect 24858 159200 24914 160000
rect 27618 159200 27674 160000
rect 29918 159200 29974 160000
rect 32218 159200 32274 160000
rect 34518 159200 34574 160000
rect 37278 159200 37334 160000
rect 39578 159200 39634 160000
rect 41878 159200 41934 160000
rect 44178 159200 44234 160000
rect 46938 159200 46994 160000
rect 49238 159200 49294 160000
rect 51538 159200 51594 160000
rect 53838 159200 53894 160000
rect 56598 159200 56654 160000
rect 58898 159200 58954 160000
rect 61198 159200 61254 160000
rect 63498 159200 63554 160000
rect 65798 159200 65854 160000
rect 68558 159200 68614 160000
rect 70858 159200 70914 160000
rect 73158 159200 73214 160000
rect 75458 159200 75514 160000
rect 78218 159200 78274 160000
rect 80518 159200 80574 160000
rect 82818 159200 82874 160000
rect 85118 159200 85174 160000
rect 87878 159200 87934 160000
rect 90178 159200 90234 160000
rect 92478 159200 92534 160000
rect 94778 159200 94834 160000
rect 97538 159200 97594 160000
rect 99838 159200 99894 160000
rect 102138 159200 102194 160000
rect 104438 159200 104494 160000
rect 107198 159200 107254 160000
rect 109498 159200 109554 160000
rect 111798 159200 111854 160000
rect 114098 159200 114154 160000
rect 116398 159200 116454 160000
rect 119158 159200 119214 160000
rect 121458 159200 121514 160000
rect 123758 159200 123814 160000
rect 126058 159200 126114 160000
rect 128818 159200 128874 160000
rect 131118 159200 131174 160000
rect 133418 159200 133474 160000
rect 135718 159200 135774 160000
rect 138478 159200 138534 160000
rect 140778 159200 140834 160000
rect 143078 159200 143134 160000
rect 145378 159200 145434 160000
rect 148138 159200 148194 160000
rect 150438 159200 150494 160000
rect 152738 159200 152794 160000
rect 155038 159200 155094 160000
rect 157338 159200 157394 160000
rect 160098 159200 160154 160000
rect 162398 159200 162454 160000
rect 164698 159200 164754 160000
rect 166998 159200 167054 160000
rect 169758 159200 169814 160000
rect 172058 159200 172114 160000
rect 174358 159200 174414 160000
rect 176658 159200 176714 160000
rect 179418 159200 179474 160000
rect 181718 159200 181774 160000
rect 184018 159200 184074 160000
rect 186318 159200 186374 160000
rect 189078 159200 189134 160000
rect 191378 159200 191434 160000
rect 193678 159200 193734 160000
rect 195978 159200 196034 160000
rect 198278 159200 198334 160000
rect 201038 159200 201094 160000
rect 203338 159200 203394 160000
rect 205638 159200 205694 160000
rect 207938 159200 207994 160000
rect 210698 159200 210754 160000
rect 212998 159200 213054 160000
rect 215298 159200 215354 160000
rect 217598 159200 217654 160000
rect 220358 159200 220414 160000
rect 222658 159200 222714 160000
rect 224958 159200 225014 160000
rect 227258 159200 227314 160000
rect 230018 159200 230074 160000
rect 232318 159200 232374 160000
rect 234618 159200 234674 160000
rect 236918 159200 236974 160000
rect 239218 159200 239274 160000
rect 478 0 534 800
rect 2778 0 2834 800
rect 5078 0 5134 800
rect 7378 0 7434 800
rect 9678 0 9734 800
rect 12438 0 12494 800
rect 14738 0 14794 800
rect 17038 0 17094 800
rect 19338 0 19394 800
rect 22098 0 22154 800
rect 24398 0 24454 800
rect 26698 0 26754 800
rect 28998 0 29054 800
rect 31758 0 31814 800
rect 34058 0 34114 800
rect 36358 0 36414 800
rect 38658 0 38714 800
rect 41418 0 41474 800
rect 43718 0 43774 800
rect 46018 0 46074 800
rect 48318 0 48374 800
rect 50618 0 50674 800
rect 53378 0 53434 800
rect 55678 0 55734 800
rect 57978 0 58034 800
rect 60278 0 60334 800
rect 63038 0 63094 800
rect 65338 0 65394 800
rect 67638 0 67694 800
rect 69938 0 69994 800
rect 72698 0 72754 800
rect 74998 0 75054 800
rect 77298 0 77354 800
rect 79598 0 79654 800
rect 82358 0 82414 800
rect 84658 0 84714 800
rect 86958 0 87014 800
rect 89258 0 89314 800
rect 91558 0 91614 800
rect 94318 0 94374 800
rect 96618 0 96674 800
rect 98918 0 98974 800
rect 101218 0 101274 800
rect 103978 0 104034 800
rect 106278 0 106334 800
rect 108578 0 108634 800
rect 110878 0 110934 800
rect 113638 0 113694 800
rect 115938 0 115994 800
rect 118238 0 118294 800
rect 120538 0 120594 800
rect 123298 0 123354 800
rect 125598 0 125654 800
rect 127898 0 127954 800
rect 130198 0 130254 800
rect 132498 0 132554 800
rect 135258 0 135314 800
rect 137558 0 137614 800
rect 139858 0 139914 800
rect 142158 0 142214 800
rect 144918 0 144974 800
rect 147218 0 147274 800
rect 149518 0 149574 800
rect 151818 0 151874 800
rect 154578 0 154634 800
rect 156878 0 156934 800
rect 159178 0 159234 800
rect 161478 0 161534 800
rect 164238 0 164294 800
rect 166538 0 166594 800
rect 168838 0 168894 800
rect 171138 0 171194 800
rect 173898 0 173954 800
rect 176198 0 176254 800
rect 178498 0 178554 800
rect 180798 0 180854 800
rect 183098 0 183154 800
rect 185858 0 185914 800
rect 188158 0 188214 800
rect 190458 0 190514 800
rect 192758 0 192814 800
rect 195518 0 195574 800
rect 197818 0 197874 800
rect 200118 0 200174 800
rect 202418 0 202474 800
rect 205178 0 205234 800
rect 207478 0 207534 800
rect 209778 0 209834 800
rect 212078 0 212134 800
rect 214838 0 214894 800
rect 217138 0 217194 800
rect 219438 0 219494 800
rect 221738 0 221794 800
rect 224038 0 224094 800
rect 226798 0 226854 800
rect 229098 0 229154 800
rect 231398 0 231454 800
rect 233698 0 233754 800
rect 236458 0 236514 800
rect 238758 0 238814 800
<< obsm2 >>
rect 480 159144 882 159200
rect 1050 159144 3182 159200
rect 3350 159144 5942 159200
rect 6110 159144 8242 159200
rect 8410 159144 10542 159200
rect 10710 159144 12842 159200
rect 13010 159144 15602 159200
rect 15770 159144 17902 159200
rect 18070 159144 20202 159200
rect 20370 159144 22502 159200
rect 22670 159144 24802 159200
rect 24970 159144 27562 159200
rect 27730 159144 29862 159200
rect 30030 159144 32162 159200
rect 32330 159144 34462 159200
rect 34630 159144 37222 159200
rect 37390 159144 39522 159200
rect 39690 159144 41822 159200
rect 41990 159144 44122 159200
rect 44290 159144 46882 159200
rect 47050 159144 49182 159200
rect 49350 159144 51482 159200
rect 51650 159144 53782 159200
rect 53950 159144 56542 159200
rect 56710 159144 58842 159200
rect 59010 159144 61142 159200
rect 61310 159144 63442 159200
rect 63610 159144 65742 159200
rect 65910 159144 68502 159200
rect 68670 159144 70802 159200
rect 70970 159144 73102 159200
rect 73270 159144 75402 159200
rect 75570 159144 78162 159200
rect 78330 159144 80462 159200
rect 80630 159144 82762 159200
rect 82930 159144 85062 159200
rect 85230 159144 87822 159200
rect 87990 159144 90122 159200
rect 90290 159144 92422 159200
rect 92590 159144 94722 159200
rect 94890 159144 97482 159200
rect 97650 159144 99782 159200
rect 99950 159144 102082 159200
rect 102250 159144 104382 159200
rect 104550 159144 107142 159200
rect 107310 159144 109442 159200
rect 109610 159144 111742 159200
rect 111910 159144 114042 159200
rect 114210 159144 116342 159200
rect 116510 159144 119102 159200
rect 119270 159144 121402 159200
rect 121570 159144 123702 159200
rect 123870 159144 126002 159200
rect 126170 159144 128762 159200
rect 128930 159144 131062 159200
rect 131230 159144 133362 159200
rect 133530 159144 135662 159200
rect 135830 159144 138422 159200
rect 138590 159144 140722 159200
rect 140890 159144 143022 159200
rect 143190 159144 145322 159200
rect 145490 159144 148082 159200
rect 148250 159144 150382 159200
rect 150550 159144 152682 159200
rect 152850 159144 154982 159200
rect 155150 159144 157282 159200
rect 157450 159144 160042 159200
rect 160210 159144 162342 159200
rect 162510 159144 164642 159200
rect 164810 159144 166942 159200
rect 167110 159144 169702 159200
rect 169870 159144 172002 159200
rect 172170 159144 174302 159200
rect 174470 159144 176602 159200
rect 176770 159144 179362 159200
rect 179530 159144 181662 159200
rect 181830 159144 183962 159200
rect 184130 159144 186262 159200
rect 186430 159144 189022 159200
rect 189190 159144 191322 159200
rect 191490 159144 193622 159200
rect 193790 159144 195922 159200
rect 196090 159144 198222 159200
rect 198390 159144 200982 159200
rect 201150 159144 203282 159200
rect 203450 159144 205582 159200
rect 205750 159144 207882 159200
rect 208050 159144 210642 159200
rect 210810 159144 212942 159200
rect 213110 159144 215242 159200
rect 215410 159144 217542 159200
rect 217710 159144 220302 159200
rect 220470 159144 222602 159200
rect 222770 159144 224902 159200
rect 225070 159144 227202 159200
rect 227370 159144 229962 159200
rect 230130 159144 232262 159200
rect 232430 159144 234562 159200
rect 234730 159144 236862 159200
rect 237030 159144 239162 159200
rect 480 856 239272 159144
rect 590 800 2722 856
rect 2890 800 5022 856
rect 5190 800 7322 856
rect 7490 800 9622 856
rect 9790 800 12382 856
rect 12550 800 14682 856
rect 14850 800 16982 856
rect 17150 800 19282 856
rect 19450 800 22042 856
rect 22210 800 24342 856
rect 24510 800 26642 856
rect 26810 800 28942 856
rect 29110 800 31702 856
rect 31870 800 34002 856
rect 34170 800 36302 856
rect 36470 800 38602 856
rect 38770 800 41362 856
rect 41530 800 43662 856
rect 43830 800 45962 856
rect 46130 800 48262 856
rect 48430 800 50562 856
rect 50730 800 53322 856
rect 53490 800 55622 856
rect 55790 800 57922 856
rect 58090 800 60222 856
rect 60390 800 62982 856
rect 63150 800 65282 856
rect 65450 800 67582 856
rect 67750 800 69882 856
rect 70050 800 72642 856
rect 72810 800 74942 856
rect 75110 800 77242 856
rect 77410 800 79542 856
rect 79710 800 82302 856
rect 82470 800 84602 856
rect 84770 800 86902 856
rect 87070 800 89202 856
rect 89370 800 91502 856
rect 91670 800 94262 856
rect 94430 800 96562 856
rect 96730 800 98862 856
rect 99030 800 101162 856
rect 101330 800 103922 856
rect 104090 800 106222 856
rect 106390 800 108522 856
rect 108690 800 110822 856
rect 110990 800 113582 856
rect 113750 800 115882 856
rect 116050 800 118182 856
rect 118350 800 120482 856
rect 120650 800 123242 856
rect 123410 800 125542 856
rect 125710 800 127842 856
rect 128010 800 130142 856
rect 130310 800 132442 856
rect 132610 800 135202 856
rect 135370 800 137502 856
rect 137670 800 139802 856
rect 139970 800 142102 856
rect 142270 800 144862 856
rect 145030 800 147162 856
rect 147330 800 149462 856
rect 149630 800 151762 856
rect 151930 800 154522 856
rect 154690 800 156822 856
rect 156990 800 159122 856
rect 159290 800 161422 856
rect 161590 800 164182 856
rect 164350 800 166482 856
rect 166650 800 168782 856
rect 168950 800 171082 856
rect 171250 800 173842 856
rect 174010 800 176142 856
rect 176310 800 178442 856
rect 178610 800 180742 856
rect 180910 800 183042 856
rect 183210 800 185802 856
rect 185970 800 188102 856
rect 188270 800 190402 856
rect 190570 800 192702 856
rect 192870 800 195462 856
rect 195630 800 197762 856
rect 197930 800 200062 856
rect 200230 800 202362 856
rect 202530 800 205122 856
rect 205290 800 207422 856
rect 207590 800 209722 856
rect 209890 800 212022 856
rect 212190 800 214782 856
rect 214950 800 217082 856
rect 217250 800 219382 856
rect 219550 800 221682 856
rect 221850 800 223982 856
rect 224150 800 226742 856
rect 226910 800 229042 856
rect 229210 800 231342 856
rect 231510 800 233642 856
rect 233810 800 236402 856
rect 236570 800 238702 856
rect 238870 800 239272 856
<< metal3 >>
rect 0 157088 800 157208
rect 239200 155728 240000 155848
rect 0 153688 800 153808
rect 239200 152328 240000 152448
rect 0 149608 800 149728
rect 239200 148928 240000 149048
rect 0 146208 800 146328
rect 239200 145528 240000 145648
rect 0 142808 800 142928
rect 239200 141448 240000 141568
rect 0 139408 800 139528
rect 239200 138048 240000 138168
rect 0 135328 800 135448
rect 239200 134648 240000 134768
rect 0 131928 800 132048
rect 239200 131248 240000 131368
rect 0 128528 800 128648
rect 239200 127168 240000 127288
rect 0 125128 800 125248
rect 239200 123768 240000 123888
rect 0 121728 800 121848
rect 239200 120368 240000 120488
rect 0 117648 800 117768
rect 239200 116968 240000 117088
rect 0 114248 800 114368
rect 239200 112888 240000 113008
rect 0 110848 800 110968
rect 239200 109488 240000 109608
rect 0 107448 800 107568
rect 239200 106088 240000 106208
rect 0 103368 800 103488
rect 239200 102688 240000 102808
rect 0 99968 800 100088
rect 239200 98608 240000 98728
rect 0 96568 800 96688
rect 239200 95208 240000 95328
rect 0 93168 800 93288
rect 239200 91808 240000 91928
rect 0 89088 800 89208
rect 239200 88408 240000 88528
rect 0 85688 800 85808
rect 239200 85008 240000 85128
rect 0 82288 800 82408
rect 239200 80928 240000 81048
rect 0 78888 800 79008
rect 239200 77528 240000 77648
rect 0 74808 800 74928
rect 239200 74128 240000 74248
rect 0 71408 800 71528
rect 239200 70728 240000 70848
rect 0 68008 800 68128
rect 239200 66648 240000 66768
rect 0 64608 800 64728
rect 239200 63248 240000 63368
rect 0 61208 800 61328
rect 239200 59848 240000 59968
rect 0 57128 800 57248
rect 239200 56448 240000 56568
rect 0 53728 800 53848
rect 239200 52368 240000 52488
rect 0 50328 800 50448
rect 239200 48968 240000 49088
rect 0 46928 800 47048
rect 239200 45568 240000 45688
rect 0 42848 800 42968
rect 239200 42168 240000 42288
rect 0 39448 800 39568
rect 239200 38088 240000 38208
rect 0 36048 800 36168
rect 239200 34688 240000 34808
rect 0 32648 800 32768
rect 239200 31288 240000 31408
rect 0 28568 800 28688
rect 239200 27888 240000 28008
rect 0 25168 800 25288
rect 239200 24488 240000 24608
rect 0 21768 800 21888
rect 239200 20408 240000 20528
rect 0 18368 800 18488
rect 239200 17008 240000 17128
rect 0 14288 800 14408
rect 239200 13608 240000 13728
rect 0 10888 800 11008
rect 239200 10208 240000 10328
rect 0 7488 800 7608
rect 239200 6128 240000 6248
rect 0 4088 800 4208
rect 239200 2728 240000 2848
<< obsm3 >>
rect 800 157288 239200 157793
rect 880 157008 239200 157288
rect 800 155928 239200 157008
rect 800 155648 239120 155928
rect 800 153888 239200 155648
rect 880 153608 239200 153888
rect 800 152528 239200 153608
rect 800 152248 239120 152528
rect 800 149808 239200 152248
rect 880 149528 239200 149808
rect 800 149128 239200 149528
rect 800 148848 239120 149128
rect 800 146408 239200 148848
rect 880 146128 239200 146408
rect 800 145728 239200 146128
rect 800 145448 239120 145728
rect 800 143008 239200 145448
rect 880 142728 239200 143008
rect 800 141648 239200 142728
rect 800 141368 239120 141648
rect 800 139608 239200 141368
rect 880 139328 239200 139608
rect 800 138248 239200 139328
rect 800 137968 239120 138248
rect 800 135528 239200 137968
rect 880 135248 239200 135528
rect 800 134848 239200 135248
rect 800 134568 239120 134848
rect 800 132128 239200 134568
rect 880 131848 239200 132128
rect 800 131448 239200 131848
rect 800 131168 239120 131448
rect 800 128728 239200 131168
rect 880 128448 239200 128728
rect 800 127368 239200 128448
rect 800 127088 239120 127368
rect 800 125328 239200 127088
rect 880 125048 239200 125328
rect 800 123968 239200 125048
rect 800 123688 239120 123968
rect 800 121928 239200 123688
rect 880 121648 239200 121928
rect 800 120568 239200 121648
rect 800 120288 239120 120568
rect 800 117848 239200 120288
rect 880 117568 239200 117848
rect 800 117168 239200 117568
rect 800 116888 239120 117168
rect 800 114448 239200 116888
rect 880 114168 239200 114448
rect 800 113088 239200 114168
rect 800 112808 239120 113088
rect 800 111048 239200 112808
rect 880 110768 239200 111048
rect 800 109688 239200 110768
rect 800 109408 239120 109688
rect 800 107648 239200 109408
rect 880 107368 239200 107648
rect 800 106288 239200 107368
rect 800 106008 239120 106288
rect 800 103568 239200 106008
rect 880 103288 239200 103568
rect 800 102888 239200 103288
rect 800 102608 239120 102888
rect 800 100168 239200 102608
rect 880 99888 239200 100168
rect 800 98808 239200 99888
rect 800 98528 239120 98808
rect 800 96768 239200 98528
rect 880 96488 239200 96768
rect 800 95408 239200 96488
rect 800 95128 239120 95408
rect 800 93368 239200 95128
rect 880 93088 239200 93368
rect 800 92008 239200 93088
rect 800 91728 239120 92008
rect 800 89288 239200 91728
rect 880 89008 239200 89288
rect 800 88608 239200 89008
rect 800 88328 239120 88608
rect 800 85888 239200 88328
rect 880 85608 239200 85888
rect 800 85208 239200 85608
rect 800 84928 239120 85208
rect 800 82488 239200 84928
rect 880 82208 239200 82488
rect 800 81128 239200 82208
rect 800 80848 239120 81128
rect 800 79088 239200 80848
rect 880 78808 239200 79088
rect 800 77728 239200 78808
rect 800 77448 239120 77728
rect 800 75008 239200 77448
rect 880 74728 239200 75008
rect 800 74328 239200 74728
rect 800 74048 239120 74328
rect 800 71608 239200 74048
rect 880 71328 239200 71608
rect 800 70928 239200 71328
rect 800 70648 239120 70928
rect 800 68208 239200 70648
rect 880 67928 239200 68208
rect 800 66848 239200 67928
rect 800 66568 239120 66848
rect 800 64808 239200 66568
rect 880 64528 239200 64808
rect 800 63448 239200 64528
rect 800 63168 239120 63448
rect 800 61408 239200 63168
rect 880 61128 239200 61408
rect 800 60048 239200 61128
rect 800 59768 239120 60048
rect 800 57328 239200 59768
rect 880 57048 239200 57328
rect 800 56648 239200 57048
rect 800 56368 239120 56648
rect 800 53928 239200 56368
rect 880 53648 239200 53928
rect 800 52568 239200 53648
rect 800 52288 239120 52568
rect 800 50528 239200 52288
rect 880 50248 239200 50528
rect 800 49168 239200 50248
rect 800 48888 239120 49168
rect 800 47128 239200 48888
rect 880 46848 239200 47128
rect 800 45768 239200 46848
rect 800 45488 239120 45768
rect 800 43048 239200 45488
rect 880 42768 239200 43048
rect 800 42368 239200 42768
rect 800 42088 239120 42368
rect 800 39648 239200 42088
rect 880 39368 239200 39648
rect 800 38288 239200 39368
rect 800 38008 239120 38288
rect 800 36248 239200 38008
rect 880 35968 239200 36248
rect 800 34888 239200 35968
rect 800 34608 239120 34888
rect 800 32848 239200 34608
rect 880 32568 239200 32848
rect 800 31488 239200 32568
rect 800 31208 239120 31488
rect 800 28768 239200 31208
rect 880 28488 239200 28768
rect 800 28088 239200 28488
rect 800 27808 239120 28088
rect 800 25368 239200 27808
rect 880 25088 239200 25368
rect 800 24688 239200 25088
rect 800 24408 239120 24688
rect 800 21968 239200 24408
rect 880 21688 239200 21968
rect 800 20608 239200 21688
rect 800 20328 239120 20608
rect 800 18568 239200 20328
rect 880 18288 239200 18568
rect 800 17208 239200 18288
rect 800 16928 239120 17208
rect 800 14488 239200 16928
rect 880 14208 239200 14488
rect 800 13808 239200 14208
rect 800 13528 239120 13808
rect 800 11088 239200 13528
rect 880 10808 239200 11088
rect 800 10408 239200 10808
rect 800 10128 239120 10408
rect 800 7688 239200 10128
rect 880 7408 239200 7688
rect 800 6328 239200 7408
rect 800 6048 239120 6328
rect 800 4288 239200 6048
rect 880 4008 239200 4288
rect 800 2928 239200 4008
rect 800 2648 239120 2928
rect 800 2143 239200 2648
<< metal4 >>
rect 4208 2128 4528 157808
rect 9208 2128 9528 157808
rect 14208 95452 14528 157808
rect 19208 95452 19528 157808
rect 24208 95452 24528 157808
rect 29208 95452 29528 157808
rect 34208 95452 34528 157808
rect 39208 95452 39528 157808
rect 44208 95452 44528 157808
rect 49208 95452 49528 157808
rect 54208 95452 54528 157808
rect 59208 95452 59528 157808
rect 64208 95452 64528 157808
rect 69208 95452 69528 157808
rect 74208 95452 74528 157808
rect 79208 95452 79528 157808
rect 84208 95452 84528 157808
rect 89208 95452 89528 157808
rect 94208 95452 94528 157808
rect 99208 95452 99528 157808
rect 104208 95452 104528 157808
rect 109208 95452 109528 157808
rect 14208 2128 14528 14048
rect 19208 2128 19528 14048
rect 24208 2128 24528 14048
rect 29208 2128 29528 14048
rect 34208 2128 34528 14048
rect 39208 2128 39528 14048
rect 44208 2128 44528 14048
rect 49208 2128 49528 14048
rect 54208 2128 54528 14048
rect 59208 2128 59528 14048
rect 64208 2128 64528 14048
rect 69208 2128 69528 14048
rect 74208 2128 74528 14048
rect 79208 2128 79528 14048
rect 84208 2128 84528 14048
rect 89208 2128 89528 14048
rect 94208 2128 94528 14048
rect 99208 2128 99528 14048
rect 104208 2128 104528 14048
rect 109208 2128 109528 14048
rect 114208 2128 114528 157808
rect 119208 2128 119528 157808
rect 124208 2128 124528 157808
rect 129208 2128 129528 157808
rect 134208 2128 134528 157808
rect 139208 2128 139528 157808
rect 144208 2128 144528 157808
rect 149208 2128 149528 157808
rect 154208 2128 154528 157808
rect 159208 2128 159528 157808
rect 164208 2128 164528 157808
rect 169208 2128 169528 157808
rect 174208 2128 174528 157808
rect 179208 2128 179528 157808
rect 184208 2128 184528 157808
rect 189208 2128 189528 157808
rect 194208 2128 194528 157808
rect 199208 2128 199528 157808
rect 204208 2128 204528 157808
rect 209208 2128 209528 157808
rect 214208 2128 214528 157808
rect 219208 2128 219528 157808
rect 224208 2128 224528 157808
rect 229208 2128 229528 157808
rect 234208 2128 234528 157808
<< obsm4 >>
rect 1814 2483 4128 141813
rect 4608 2483 9128 141813
rect 9608 95372 14128 141813
rect 14608 95372 19128 141813
rect 19608 95372 24128 141813
rect 24608 95372 29128 141813
rect 29608 95372 34128 141813
rect 34608 95372 39128 141813
rect 39608 95372 44128 141813
rect 44608 95372 49128 141813
rect 49608 95372 54128 141813
rect 54608 95372 59128 141813
rect 59608 95372 64128 141813
rect 64608 95372 69128 141813
rect 69608 95372 74128 141813
rect 74608 95372 79128 141813
rect 79608 95372 84128 141813
rect 84608 95372 89128 141813
rect 89608 95372 94128 141813
rect 94608 95372 99128 141813
rect 99608 95372 104128 141813
rect 104608 95372 109128 141813
rect 109608 95372 114128 141813
rect 9608 14128 114128 95372
rect 9608 2483 14128 14128
rect 14608 2483 19128 14128
rect 19608 2483 24128 14128
rect 24608 2483 29128 14128
rect 29608 2483 34128 14128
rect 34608 2483 39128 14128
rect 39608 2483 44128 14128
rect 44608 2483 49128 14128
rect 49608 2483 54128 14128
rect 54608 2483 59128 14128
rect 59608 2483 64128 14128
rect 64608 2483 69128 14128
rect 69608 2483 74128 14128
rect 74608 2483 79128 14128
rect 79608 2483 84128 14128
rect 84608 2483 89128 14128
rect 89608 2483 94128 14128
rect 94608 2483 99128 14128
rect 99608 2483 104128 14128
rect 104608 2483 109128 14128
rect 109608 2483 114128 14128
rect 114608 2483 119128 141813
rect 119608 2483 124128 141813
rect 124608 2483 129128 141813
rect 129608 2483 134128 141813
rect 134608 2483 139128 141813
rect 139608 2483 144128 141813
rect 144608 2483 149128 141813
rect 149608 2483 154128 141813
rect 154608 2483 159128 141813
rect 159608 2483 164128 141813
rect 164608 2483 169128 141813
rect 169608 2483 174128 141813
rect 174608 2483 179128 141813
rect 179608 2483 184128 141813
rect 184608 2483 189128 141813
rect 189608 2483 194128 141813
rect 194608 2483 199128 141813
rect 199608 2483 204128 141813
rect 204608 2483 209128 141813
rect 209608 2483 214128 141813
rect 214608 2483 215037 141813
<< metal5 >>
rect 1104 143160 238832 143480
rect 1104 127842 238832 128162
rect 1104 112524 238832 112844
rect 1104 97206 238832 97526
rect 1104 81888 238832 82208
rect 1104 66570 238832 66890
rect 1104 51252 238832 51572
rect 1104 35934 238832 36254
rect 1104 20616 238832 20936
rect 1104 5298 238832 5618
<< obsm5 >>
rect 1772 97846 167140 98420
rect 1772 82528 167140 96886
rect 1772 67210 167140 81568
rect 1772 51892 167140 66250
rect 1772 36574 167140 50932
rect 1772 21256 167140 35614
rect 1772 15140 167140 20296
<< labels >>
rlabel metal3 s 0 25168 800 25288 6 clk_i
port 1 nsew signal input
rlabel metal3 s 239200 109488 240000 109608 6 debug_req_i
port 2 nsew signal input
rlabel metal2 s 234618 159200 234674 160000 6 eFPGA_delay_o[0]
port 3 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 eFPGA_delay_o[1]
port 4 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 eFPGA_delay_o[2]
port 5 nsew signal output
rlabel metal2 s 181718 159200 181774 160000 6 eFPGA_delay_o[3]
port 6 nsew signal output
rlabel metal2 s 109498 159200 109554 160000 6 eFPGA_en_o
port 7 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 eFPGA_fpga_done_i
port 8 nsew signal input
rlabel metal3 s 239200 102688 240000 102808 6 eFPGA_operand_a_o[0]
port 9 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 eFPGA_operand_a_o[10]
port 10 nsew signal output
rlabel metal2 s 27618 159200 27674 160000 6 eFPGA_operand_a_o[11]
port 11 nsew signal output
rlabel metal2 s 202418 0 202474 800 6 eFPGA_operand_a_o[12]
port 12 nsew signal output
rlabel metal2 s 63038 0 63094 800 6 eFPGA_operand_a_o[13]
port 13 nsew signal output
rlabel metal2 s 127898 0 127954 800 6 eFPGA_operand_a_o[14]
port 14 nsew signal output
rlabel metal2 s 230018 159200 230074 160000 6 eFPGA_operand_a_o[15]
port 15 nsew signal output
rlabel metal3 s 239200 42168 240000 42288 6 eFPGA_operand_a_o[16]
port 16 nsew signal output
rlabel metal2 s 207938 159200 207994 160000 6 eFPGA_operand_a_o[17]
port 17 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 eFPGA_operand_a_o[18]
port 18 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 eFPGA_operand_a_o[19]
port 19 nsew signal output
rlabel metal2 s 46938 159200 46994 160000 6 eFPGA_operand_a_o[1]
port 20 nsew signal output
rlabel metal3 s 0 57128 800 57248 6 eFPGA_operand_a_o[20]
port 21 nsew signal output
rlabel metal3 s 239200 88408 240000 88528 6 eFPGA_operand_a_o[21]
port 22 nsew signal output
rlabel metal2 s 226798 0 226854 800 6 eFPGA_operand_a_o[22]
port 23 nsew signal output
rlabel metal2 s 233698 0 233754 800 6 eFPGA_operand_a_o[23]
port 24 nsew signal output
rlabel metal2 s 15658 159200 15714 160000 6 eFPGA_operand_a_o[24]
port 25 nsew signal output
rlabel metal2 s 91558 0 91614 800 6 eFPGA_operand_a_o[25]
port 26 nsew signal output
rlabel metal3 s 239200 127168 240000 127288 6 eFPGA_operand_a_o[26]
port 27 nsew signal output
rlabel metal3 s 239200 120368 240000 120488 6 eFPGA_operand_a_o[27]
port 28 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 eFPGA_operand_a_o[28]
port 29 nsew signal output
rlabel metal2 s 176658 159200 176714 160000 6 eFPGA_operand_a_o[29]
port 30 nsew signal output
rlabel metal3 s 239200 6128 240000 6248 6 eFPGA_operand_a_o[2]
port 31 nsew signal output
rlabel metal2 s 173898 0 173954 800 6 eFPGA_operand_a_o[30]
port 32 nsew signal output
rlabel metal2 s 157338 159200 157394 160000 6 eFPGA_operand_a_o[31]
port 33 nsew signal output
rlabel metal2 s 197818 0 197874 800 6 eFPGA_operand_a_o[3]
port 34 nsew signal output
rlabel metal2 s 224958 159200 225014 160000 6 eFPGA_operand_a_o[4]
port 35 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 eFPGA_operand_a_o[5]
port 36 nsew signal output
rlabel metal3 s 0 32648 800 32768 6 eFPGA_operand_a_o[6]
port 37 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 eFPGA_operand_a_o[7]
port 38 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 eFPGA_operand_a_o[8]
port 39 nsew signal output
rlabel metal2 s 128818 159200 128874 160000 6 eFPGA_operand_a_o[9]
port 40 nsew signal output
rlabel metal3 s 239200 134648 240000 134768 6 eFPGA_operand_b_o[0]
port 41 nsew signal output
rlabel metal3 s 239200 141448 240000 141568 6 eFPGA_operand_b_o[10]
port 42 nsew signal output
rlabel metal2 s 145378 159200 145434 160000 6 eFPGA_operand_b_o[11]
port 43 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 eFPGA_operand_b_o[12]
port 44 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 eFPGA_operand_b_o[13]
port 45 nsew signal output
rlabel metal2 s 162398 159200 162454 160000 6 eFPGA_operand_b_o[14]
port 46 nsew signal output
rlabel metal2 s 107198 159200 107254 160000 6 eFPGA_operand_b_o[15]
port 47 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 eFPGA_operand_b_o[16]
port 48 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 eFPGA_operand_b_o[17]
port 49 nsew signal output
rlabel metal2 s 192758 0 192814 800 6 eFPGA_operand_b_o[18]
port 50 nsew signal output
rlabel metal2 s 68558 159200 68614 160000 6 eFPGA_operand_b_o[19]
port 51 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 eFPGA_operand_b_o[1]
port 52 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 eFPGA_operand_b_o[20]
port 53 nsew signal output
rlabel metal3 s 239200 52368 240000 52488 6 eFPGA_operand_b_o[21]
port 54 nsew signal output
rlabel metal2 s 169758 159200 169814 160000 6 eFPGA_operand_b_o[22]
port 55 nsew signal output
rlabel metal2 s 131118 159200 131174 160000 6 eFPGA_operand_b_o[23]
port 56 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 eFPGA_operand_b_o[24]
port 57 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 eFPGA_operand_b_o[25]
port 58 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 eFPGA_operand_b_o[26]
port 59 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 eFPGA_operand_b_o[27]
port 60 nsew signal output
rlabel metal2 s 58898 159200 58954 160000 6 eFPGA_operand_b_o[28]
port 61 nsew signal output
rlabel metal2 s 144918 0 144974 800 6 eFPGA_operand_b_o[29]
port 62 nsew signal output
rlabel metal3 s 239200 77528 240000 77648 6 eFPGA_operand_b_o[2]
port 63 nsew signal output
rlabel metal3 s 239200 10208 240000 10328 6 eFPGA_operand_b_o[30]
port 64 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 eFPGA_operand_b_o[31]
port 65 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 eFPGA_operand_b_o[3]
port 66 nsew signal output
rlabel metal3 s 0 157088 800 157208 6 eFPGA_operand_b_o[4]
port 67 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 eFPGA_operand_b_o[5]
port 68 nsew signal output
rlabel metal2 s 166998 159200 167054 160000 6 eFPGA_operand_b_o[6]
port 69 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 eFPGA_operand_b_o[7]
port 70 nsew signal output
rlabel metal2 s 193678 159200 193734 160000 6 eFPGA_operand_b_o[8]
port 71 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 eFPGA_operand_b_o[9]
port 72 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 eFPGA_operator_o[0]
port 73 nsew signal output
rlabel metal3 s 239200 74128 240000 74248 6 eFPGA_operator_o[1]
port 74 nsew signal output
rlabel metal2 s 82818 159200 82874 160000 6 eFPGA_result_a_i[0]
port 75 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 eFPGA_result_a_i[10]
port 76 nsew signal input
rlabel metal2 s 164698 159200 164754 160000 6 eFPGA_result_a_i[11]
port 77 nsew signal input
rlabel metal2 s 17958 159200 18014 160000 6 eFPGA_result_a_i[12]
port 78 nsew signal input
rlabel metal3 s 239200 138048 240000 138168 6 eFPGA_result_a_i[13]
port 79 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 eFPGA_result_a_i[14]
port 80 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 eFPGA_result_a_i[15]
port 81 nsew signal input
rlabel metal2 s 191378 159200 191434 160000 6 eFPGA_result_a_i[16]
port 82 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 eFPGA_result_a_i[17]
port 83 nsew signal input
rlabel metal2 s 80518 159200 80574 160000 6 eFPGA_result_a_i[18]
port 84 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 eFPGA_result_a_i[19]
port 85 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 eFPGA_result_a_i[1]
port 86 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 eFPGA_result_a_i[20]
port 87 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 eFPGA_result_a_i[21]
port 88 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 eFPGA_result_a_i[22]
port 89 nsew signal input
rlabel metal3 s 0 139408 800 139528 6 eFPGA_result_a_i[23]
port 90 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 eFPGA_result_a_i[24]
port 91 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 eFPGA_result_a_i[25]
port 92 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 eFPGA_result_a_i[26]
port 93 nsew signal input
rlabel metal2 s 8298 159200 8354 160000 6 eFPGA_result_a_i[27]
port 94 nsew signal input
rlabel metal2 s 135718 159200 135774 160000 6 eFPGA_result_a_i[28]
port 95 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 eFPGA_result_a_i[29]
port 96 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 eFPGA_result_a_i[2]
port 97 nsew signal input
rlabel metal3 s 239200 112888 240000 113008 6 eFPGA_result_a_i[30]
port 98 nsew signal input
rlabel metal2 s 133418 159200 133474 160000 6 eFPGA_result_a_i[31]
port 99 nsew signal input
rlabel metal2 s 195978 159200 196034 160000 6 eFPGA_result_a_i[3]
port 100 nsew signal input
rlabel metal2 s 121458 159200 121514 160000 6 eFPGA_result_a_i[4]
port 101 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 eFPGA_result_a_i[5]
port 102 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 eFPGA_result_a_i[6]
port 103 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 eFPGA_result_a_i[7]
port 104 nsew signal input
rlabel metal2 s 220358 159200 220414 160000 6 eFPGA_result_a_i[8]
port 105 nsew signal input
rlabel metal2 s 123758 159200 123814 160000 6 eFPGA_result_a_i[9]
port 106 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 eFPGA_result_b_i[0]
port 107 nsew signal input
rlabel metal3 s 239200 48968 240000 49088 6 eFPGA_result_b_i[10]
port 108 nsew signal input
rlabel metal2 s 205638 159200 205694 160000 6 eFPGA_result_b_i[11]
port 109 nsew signal input
rlabel metal3 s 239200 38088 240000 38208 6 eFPGA_result_b_i[12]
port 110 nsew signal input
rlabel metal2 s 119158 159200 119214 160000 6 eFPGA_result_b_i[13]
port 111 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 eFPGA_result_b_i[14]
port 112 nsew signal input
rlabel metal2 s 39578 159200 39634 160000 6 eFPGA_result_b_i[15]
port 113 nsew signal input
rlabel metal3 s 239200 145528 240000 145648 6 eFPGA_result_b_i[16]
port 114 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 eFPGA_result_b_i[17]
port 115 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 eFPGA_result_b_i[18]
port 116 nsew signal input
rlabel metal2 s 189078 159200 189134 160000 6 eFPGA_result_b_i[19]
port 117 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 eFPGA_result_b_i[1]
port 118 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 eFPGA_result_b_i[20]
port 119 nsew signal input
rlabel metal2 s 152738 159200 152794 160000 6 eFPGA_result_b_i[21]
port 120 nsew signal input
rlabel metal2 s 32218 159200 32274 160000 6 eFPGA_result_b_i[22]
port 121 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 eFPGA_result_b_i[23]
port 122 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 eFPGA_result_b_i[24]
port 123 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 eFPGA_result_b_i[25]
port 124 nsew signal input
rlabel metal2 s 140778 159200 140834 160000 6 eFPGA_result_b_i[26]
port 125 nsew signal input
rlabel metal2 s 24858 159200 24914 160000 6 eFPGA_result_b_i[27]
port 126 nsew signal input
rlabel metal3 s 239200 116968 240000 117088 6 eFPGA_result_b_i[28]
port 127 nsew signal input
rlabel metal3 s 239200 123768 240000 123888 6 eFPGA_result_b_i[29]
port 128 nsew signal input
rlabel metal2 s 73158 159200 73214 160000 6 eFPGA_result_b_i[2]
port 129 nsew signal input
rlabel metal2 s 41878 159200 41934 160000 6 eFPGA_result_b_i[30]
port 130 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 eFPGA_result_b_i[31]
port 131 nsew signal input
rlabel metal2 s 222658 159200 222714 160000 6 eFPGA_result_b_i[3]
port 132 nsew signal input
rlabel metal3 s 239200 131248 240000 131368 6 eFPGA_result_b_i[4]
port 133 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 eFPGA_result_b_i[5]
port 134 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 eFPGA_result_b_i[6]
port 135 nsew signal input
rlabel metal2 s 212078 0 212134 800 6 eFPGA_result_b_i[7]
port 136 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 eFPGA_result_b_i[8]
port 137 nsew signal input
rlabel metal2 s 116398 159200 116454 160000 6 eFPGA_result_b_i[9]
port 138 nsew signal input
rlabel metal2 s 148138 159200 148194 160000 6 eFPGA_result_c_i[0]
port 139 nsew signal input
rlabel metal2 s 186318 159200 186374 160000 6 eFPGA_result_c_i[10]
port 140 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 eFPGA_result_c_i[11]
port 141 nsew signal input
rlabel metal3 s 0 99968 800 100088 6 eFPGA_result_c_i[12]
port 142 nsew signal input
rlabel metal2 s 180798 0 180854 800 6 eFPGA_result_c_i[13]
port 143 nsew signal input
rlabel metal2 s 160098 159200 160154 160000 6 eFPGA_result_c_i[14]
port 144 nsew signal input
rlabel metal2 s 231398 0 231454 800 6 eFPGA_result_c_i[15]
port 145 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 eFPGA_result_c_i[16]
port 146 nsew signal input
rlabel metal2 s 938 159200 994 160000 6 eFPGA_result_c_i[17]
port 147 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 eFPGA_result_c_i[18]
port 148 nsew signal input
rlabel metal2 s 166538 0 166594 800 6 eFPGA_result_c_i[19]
port 149 nsew signal input
rlabel metal2 s 185858 0 185914 800 6 eFPGA_result_c_i[1]
port 150 nsew signal input
rlabel metal2 s 221738 0 221794 800 6 eFPGA_result_c_i[20]
port 151 nsew signal input
rlabel metal2 s 238758 0 238814 800 6 eFPGA_result_c_i[21]
port 152 nsew signal input
rlabel metal2 s 478 0 534 800 6 eFPGA_result_c_i[22]
port 153 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 eFPGA_result_c_i[23]
port 154 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 eFPGA_result_c_i[24]
port 155 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 eFPGA_result_c_i[25]
port 156 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 eFPGA_result_c_i[26]
port 157 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 eFPGA_result_c_i[27]
port 158 nsew signal input
rlabel metal2 s 94778 159200 94834 160000 6 eFPGA_result_c_i[28]
port 159 nsew signal input
rlabel metal2 s 61198 159200 61254 160000 6 eFPGA_result_c_i[29]
port 160 nsew signal input
rlabel metal2 s 154578 0 154634 800 6 eFPGA_result_c_i[2]
port 161 nsew signal input
rlabel metal2 s 217598 159200 217654 160000 6 eFPGA_result_c_i[30]
port 162 nsew signal input
rlabel metal2 s 5998 159200 6054 160000 6 eFPGA_result_c_i[31]
port 163 nsew signal input
rlabel metal2 s 53838 159200 53894 160000 6 eFPGA_result_c_i[3]
port 164 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 eFPGA_result_c_i[4]
port 165 nsew signal input
rlabel metal3 s 239200 34688 240000 34808 6 eFPGA_result_c_i[5]
port 166 nsew signal input
rlabel metal2 s 150438 159200 150494 160000 6 eFPGA_result_c_i[6]
port 167 nsew signal input
rlabel metal2 s 236918 159200 236974 160000 6 eFPGA_result_c_i[7]
port 168 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 eFPGA_result_c_i[8]
port 169 nsew signal input
rlabel metal3 s 239200 24488 240000 24608 6 eFPGA_result_c_i[9]
port 170 nsew signal input
rlabel metal2 s 99838 159200 99894 160000 6 eFPGA_write_strobe_o
port 171 nsew signal output
rlabel metal2 s 200118 0 200174 800 6 ext_data_addr_i[0]
port 172 nsew signal input
rlabel metal3 s 239200 155728 240000 155848 6 ext_data_addr_i[10]
port 173 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 ext_data_addr_i[11]
port 174 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 ext_data_addr_i[12]
port 175 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 ext_data_addr_i[13]
port 176 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 ext_data_addr_i[14]
port 177 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 ext_data_addr_i[15]
port 178 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 ext_data_addr_i[16]
port 179 nsew signal input
rlabel metal2 s 102138 159200 102194 160000 6 ext_data_addr_i[17]
port 180 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 ext_data_addr_i[18]
port 181 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 ext_data_addr_i[19]
port 182 nsew signal input
rlabel metal3 s 239200 56448 240000 56568 6 ext_data_addr_i[1]
port 183 nsew signal input
rlabel metal2 s 49238 159200 49294 160000 6 ext_data_addr_i[20]
port 184 nsew signal input
rlabel metal3 s 239200 95208 240000 95328 6 ext_data_addr_i[21]
port 185 nsew signal input
rlabel metal2 s 92478 159200 92534 160000 6 ext_data_addr_i[22]
port 186 nsew signal input
rlabel metal3 s 239200 2728 240000 2848 6 ext_data_addr_i[23]
port 187 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 ext_data_addr_i[24]
port 188 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 ext_data_addr_i[25]
port 189 nsew signal input
rlabel metal3 s 239200 152328 240000 152448 6 ext_data_addr_i[26]
port 190 nsew signal input
rlabel metal2 s 75458 159200 75514 160000 6 ext_data_addr_i[27]
port 191 nsew signal input
rlabel metal2 s 179418 159200 179474 160000 6 ext_data_addr_i[28]
port 192 nsew signal input
rlabel metal2 s 198278 159200 198334 160000 6 ext_data_addr_i[29]
port 193 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 ext_data_addr_i[2]
port 194 nsew signal input
rlabel metal2 s 104438 159200 104494 160000 6 ext_data_addr_i[30]
port 195 nsew signal input
rlabel metal2 s 126058 159200 126114 160000 6 ext_data_addr_i[31]
port 196 nsew signal input
rlabel metal2 s 85118 159200 85174 160000 6 ext_data_addr_i[3]
port 197 nsew signal input
rlabel metal2 s 227258 159200 227314 160000 6 ext_data_addr_i[4]
port 198 nsew signal input
rlabel metal2 s 224038 0 224094 800 6 ext_data_addr_i[5]
port 199 nsew signal input
rlabel metal2 s 70858 159200 70914 160000 6 ext_data_addr_i[6]
port 200 nsew signal input
rlabel metal2 s 97538 159200 97594 160000 6 ext_data_addr_i[7]
port 201 nsew signal input
rlabel metal2 s 12898 159200 12954 160000 6 ext_data_addr_i[8]
port 202 nsew signal input
rlabel metal2 s 10598 159200 10654 160000 6 ext_data_addr_i[9]
port 203 nsew signal input
rlabel metal2 s 56598 159200 56654 160000 6 ext_data_be_i[0]
port 204 nsew signal input
rlabel metal2 s 219438 0 219494 800 6 ext_data_be_i[1]
port 205 nsew signal input
rlabel metal2 s 44178 159200 44234 160000 6 ext_data_be_i[2]
port 206 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 ext_data_be_i[3]
port 207 nsew signal input
rlabel metal2 s 20258 159200 20314 160000 6 ext_data_rdata_o[0]
port 208 nsew signal output
rlabel metal2 s 190458 0 190514 800 6 ext_data_rdata_o[10]
port 209 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 ext_data_rdata_o[11]
port 210 nsew signal output
rlabel metal3 s 239200 80928 240000 81048 6 ext_data_rdata_o[12]
port 211 nsew signal output
rlabel metal2 s 138478 159200 138534 160000 6 ext_data_rdata_o[13]
port 212 nsew signal output
rlabel metal3 s 239200 91808 240000 91928 6 ext_data_rdata_o[14]
port 213 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 ext_data_rdata_o[15]
port 214 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 ext_data_rdata_o[16]
port 215 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 ext_data_rdata_o[17]
port 216 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 ext_data_rdata_o[18]
port 217 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 ext_data_rdata_o[19]
port 218 nsew signal output
rlabel metal3 s 239200 66648 240000 66768 6 ext_data_rdata_o[1]
port 219 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 ext_data_rdata_o[20]
port 220 nsew signal output
rlabel metal2 s 209778 0 209834 800 6 ext_data_rdata_o[21]
port 221 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 ext_data_rdata_o[22]
port 222 nsew signal output
rlabel metal3 s 239200 13608 240000 13728 6 ext_data_rdata_o[23]
port 223 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 ext_data_rdata_o[24]
port 224 nsew signal output
rlabel metal2 s 201038 159200 201094 160000 6 ext_data_rdata_o[25]
port 225 nsew signal output
rlabel metal2 s 22558 159200 22614 160000 6 ext_data_rdata_o[26]
port 226 nsew signal output
rlabel metal2 s 65798 159200 65854 160000 6 ext_data_rdata_o[27]
port 227 nsew signal output
rlabel metal2 s 161478 0 161534 800 6 ext_data_rdata_o[28]
port 228 nsew signal output
rlabel metal2 s 239218 159200 239274 160000 6 ext_data_rdata_o[29]
port 229 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 ext_data_rdata_o[2]
port 230 nsew signal output
rlabel metal2 s 205178 0 205234 800 6 ext_data_rdata_o[30]
port 231 nsew signal output
rlabel metal2 s 51538 159200 51594 160000 6 ext_data_rdata_o[31]
port 232 nsew signal output
rlabel metal2 s 229098 0 229154 800 6 ext_data_rdata_o[3]
port 233 nsew signal output
rlabel metal3 s 239200 70728 240000 70848 6 ext_data_rdata_o[4]
port 234 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 ext_data_rdata_o[5]
port 235 nsew signal output
rlabel metal3 s 239200 17008 240000 17128 6 ext_data_rdata_o[6]
port 236 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 ext_data_rdata_o[7]
port 237 nsew signal output
rlabel metal2 s 184018 159200 184074 160000 6 ext_data_rdata_o[8]
port 238 nsew signal output
rlabel metal2 s 174358 159200 174414 160000 6 ext_data_rdata_o[9]
port 239 nsew signal output
rlabel metal2 s 34518 159200 34574 160000 6 ext_data_req_i
port 240 nsew signal input
rlabel metal2 s 90178 159200 90234 160000 6 ext_data_rvalid_o
port 241 nsew signal output
rlabel metal2 s 63498 159200 63554 160000 6 ext_data_wdata_i[0]
port 242 nsew signal input
rlabel metal3 s 239200 148928 240000 149048 6 ext_data_wdata_i[10]
port 243 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 ext_data_wdata_i[11]
port 244 nsew signal input
rlabel metal3 s 239200 45568 240000 45688 6 ext_data_wdata_i[12]
port 245 nsew signal input
rlabel metal3 s 239200 20408 240000 20528 6 ext_data_wdata_i[13]
port 246 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 ext_data_wdata_i[14]
port 247 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 ext_data_wdata_i[15]
port 248 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 ext_data_wdata_i[16]
port 249 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 ext_data_wdata_i[17]
port 250 nsew signal input
rlabel metal3 s 239200 63248 240000 63368 6 ext_data_wdata_i[18]
port 251 nsew signal input
rlabel metal2 s 210698 159200 210754 160000 6 ext_data_wdata_i[19]
port 252 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 ext_data_wdata_i[1]
port 253 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 ext_data_wdata_i[20]
port 254 nsew signal input
rlabel metal3 s 239200 98608 240000 98728 6 ext_data_wdata_i[21]
port 255 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 ext_data_wdata_i[22]
port 256 nsew signal input
rlabel metal2 s 29918 159200 29974 160000 6 ext_data_wdata_i[23]
port 257 nsew signal input
rlabel metal2 s 232318 159200 232374 160000 6 ext_data_wdata_i[24]
port 258 nsew signal input
rlabel metal2 s 172058 159200 172114 160000 6 ext_data_wdata_i[25]
port 259 nsew signal input
rlabel metal2 s 143078 159200 143134 160000 6 ext_data_wdata_i[26]
port 260 nsew signal input
rlabel metal2 s 188158 0 188214 800 6 ext_data_wdata_i[27]
port 261 nsew signal input
rlabel metal3 s 239200 59848 240000 59968 6 ext_data_wdata_i[28]
port 262 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 ext_data_wdata_i[29]
port 263 nsew signal input
rlabel metal3 s 239200 31288 240000 31408 6 ext_data_wdata_i[2]
port 264 nsew signal input
rlabel metal2 s 215298 159200 215354 160000 6 ext_data_wdata_i[30]
port 265 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 ext_data_wdata_i[31]
port 266 nsew signal input
rlabel metal2 s 78218 159200 78274 160000 6 ext_data_wdata_i[3]
port 267 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 ext_data_wdata_i[4]
port 268 nsew signal input
rlabel metal3 s 239200 106088 240000 106208 6 ext_data_wdata_i[5]
port 269 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 ext_data_wdata_i[6]
port 270 nsew signal input
rlabel metal2 s 37278 159200 37334 160000 6 ext_data_wdata_i[7]
port 271 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 ext_data_wdata_i[8]
port 272 nsew signal input
rlabel metal2 s 87878 159200 87934 160000 6 ext_data_wdata_i[9]
port 273 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 ext_data_we_i
port 274 nsew signal input
rlabel metal2 s 207478 0 207534 800 6 fetch_enable_i
port 275 nsew signal input
rlabel metal2 s 111798 159200 111854 160000 6 irq_ack_o
port 276 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 irq_i
port 277 nsew signal input
rlabel metal2 s 203338 159200 203394 160000 6 irq_id_i[0]
port 278 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 irq_id_i[1]
port 279 nsew signal input
rlabel metal2 s 114098 159200 114154 160000 6 irq_id_i[2]
port 280 nsew signal input
rlabel metal3 s 239200 27888 240000 28008 6 irq_id_i[3]
port 281 nsew signal input
rlabel metal2 s 214838 0 214894 800 6 irq_id_i[4]
port 282 nsew signal input
rlabel metal2 s 155038 159200 155094 160000 6 irq_id_o[0]
port 283 nsew signal output
rlabel metal2 s 236458 0 236514 800 6 irq_id_o[1]
port 284 nsew signal output
rlabel metal2 s 212998 159200 213054 160000 6 irq_id_o[2]
port 285 nsew signal output
rlabel metal2 s 3238 159200 3294 160000 6 irq_id_o[3]
port 286 nsew signal output
rlabel metal3 s 239200 85008 240000 85128 6 irq_id_o[4]
port 287 nsew signal output
rlabel metal2 s 115938 0 115994 800 6 reset
port 288 nsew signal input
rlabel metal4 s 234208 2128 234528 157808 6 VPWR
port 289 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 157808 6 VPWR
port 290 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 157808 6 VPWR
port 291 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 157808 6 VPWR
port 292 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 157808 6 VPWR
port 293 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 157808 6 VPWR
port 294 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 157808 6 VPWR
port 295 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 157808 6 VPWR
port 296 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 157808 6 VPWR
port 297 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 157808 6 VPWR
port 298 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 157808 6 VPWR
port 299 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 157808 6 VPWR
port 300 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 157808 6 VPWR
port 301 nsew power bidirectional
rlabel metal4 s 104208 95452 104528 157808 6 VPWR
port 302 nsew power bidirectional
rlabel metal4 s 94208 95452 94528 157808 6 VPWR
port 303 nsew power bidirectional
rlabel metal4 s 84208 95452 84528 157808 6 VPWR
port 304 nsew power bidirectional
rlabel metal4 s 74208 95452 74528 157808 6 VPWR
port 305 nsew power bidirectional
rlabel metal4 s 64208 95452 64528 157808 6 VPWR
port 306 nsew power bidirectional
rlabel metal4 s 54208 95452 54528 157808 6 VPWR
port 307 nsew power bidirectional
rlabel metal4 s 44208 95452 44528 157808 6 VPWR
port 308 nsew power bidirectional
rlabel metal4 s 34208 95452 34528 157808 6 VPWR
port 309 nsew power bidirectional
rlabel metal4 s 24208 95452 24528 157808 6 VPWR
port 310 nsew power bidirectional
rlabel metal4 s 14208 95452 14528 157808 6 VPWR
port 311 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 157808 6 VPWR
port 312 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 14048 6 VPWR
port 313 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 14048 6 VPWR
port 314 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 14048 6 VPWR
port 315 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 14048 6 VPWR
port 316 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 14048 6 VPWR
port 317 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 14048 6 VPWR
port 318 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 14048 6 VPWR
port 319 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 14048 6 VPWR
port 320 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 14048 6 VPWR
port 321 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 14048 6 VPWR
port 322 nsew power bidirectional
rlabel metal5 s 1104 127842 238832 128162 6 VPWR
port 323 nsew power bidirectional
rlabel metal5 s 1104 97206 238832 97526 6 VPWR
port 324 nsew power bidirectional
rlabel metal5 s 1104 66570 238832 66890 6 VPWR
port 325 nsew power bidirectional
rlabel metal5 s 1104 35934 238832 36254 6 VPWR
port 326 nsew power bidirectional
rlabel metal5 s 1104 5298 238832 5618 6 VPWR
port 327 nsew power bidirectional
rlabel metal4 s 229208 2128 229528 157808 6 VGND
port 328 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 157808 6 VGND
port 329 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 157808 6 VGND
port 330 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 157808 6 VGND
port 331 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 157808 6 VGND
port 332 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 157808 6 VGND
port 333 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 157808 6 VGND
port 334 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 157808 6 VGND
port 335 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 157808 6 VGND
port 336 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 157808 6 VGND
port 337 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 157808 6 VGND
port 338 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 157808 6 VGND
port 339 nsew ground bidirectional
rlabel metal4 s 109208 95452 109528 157808 6 VGND
port 340 nsew ground bidirectional
rlabel metal4 s 99208 95452 99528 157808 6 VGND
port 341 nsew ground bidirectional
rlabel metal4 s 89208 95452 89528 157808 6 VGND
port 342 nsew ground bidirectional
rlabel metal4 s 79208 95452 79528 157808 6 VGND
port 343 nsew ground bidirectional
rlabel metal4 s 69208 95452 69528 157808 6 VGND
port 344 nsew ground bidirectional
rlabel metal4 s 59208 95452 59528 157808 6 VGND
port 345 nsew ground bidirectional
rlabel metal4 s 49208 95452 49528 157808 6 VGND
port 346 nsew ground bidirectional
rlabel metal4 s 39208 95452 39528 157808 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 29208 95452 29528 157808 6 VGND
port 348 nsew ground bidirectional
rlabel metal4 s 19208 95452 19528 157808 6 VGND
port 349 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 157808 6 VGND
port 350 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 14048 6 VGND
port 351 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 14048 6 VGND
port 352 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 14048 6 VGND
port 353 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 14048 6 VGND
port 354 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 14048 6 VGND
port 355 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 14048 6 VGND
port 356 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 14048 6 VGND
port 357 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 14048 6 VGND
port 358 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 14048 6 VGND
port 359 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 14048 6 VGND
port 360 nsew ground bidirectional
rlabel metal5 s 1104 143160 238832 143480 6 VGND
port 361 nsew ground bidirectional
rlabel metal5 s 1104 112524 238832 112844 6 VGND
port 362 nsew ground bidirectional
rlabel metal5 s 1104 81888 238832 82208 6 VGND
port 363 nsew ground bidirectional
rlabel metal5 s 1104 51252 238832 51572 6 VGND
port 364 nsew ground bidirectional
rlabel metal5 s 1104 20616 238832 20936 6 VGND
port 365 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 240000 160000
string LEFview TRUE
string GDS_FILE /project/openlane/core_sram/runs/core_sram/results/magic/core_sram.gds
string GDS_END 67747250
string GDS_START 10596454
<< end >>

