magic
tech sky130A
magscale 1 2
timestamp 1624390257
<< locali >>
rect 29285 26231 29319 26401
rect 19993 22967 20027 23137
rect 50813 20927 50847 21029
rect 29929 4471 29963 4641
rect 40877 4063 40911 4233
rect 48329 2363 48363 2533
rect 48329 1751 48363 1921
<< viali >>
rect 3157 27625 3191 27659
rect 8033 27625 8067 27659
rect 13829 27625 13863 27659
rect 22017 27625 22051 27659
rect 29929 27625 29963 27659
rect 37381 27625 37415 27659
rect 43177 27625 43211 27659
rect 47041 27625 47075 27659
rect 50537 27625 50571 27659
rect 56517 27625 56551 27659
rect 2605 27557 2639 27591
rect 5549 27557 5583 27591
rect 5733 27557 5767 27591
rect 7941 27557 7975 27591
rect 8585 27557 8619 27591
rect 9689 27557 9723 27591
rect 10609 27557 10643 27591
rect 11989 27557 12023 27591
rect 12449 27557 12483 27591
rect 14933 27557 14967 27591
rect 15945 27557 15979 27591
rect 16497 27557 16531 27591
rect 16681 27557 16715 27591
rect 19349 27557 19383 27591
rect 20637 27557 20671 27591
rect 23949 27557 23983 27591
rect 25605 27557 25639 27591
rect 25789 27557 25823 27591
rect 28089 27557 28123 27591
rect 28641 27557 28675 27591
rect 32229 27557 32263 27591
rect 33977 27557 34011 27591
rect 34161 27557 34195 27591
rect 36277 27557 36311 27591
rect 37544 27557 37578 27591
rect 37749 27557 37783 27591
rect 39497 27557 39531 27591
rect 42441 27557 42475 27591
rect 42625 27557 42659 27591
rect 44281 27557 44315 27591
rect 45293 27557 45327 27591
rect 46029 27557 46063 27591
rect 47133 27557 47167 27591
rect 47685 27557 47719 27591
rect 48513 27557 48547 27591
rect 49617 27557 49651 27591
rect 51273 27557 51307 27591
rect 52469 27557 52503 27591
rect 53573 27557 53607 27591
rect 54953 27557 54987 27591
rect 55689 27557 55723 27591
rect 58081 27557 58115 27591
rect 1409 27489 1443 27523
rect 2421 27489 2455 27523
rect 3249 27489 3283 27523
rect 4629 27489 4663 27523
rect 4721 27489 4755 27523
rect 7113 27489 7147 27523
rect 9873 27489 9907 27523
rect 10793 27489 10827 27523
rect 12633 27489 12667 27523
rect 13921 27489 13955 27523
rect 15117 27489 15151 27523
rect 15761 27489 15795 27523
rect 17693 27489 17727 27523
rect 17877 27489 17911 27523
rect 18613 27489 18647 27523
rect 19165 27489 19199 27523
rect 20269 27489 20303 27523
rect 20453 27489 20487 27523
rect 21281 27489 21315 27523
rect 21833 27489 21867 27523
rect 22569 27489 22603 27523
rect 23305 27489 23339 27523
rect 24133 27489 24167 27523
rect 26801 27489 26835 27523
rect 26893 27489 26927 27523
rect 27077 27489 27111 27523
rect 29837 27489 29871 27523
rect 31585 27489 31619 27523
rect 32413 27489 32447 27523
rect 34989 27489 35023 27523
rect 36461 27489 36495 27523
rect 39313 27489 39347 27523
rect 40325 27489 40359 27523
rect 41613 27489 41647 27523
rect 43269 27489 43303 27523
rect 44465 27489 44499 27523
rect 45109 27489 45143 27523
rect 45845 27489 45879 27523
rect 49801 27489 49835 27523
rect 50445 27489 50479 27523
rect 55137 27489 55171 27523
rect 55873 27489 55907 27523
rect 56609 27489 56643 27523
rect 4905 27421 4939 27455
rect 17601 27421 17635 27455
rect 21097 27421 21131 27455
rect 34253 27421 34287 27455
rect 39589 27421 39623 27455
rect 6929 27353 6963 27387
rect 13277 27353 13311 27387
rect 31769 27353 31803 27387
rect 39037 27353 39071 27387
rect 40141 27353 40175 27387
rect 1593 27285 1627 27319
rect 4261 27285 4295 27319
rect 18429 27285 18463 27319
rect 23397 27285 23431 27319
rect 28733 27285 28767 27319
rect 30573 27285 30607 27319
rect 33701 27285 33735 27319
rect 34897 27285 34931 27319
rect 37565 27285 37599 27319
rect 41797 27285 41831 27319
rect 48421 27285 48455 27319
rect 51181 27285 51215 27319
rect 52377 27285 52411 27319
rect 53481 27285 53515 27319
rect 57805 27285 57839 27319
rect 23305 27081 23339 27115
rect 48697 27081 48731 27115
rect 52101 27081 52135 27115
rect 53757 27081 53791 27115
rect 2145 27013 2179 27047
rect 3065 27013 3099 27047
rect 4261 27013 4295 27047
rect 8677 27013 8711 27047
rect 16313 27013 16347 27047
rect 17969 27013 18003 27047
rect 22569 27013 22603 27047
rect 26893 27013 26927 27047
rect 29009 27013 29043 27047
rect 29561 27013 29595 27047
rect 30849 27013 30883 27047
rect 38485 27013 38519 27047
rect 40417 27013 40451 27047
rect 41889 27013 41923 27047
rect 44097 27013 44131 27047
rect 44649 27013 44683 27047
rect 45385 27013 45419 27047
rect 47869 27013 47903 27047
rect 49709 27013 49743 27047
rect 50169 27013 50203 27047
rect 51089 27013 51123 27047
rect 56149 27013 56183 27047
rect 57437 27013 57471 27047
rect 4721 26945 4755 26979
rect 6837 26945 6871 26979
rect 9321 26945 9355 26979
rect 19073 26945 19107 26979
rect 26065 26945 26099 26979
rect 30021 26945 30055 26979
rect 33517 26945 33551 26979
rect 33609 26945 33643 26979
rect 35725 26945 35759 26979
rect 39589 26945 39623 26979
rect 55045 26945 55079 26979
rect 1501 26877 1535 26911
rect 2881 26877 2915 26911
rect 3525 26877 3559 26911
rect 5549 26877 5583 26911
rect 7021 26877 7055 26911
rect 7573 26877 7607 26911
rect 8493 26877 8527 26911
rect 9413 26877 9447 26911
rect 10609 26877 10643 26911
rect 11161 26877 11195 26911
rect 12081 26877 12115 26911
rect 12909 26877 12943 26911
rect 13553 26877 13587 26911
rect 14289 26877 14323 26911
rect 14933 26877 14967 26911
rect 15761 26877 15795 26911
rect 16405 26877 16439 26911
rect 17417 26877 17451 26911
rect 20545 26877 20579 26911
rect 21097 26877 21131 26911
rect 23305 26877 23339 26911
rect 23489 26877 23523 26911
rect 24133 26877 24167 26911
rect 24869 26877 24903 26911
rect 25329 26877 25363 26911
rect 25973 26877 26007 26911
rect 26157 26877 26191 26911
rect 27813 26877 27847 26911
rect 28089 26877 28123 26911
rect 30113 26877 30147 26911
rect 31953 26877 31987 26911
rect 34437 26877 34471 26911
rect 34713 26877 34747 26911
rect 35541 26877 35575 26911
rect 35817 26877 35851 26911
rect 36553 26877 36587 26911
rect 36737 26877 36771 26911
rect 37381 26877 37415 26911
rect 38301 26877 38335 26911
rect 39865 26877 39899 26911
rect 41153 26877 41187 26911
rect 43177 26877 43211 26911
rect 45569 26877 45603 26911
rect 46029 26877 46063 26911
rect 50353 26877 50387 26911
rect 54401 26877 54435 26911
rect 55689 26877 55723 26911
rect 57253 26877 57287 26911
rect 58081 26877 58115 26911
rect 1685 26809 1719 26843
rect 2329 26809 2363 26843
rect 4813 26809 4847 26843
rect 9505 26809 9539 26843
rect 17509 26809 17543 26843
rect 17693 26809 17727 26843
rect 21557 26809 21591 26843
rect 22753 26809 22787 26843
rect 26709 26809 26743 26843
rect 28181 26809 28215 26843
rect 28825 26809 28859 26843
rect 30021 26809 30055 26843
rect 31033 26809 31067 26843
rect 33425 26809 33459 26843
rect 40601 26809 40635 26843
rect 42073 26809 42107 26843
rect 44833 26809 44867 26843
rect 47685 26809 47719 26843
rect 49525 26809 49559 26843
rect 51273 26809 51307 26843
rect 56333 26809 56367 26843
rect 57897 26809 57931 26843
rect 4721 26741 4755 26775
rect 5365 26741 5399 26775
rect 7757 26741 7791 26775
rect 9873 26741 9907 26775
rect 11069 26741 11103 26775
rect 12265 26741 12299 26775
rect 13093 26741 13127 26775
rect 14473 26741 14507 26775
rect 15577 26741 15611 26775
rect 19257 26741 19291 26775
rect 19349 26741 19383 26775
rect 19717 26741 19751 26775
rect 21005 26741 21039 26775
rect 23949 26741 23983 26775
rect 25513 26741 25547 26775
rect 31769 26741 31803 26775
rect 33057 26741 33091 26775
rect 34529 26741 34563 26775
rect 36737 26741 36771 26775
rect 41337 26741 41371 26775
rect 55505 26741 55539 26775
rect 1501 26537 1535 26571
rect 5181 26537 5215 26571
rect 5733 26537 5767 26571
rect 7389 26537 7423 26571
rect 8033 26537 8067 26571
rect 8585 26537 8619 26571
rect 10333 26537 10367 26571
rect 11713 26537 11747 26571
rect 12357 26537 12391 26571
rect 15853 26537 15887 26571
rect 17049 26537 17083 26571
rect 17693 26537 17727 26571
rect 23765 26537 23799 26571
rect 29469 26537 29503 26571
rect 32045 26537 32079 26571
rect 34161 26537 34195 26571
rect 35817 26537 35851 26571
rect 36369 26537 36403 26571
rect 41613 26537 41647 26571
rect 51549 26537 51583 26571
rect 54677 26537 54711 26571
rect 55781 26537 55815 26571
rect 1593 26469 1627 26503
rect 2973 26469 3007 26503
rect 4261 26469 4295 26503
rect 4445 26469 4479 26503
rect 9505 26469 9539 26503
rect 9689 26469 9723 26503
rect 11805 26469 11839 26503
rect 20269 26469 20303 26503
rect 21189 26469 21223 26503
rect 21373 26469 21407 26503
rect 27077 26469 27111 26503
rect 27629 26469 27663 26503
rect 33149 26469 33183 26503
rect 33333 26469 33367 26503
rect 38761 26469 38795 26503
rect 38853 26469 38887 26503
rect 55137 26469 55171 26503
rect 56701 26469 56735 26503
rect 58173 26469 58207 26503
rect 2329 26401 2363 26435
rect 10241 26401 10275 26435
rect 12541 26401 12575 26435
rect 13001 26401 13035 26435
rect 16957 26401 16991 26435
rect 17141 26401 17175 26435
rect 17693 26401 17727 26435
rect 17969 26401 18003 26435
rect 18889 26401 18923 26435
rect 19625 26401 19659 26435
rect 20453 26401 20487 26435
rect 22293 26401 22327 26435
rect 25881 26401 25915 26435
rect 26525 26401 26559 26435
rect 27169 26401 27203 26435
rect 27813 26401 27847 26435
rect 29285 26401 29319 26435
rect 29537 26401 29571 26435
rect 30665 26401 30699 26435
rect 31125 26401 31159 26435
rect 33977 26401 34011 26435
rect 34621 26401 34655 26435
rect 35725 26401 35759 26435
rect 36553 26401 36587 26435
rect 37381 26401 37415 26435
rect 37565 26401 37599 26435
rect 39589 26401 39623 26435
rect 41153 26401 41187 26435
rect 56885 26401 56919 26435
rect 57989 26401 58023 26435
rect 11713 26333 11747 26367
rect 2513 26265 2547 26299
rect 16497 26265 16531 26299
rect 26341 26265 26375 26299
rect 38669 26333 38703 26367
rect 37657 26265 37691 26299
rect 39405 26265 39439 26299
rect 49433 26265 49467 26299
rect 6377 26197 6411 26231
rect 11253 26197 11287 26231
rect 13553 26197 13587 26231
rect 15301 26197 15335 26231
rect 19073 26197 19107 26231
rect 22385 26197 22419 26231
rect 23213 26197 23247 26231
rect 25329 26197 25363 26231
rect 28365 26197 28399 26231
rect 29285 26197 29319 26231
rect 30481 26197 30515 26231
rect 32597 26197 32631 26231
rect 34713 26197 34747 26231
rect 38301 26197 38335 26231
rect 40969 26197 41003 26231
rect 42349 26197 42383 26231
rect 44465 26197 44499 26231
rect 45845 26197 45879 26231
rect 49985 26197 50019 26231
rect 2605 25993 2639 26027
rect 3433 25993 3467 26027
rect 33977 25993 34011 26027
rect 34437 25993 34471 26027
rect 36645 25993 36679 26027
rect 37197 25993 37231 26027
rect 38485 25993 38519 26027
rect 39221 25993 39255 26027
rect 40325 25993 40359 26027
rect 40969 25993 41003 26027
rect 41521 25993 41555 26027
rect 57253 25993 57287 26027
rect 5181 25925 5215 25959
rect 8769 25925 8803 25959
rect 9321 25925 9355 25959
rect 11069 25925 11103 25959
rect 11805 25925 11839 25959
rect 17509 25925 17543 25959
rect 18337 25925 18371 25959
rect 18889 25925 18923 25959
rect 34989 25925 35023 25959
rect 38669 25925 38703 25959
rect 55045 25925 55079 25959
rect 56701 25925 56735 25959
rect 1409 25857 1443 25891
rect 10517 25857 10551 25891
rect 17049 25857 17083 25891
rect 20085 25857 20119 25891
rect 55505 25857 55539 25891
rect 56149 25857 56183 25891
rect 57713 25857 57747 25891
rect 1593 25789 1627 25823
rect 5641 25789 5675 25823
rect 9787 25789 9821 25823
rect 9965 25789 9999 25823
rect 17693 25789 17727 25823
rect 19441 25789 19475 25823
rect 19533 25789 19567 25823
rect 21189 25789 21223 25823
rect 23673 25789 23707 25823
rect 26341 25789 26375 25823
rect 26801 25789 26835 25823
rect 29377 25789 29411 25823
rect 32781 25789 32815 25823
rect 33333 25789 33367 25823
rect 35173 25789 35207 25823
rect 35633 25789 35667 25823
rect 37197 25789 37231 25823
rect 37381 25789 37415 25823
rect 39865 25789 39899 25823
rect 38301 25721 38335 25755
rect 38517 25721 38551 25755
rect 57805 25721 57839 25755
rect 9873 25653 9907 25687
rect 26617 25653 26651 25687
rect 57713 25653 57747 25687
rect 2789 25449 2823 25483
rect 9965 25449 9999 25483
rect 16957 25449 16991 25483
rect 17785 25449 17819 25483
rect 34253 25449 34287 25483
rect 35633 25449 35667 25483
rect 37657 25449 37691 25483
rect 39681 25449 39715 25483
rect 57437 25449 57471 25483
rect 57989 25381 58023 25415
rect 58173 25381 58207 25415
rect 1593 25313 1627 25347
rect 18797 25313 18831 25347
rect 38209 25313 38243 25347
rect 38393 25313 38427 25347
rect 39025 25313 39059 25347
rect 39221 25313 39255 25347
rect 40601 25313 40635 25347
rect 56793 25313 56827 25347
rect 57253 25313 57287 25347
rect 33517 25245 33551 25279
rect 39129 25245 39163 25279
rect 1409 25177 1443 25211
rect 2237 25177 2271 25211
rect 36185 25177 36219 25211
rect 38485 25177 38519 25211
rect 36921 25109 36955 25143
rect 55689 25109 55723 25143
rect 1501 24905 1535 24939
rect 1961 24905 1995 24939
rect 34437 24905 34471 24939
rect 56425 24905 56459 24939
rect 56977 24905 57011 24939
rect 38025 24837 38059 24871
rect 39129 24837 39163 24871
rect 39681 24837 39715 24871
rect 38577 24769 38611 24803
rect 40141 24769 40175 24803
rect 23581 24701 23615 24735
rect 29009 24701 29043 24735
rect 57529 24701 57563 24735
rect 58173 24701 58207 24735
rect 23489 24565 23523 24599
rect 28917 24565 28951 24599
rect 36737 24565 36771 24599
rect 37289 24565 37323 24599
rect 57989 24565 58023 24599
rect 39037 24361 39071 24395
rect 56885 24361 56919 24395
rect 22661 24225 22695 24259
rect 22845 24225 22879 24259
rect 28181 24225 28215 24259
rect 28365 24225 28399 24259
rect 37749 24225 37783 24259
rect 38301 24225 38335 24259
rect 39129 24225 39163 24259
rect 39773 24225 39807 24259
rect 57529 24225 57563 24259
rect 58173 24225 58207 24259
rect 38485 24157 38519 24191
rect 39681 24157 39715 24191
rect 22569 24089 22603 24123
rect 28365 24089 28399 24123
rect 40693 24021 40727 24055
rect 57989 24021 58023 24055
rect 1501 23817 1535 23851
rect 22569 23817 22603 23851
rect 39221 23817 39255 23851
rect 37013 23749 37047 23783
rect 22569 23613 22603 23647
rect 22753 23613 22787 23647
rect 25789 23613 25823 23647
rect 25973 23613 26007 23647
rect 28089 23613 28123 23647
rect 28549 23613 28583 23647
rect 57529 23613 57563 23647
rect 58173 23613 58207 23647
rect 1593 23545 1627 23579
rect 26157 23545 26191 23579
rect 36829 23545 36863 23579
rect 2145 23477 2179 23511
rect 28273 23477 28307 23511
rect 57989 23477 58023 23511
rect 27445 23205 27479 23239
rect 27629 23205 27663 23239
rect 1409 23137 1443 23171
rect 1593 23137 1627 23171
rect 5089 23137 5123 23171
rect 19993 23137 20027 23171
rect 20637 23137 20671 23171
rect 20729 23137 20763 23171
rect 21557 23137 21591 23171
rect 21833 23137 21867 23171
rect 4905 23069 4939 23103
rect 2237 23001 2271 23035
rect 21557 23001 21591 23035
rect 19993 22933 20027 22967
rect 20085 22933 20119 22967
rect 4169 22729 4203 22763
rect 34897 22729 34931 22763
rect 36461 22729 36495 22763
rect 21189 22525 21223 22559
rect 21465 22525 21499 22559
rect 26433 22525 26467 22559
rect 35449 22525 35483 22559
rect 35541 22525 35575 22559
rect 36461 22525 36495 22559
rect 36645 22525 36679 22559
rect 57529 22525 57563 22559
rect 58173 22525 58207 22559
rect 1409 22457 1443 22491
rect 1593 22457 1627 22491
rect 2237 22457 2271 22491
rect 21097 22457 21131 22491
rect 26525 22389 26559 22423
rect 57989 22389 58023 22423
rect 27353 22185 27387 22219
rect 27261 22049 27295 22083
rect 27445 22049 27479 22083
rect 36277 22049 36311 22083
rect 36921 22049 36955 22083
rect 57989 22049 58023 22083
rect 36461 21913 36495 21947
rect 37105 21913 37139 21947
rect 57345 21913 57379 21947
rect 58173 21913 58207 21947
rect 19809 21641 19843 21675
rect 20453 21641 20487 21675
rect 29469 21641 29503 21675
rect 31401 21641 31435 21675
rect 36737 21573 36771 21607
rect 19809 21437 19843 21471
rect 19993 21437 20027 21471
rect 20453 21437 20487 21471
rect 20637 21437 20671 21471
rect 28733 21437 28767 21471
rect 31217 21437 31251 21471
rect 31401 21437 31435 21471
rect 35909 21437 35943 21471
rect 36829 21437 36863 21471
rect 36921 21437 36955 21471
rect 38301 21437 38335 21471
rect 38761 21437 38795 21471
rect 30573 21369 30607 21403
rect 30757 21369 30791 21403
rect 39037 21369 39071 21403
rect 28917 21301 28951 21335
rect 36093 21301 36127 21335
rect 1501 21097 1535 21131
rect 20085 21097 20119 21131
rect 28917 21029 28951 21063
rect 29285 21029 29319 21063
rect 32413 21029 32447 21063
rect 50813 21029 50847 21063
rect 1593 20961 1627 20995
rect 20177 20961 20211 20995
rect 20637 20961 20671 20995
rect 27905 20961 27939 20995
rect 28181 20961 28215 20995
rect 30941 20961 30975 20995
rect 31677 20961 31711 20995
rect 32229 20961 32263 20995
rect 36001 20961 36035 20995
rect 36553 20961 36587 20995
rect 37197 20961 37231 20995
rect 37381 20961 37415 20995
rect 37841 20961 37875 20995
rect 38025 20961 38059 20995
rect 38853 20961 38887 20995
rect 48145 20961 48179 20995
rect 48237 20961 48271 20995
rect 57529 20961 57563 20995
rect 58173 20961 58207 20995
rect 27721 20893 27755 20927
rect 30665 20893 30699 20927
rect 36093 20893 36127 20927
rect 37013 20893 37047 20927
rect 38761 20893 38795 20927
rect 48329 20893 48363 20927
rect 50813 20893 50847 20927
rect 38117 20825 38151 20859
rect 57989 20825 58023 20859
rect 47225 20757 47259 20791
rect 47777 20757 47811 20791
rect 1593 20553 1627 20587
rect 38393 20553 38427 20587
rect 47409 20553 47443 20587
rect 1409 20349 1443 20383
rect 2053 20349 2087 20383
rect 22845 20349 22879 20383
rect 23121 20349 23155 20383
rect 31401 20349 31435 20383
rect 31677 20349 31711 20383
rect 36553 20349 36587 20383
rect 36829 20349 36863 20383
rect 38485 20349 38519 20383
rect 31769 20281 31803 20315
rect 2697 20213 2731 20247
rect 23305 20213 23339 20247
rect 36369 20213 36403 20247
rect 38945 20213 38979 20247
rect 2421 20009 2455 20043
rect 3065 20009 3099 20043
rect 15945 20009 15979 20043
rect 17877 20009 17911 20043
rect 21925 20009 21959 20043
rect 32689 19941 32723 19975
rect 36461 19941 36495 19975
rect 2329 19873 2363 19907
rect 2513 19873 2547 19907
rect 2973 19873 3007 19907
rect 3157 19873 3191 19907
rect 15853 19873 15887 19907
rect 16037 19873 16071 19907
rect 16773 19873 16807 19907
rect 17785 19873 17819 19907
rect 21833 19873 21867 19907
rect 22477 19873 22511 19907
rect 31125 19873 31159 19907
rect 31401 19873 31435 19907
rect 32045 19873 32079 19907
rect 32137 19873 32171 19907
rect 32597 19873 32631 19907
rect 36369 19873 36403 19907
rect 37013 19873 37047 19907
rect 37289 19873 37323 19907
rect 57989 19873 58023 19907
rect 31401 19737 31435 19771
rect 37289 19737 37323 19771
rect 57345 19737 57379 19771
rect 58173 19737 58207 19771
rect 3985 19669 4019 19703
rect 18521 19669 18555 19703
rect 35817 19669 35851 19703
rect 2329 19465 2363 19499
rect 16221 19329 16255 19363
rect 1409 19261 1443 19295
rect 2237 19261 2271 19295
rect 8677 19261 8711 19295
rect 8769 19261 8803 19295
rect 57989 19193 58023 19227
rect 58173 19193 58207 19227
rect 1593 19125 1627 19159
rect 32781 19125 32815 19159
rect 57345 19125 57379 19159
rect 1409 18921 1443 18955
rect 2329 18921 2363 18955
rect 26525 18921 26559 18955
rect 26433 18785 26467 18819
rect 26617 18785 26651 18819
rect 27445 18785 27479 18819
rect 27905 18785 27939 18819
rect 2421 18717 2455 18751
rect 2605 18717 2639 18751
rect 28181 18717 28215 18751
rect 3249 18649 3283 18683
rect 1961 18581 1995 18615
rect 1593 18377 1627 18411
rect 2605 18377 2639 18411
rect 1409 18173 1443 18207
rect 2053 18173 2087 18207
rect 27077 17833 27111 17867
rect 27905 17833 27939 17867
rect 55229 17833 55263 17867
rect 57989 17833 58023 17867
rect 26341 17765 26375 17799
rect 27813 17765 27847 17799
rect 1409 17697 1443 17731
rect 1593 17697 1627 17731
rect 27261 17697 27295 17731
rect 54217 17697 54251 17731
rect 55137 17697 55171 17731
rect 57529 17697 57563 17731
rect 58173 17697 58207 17731
rect 26525 17629 26559 17663
rect 55321 17629 55355 17663
rect 2237 17493 2271 17527
rect 54769 17493 54803 17527
rect 25421 17289 25455 17323
rect 54401 17289 54435 17323
rect 26065 17153 26099 17187
rect 8033 17085 8067 17119
rect 24869 17085 24903 17119
rect 25329 17085 25363 17119
rect 26617 17085 26651 17119
rect 36277 17085 36311 17119
rect 57897 17085 57931 17119
rect 36553 17017 36587 17051
rect 57437 17017 57471 17051
rect 58081 17017 58115 17051
rect 8125 16949 8159 16983
rect 10333 16745 10367 16779
rect 21281 16745 21315 16779
rect 22017 16677 22051 16711
rect 1501 16609 1535 16643
rect 10333 16609 10367 16643
rect 10609 16609 10643 16643
rect 21097 16609 21131 16643
rect 21741 16609 21775 16643
rect 22753 16609 22787 16643
rect 25697 16609 25731 16643
rect 26801 16609 26835 16643
rect 28641 16609 28675 16643
rect 29193 16609 29227 16643
rect 29377 16609 29411 16643
rect 37105 16609 37139 16643
rect 38025 16609 38059 16643
rect 44649 16609 44683 16643
rect 57989 16609 58023 16643
rect 11161 16541 11195 16575
rect 37381 16541 37415 16575
rect 29377 16473 29411 16507
rect 58173 16473 58207 16507
rect 1593 16405 1627 16439
rect 20637 16405 20671 16439
rect 23029 16405 23063 16439
rect 25513 16405 25547 16439
rect 26617 16405 26651 16439
rect 38209 16405 38243 16439
rect 44557 16405 44591 16439
rect 45201 16405 45235 16439
rect 1409 16201 1443 16235
rect 29929 16201 29963 16235
rect 18337 16133 18371 16167
rect 25973 16133 26007 16167
rect 29377 16133 29411 16167
rect 21097 16065 21131 16099
rect 23305 16065 23339 16099
rect 40877 16065 40911 16099
rect 43545 16065 43579 16099
rect 8493 15997 8527 16031
rect 8769 15997 8803 16031
rect 18521 15997 18555 16031
rect 21373 15997 21407 16031
rect 23213 15997 23247 16031
rect 23765 15997 23799 16031
rect 29101 15997 29135 16031
rect 29285 15997 29319 16031
rect 30113 15997 30147 16031
rect 30573 15997 30607 16031
rect 36001 15997 36035 16031
rect 37013 15997 37047 16031
rect 38761 15997 38795 16031
rect 38853 15997 38887 16031
rect 40693 15997 40727 16031
rect 40969 15997 41003 16031
rect 43637 15997 43671 16031
rect 43821 15997 43855 16031
rect 44373 15997 44407 16031
rect 44557 15997 44591 16031
rect 8401 15929 8435 15963
rect 9321 15929 9355 15963
rect 22569 15929 22603 15963
rect 26249 15929 26283 15963
rect 39037 15929 39071 15963
rect 44741 15929 44775 15963
rect 28549 15861 28583 15895
rect 35909 15861 35943 15895
rect 37289 15861 37323 15895
rect 1593 15657 1627 15691
rect 22017 15657 22051 15691
rect 28549 15657 28583 15691
rect 36093 15657 36127 15691
rect 37105 15657 37139 15691
rect 37749 15657 37783 15691
rect 33701 15589 33735 15623
rect 1409 15521 1443 15555
rect 17693 15521 17727 15555
rect 17877 15521 17911 15555
rect 18797 15521 18831 15555
rect 22109 15521 22143 15555
rect 25237 15521 25271 15555
rect 28457 15521 28491 15555
rect 29101 15521 29135 15555
rect 32413 15521 32447 15555
rect 32965 15521 32999 15555
rect 33057 15521 33091 15555
rect 37657 15521 37691 15555
rect 38577 15521 38611 15555
rect 38853 15521 38887 15555
rect 40969 15521 41003 15555
rect 41521 15521 41555 15555
rect 17601 15453 17635 15487
rect 25421 15453 25455 15487
rect 33241 15453 33275 15487
rect 38669 15453 38703 15487
rect 41429 15453 41463 15487
rect 18981 15317 19015 15351
rect 1409 15113 1443 15147
rect 18889 15113 18923 15147
rect 18153 14977 18187 15011
rect 17877 14909 17911 14943
rect 18061 14909 18095 14943
rect 36829 14909 36863 14943
rect 37013 14909 37047 14943
rect 57437 14909 57471 14943
rect 58173 14909 58207 14943
rect 36645 14841 36679 14875
rect 57989 14773 58023 14807
rect 23673 14501 23707 14535
rect 52469 14501 52503 14535
rect 1409 14433 1443 14467
rect 2053 14433 2087 14467
rect 14933 14433 14967 14467
rect 15485 14433 15519 14467
rect 22477 14433 22511 14467
rect 37105 14433 37139 14467
rect 52009 14433 52043 14467
rect 52929 14433 52963 14467
rect 53113 14433 53147 14467
rect 57529 14433 57563 14467
rect 58173 14433 58207 14467
rect 53205 14365 53239 14399
rect 1593 14297 1627 14331
rect 22569 14297 22603 14331
rect 37013 14297 37047 14331
rect 57989 14297 58023 14331
rect 14841 14229 14875 14263
rect 23581 14229 23615 14263
rect 1409 13821 1443 13855
rect 2053 13821 2087 13855
rect 10609 13821 10643 13855
rect 10793 13821 10827 13855
rect 11805 13821 11839 13855
rect 13553 13821 13587 13855
rect 13737 13821 13771 13855
rect 14381 13821 14415 13855
rect 22845 13821 22879 13855
rect 23029 13821 23063 13855
rect 35357 13821 35391 13855
rect 35633 13821 35667 13855
rect 10425 13753 10459 13787
rect 13829 13753 13863 13787
rect 22661 13753 22695 13787
rect 1593 13685 1627 13719
rect 23581 13685 23615 13719
rect 34621 13685 34655 13719
rect 35817 13685 35851 13719
rect 2421 13481 2455 13515
rect 1501 13413 1535 13447
rect 11253 13413 11287 13447
rect 2329 13345 2363 13379
rect 10333 13345 10367 13379
rect 10517 13345 10551 13379
rect 11345 13345 11379 13379
rect 12817 13345 12851 13379
rect 13001 13345 13035 13379
rect 13553 13345 13587 13379
rect 2513 13277 2547 13311
rect 12633 13277 12667 13311
rect 10241 13209 10275 13243
rect 1961 13141 1995 13175
rect 3249 13141 3283 13175
rect 11897 13141 11931 13175
rect 10609 12937 10643 12971
rect 1409 12801 1443 12835
rect 57437 12801 57471 12835
rect 58081 12733 58115 12767
rect 1593 12665 1627 12699
rect 57897 12665 57931 12699
rect 2145 12597 2179 12631
rect 57437 12257 57471 12291
rect 58173 12257 58207 12291
rect 57989 12121 58023 12155
rect 1409 11577 1443 11611
rect 1593 11577 1627 11611
rect 2237 11577 2271 11611
rect 57989 11577 58023 11611
rect 58173 11577 58207 11611
rect 57897 11305 57931 11339
rect 57529 11237 57563 11271
rect 1593 11169 1627 11203
rect 2237 11169 2271 11203
rect 57253 11101 57287 11135
rect 57437 11101 57471 11135
rect 1501 10965 1535 10999
rect 56701 10965 56735 10999
rect 23857 10761 23891 10795
rect 24593 10557 24627 10591
rect 24777 10557 24811 10591
rect 24409 10489 24443 10523
rect 56793 10421 56827 10455
rect 57437 10149 57471 10183
rect 57989 10149 58023 10183
rect 58173 10149 58207 10183
rect 1501 9877 1535 9911
rect 34621 9605 34655 9639
rect 58173 9537 58207 9571
rect 1501 9469 1535 9503
rect 35173 9469 35207 9503
rect 35357 9469 35391 9503
rect 57989 9401 58023 9435
rect 1593 9333 1627 9367
rect 35449 9333 35483 9367
rect 57345 9333 57379 9367
rect 1593 9061 1627 9095
rect 1409 8857 1443 8891
rect 9229 8585 9263 8619
rect 10517 8585 10551 8619
rect 26525 8585 26559 8619
rect 8769 8449 8803 8483
rect 9873 8449 9907 8483
rect 9597 8381 9631 8415
rect 1593 8313 1627 8347
rect 2237 8313 2271 8347
rect 57345 8313 57379 8347
rect 57989 8313 58023 8347
rect 58173 8313 58207 8347
rect 1501 8245 1535 8279
rect 9689 8245 9723 8279
rect 25789 8041 25823 8075
rect 25789 7905 25823 7939
rect 26065 7905 26099 7939
rect 26893 7905 26927 7939
rect 26985 7905 27019 7939
rect 26709 7837 26743 7871
rect 26249 7497 26283 7531
rect 28089 7497 28123 7531
rect 1409 7293 1443 7327
rect 2053 7293 2087 7327
rect 28181 7293 28215 7327
rect 57529 7293 57563 7327
rect 58173 7293 58207 7327
rect 28733 7225 28767 7259
rect 1593 7157 1627 7191
rect 57989 7157 58023 7191
rect 1501 6953 1535 6987
rect 2421 6953 2455 6987
rect 57897 6885 57931 6919
rect 2329 6817 2363 6851
rect 54125 6817 54159 6851
rect 58081 6817 58115 6851
rect 2513 6749 2547 6783
rect 57437 6749 57471 6783
rect 3249 6681 3283 6715
rect 1961 6613 1995 6647
rect 54033 6613 54067 6647
rect 1593 6205 1627 6239
rect 1409 6137 1443 6171
rect 57713 6069 57747 6103
rect 57989 5729 58023 5763
rect 58173 5593 58207 5627
rect 40785 5525 40819 5559
rect 57069 5525 57103 5559
rect 17049 5321 17083 5355
rect 33977 5321 34011 5355
rect 2053 5253 2087 5287
rect 34805 5185 34839 5219
rect 35725 5185 35759 5219
rect 39589 5185 39623 5219
rect 40233 5185 40267 5219
rect 41429 5185 41463 5219
rect 56425 5185 56459 5219
rect 57529 5185 57563 5219
rect 25329 5117 25363 5151
rect 25421 5117 25455 5151
rect 34621 5117 34655 5151
rect 58173 5117 58207 5151
rect 1409 4981 1443 5015
rect 34713 4981 34747 5015
rect 35191 4981 35225 5015
rect 40785 4981 40819 5015
rect 56977 4981 57011 5015
rect 57989 4981 58023 5015
rect 2421 4777 2455 4811
rect 26433 4777 26467 4811
rect 1501 4709 1535 4743
rect 37657 4709 37691 4743
rect 42625 4709 42659 4743
rect 56793 4709 56827 4743
rect 58081 4709 58115 4743
rect 27445 4641 27479 4675
rect 29929 4641 29963 4675
rect 40969 4641 41003 4675
rect 57437 4641 57471 4675
rect 29285 4573 29319 4607
rect 1685 4505 1719 4539
rect 38761 4505 38795 4539
rect 57897 4505 57931 4539
rect 15853 4437 15887 4471
rect 16497 4437 16531 4471
rect 17509 4437 17543 4471
rect 28733 4437 28767 4471
rect 29929 4437 29963 4471
rect 37105 4437 37139 4471
rect 39773 4437 39807 4471
rect 41153 4437 41187 4471
rect 42165 4437 42199 4471
rect 43269 4437 43303 4471
rect 43821 4437 43855 4471
rect 44373 4437 44407 4471
rect 57253 4437 57287 4471
rect 3801 4233 3835 4267
rect 10333 4233 10367 4267
rect 19349 4233 19383 4267
rect 22753 4233 22787 4267
rect 26341 4233 26375 4267
rect 28917 4233 28951 4267
rect 29469 4233 29503 4267
rect 37013 4233 37047 4267
rect 40877 4233 40911 4267
rect 57989 4233 58023 4267
rect 15393 4165 15427 4199
rect 1409 4097 1443 4131
rect 45201 4097 45235 4131
rect 55137 4097 55171 4131
rect 1593 4029 1627 4063
rect 2329 4029 2363 4063
rect 15209 4029 15243 4063
rect 15853 4029 15887 4063
rect 17693 4029 17727 4063
rect 18153 4029 18187 4063
rect 25053 4029 25087 4063
rect 25237 4029 25271 4063
rect 25697 4029 25731 4063
rect 25881 4029 25915 4063
rect 36829 4029 36863 4063
rect 40049 4029 40083 4063
rect 40233 4029 40267 4063
rect 40877 4029 40911 4063
rect 40969 4029 41003 4063
rect 41153 4029 41187 4063
rect 41705 4029 41739 4063
rect 41797 4029 41831 4063
rect 42441 4029 42475 4063
rect 44097 4029 44131 4063
rect 56333 4029 56367 4063
rect 57345 4029 57379 4063
rect 58173 4029 58207 4063
rect 2145 3961 2179 3995
rect 17049 3961 17083 3995
rect 24593 3961 24627 3995
rect 36185 3961 36219 3995
rect 45753 3961 45787 3995
rect 56885 3961 56919 3995
rect 3157 3893 3191 3927
rect 17509 3893 17543 3927
rect 18705 3893 18739 3927
rect 21189 3893 21223 3927
rect 25145 3893 25179 3927
rect 25789 3893 25823 3927
rect 27629 3893 27663 3927
rect 28181 3893 28215 3927
rect 35541 3893 35575 3927
rect 38301 3893 38335 3927
rect 38945 3893 38979 3927
rect 39497 3893 39531 3927
rect 40141 3893 40175 3927
rect 41061 3893 41095 3927
rect 42257 3893 42291 3927
rect 43453 3893 43487 3927
rect 44557 3893 44591 3927
rect 46305 3893 46339 3927
rect 46857 3893 46891 3927
rect 47593 3893 47627 3927
rect 55689 3893 55723 3927
rect 57529 3893 57563 3927
rect 11529 3689 11563 3723
rect 14381 3689 14415 3723
rect 15577 3689 15611 3723
rect 22569 3689 22603 3723
rect 25789 3689 25823 3723
rect 30481 3689 30515 3723
rect 31677 3689 31711 3723
rect 32413 3689 32447 3723
rect 35725 3689 35759 3723
rect 38853 3689 38887 3723
rect 43913 3689 43947 3723
rect 2329 3621 2363 3655
rect 3065 3621 3099 3655
rect 47869 3621 47903 3655
rect 57989 3621 58023 3655
rect 1593 3553 1627 3587
rect 4445 3553 4479 3587
rect 9505 3553 9539 3587
rect 10149 3553 10183 3587
rect 14933 3553 14967 3587
rect 15117 3553 15151 3587
rect 16221 3553 16255 3587
rect 16313 3553 16347 3587
rect 16773 3553 16807 3587
rect 17417 3553 17451 3587
rect 18429 3553 18463 3587
rect 22753 3553 22787 3587
rect 23213 3553 23247 3587
rect 25237 3553 25271 3587
rect 25881 3553 25915 3587
rect 27353 3553 27387 3587
rect 27905 3553 27939 3587
rect 28733 3553 28767 3587
rect 29285 3553 29319 3587
rect 30665 3553 30699 3587
rect 31125 3553 31159 3587
rect 32229 3553 32263 3587
rect 32873 3553 32907 3587
rect 34069 3553 34103 3587
rect 34713 3553 34747 3587
rect 35909 3553 35943 3587
rect 36553 3553 36587 3587
rect 37289 3553 37323 3587
rect 38025 3553 38059 3587
rect 38669 3553 38703 3587
rect 39773 3553 39807 3587
rect 41153 3553 41187 3587
rect 42073 3553 42107 3587
rect 43361 3553 43395 3587
rect 44005 3553 44039 3587
rect 44649 3553 44683 3587
rect 48053 3553 48087 3587
rect 57253 3553 57287 3587
rect 45109 3485 45143 3519
rect 48605 3485 48639 3519
rect 55781 3485 55815 3519
rect 2881 3417 2915 3451
rect 9689 3417 9723 3451
rect 16957 3417 16991 3451
rect 26617 3417 26651 3451
rect 27169 3417 27203 3451
rect 28089 3417 28123 3451
rect 36369 3417 36403 3451
rect 39589 3417 39623 3451
rect 41889 3417 41923 3451
rect 54309 3417 54343 3451
rect 57437 3417 57471 3451
rect 58173 3417 58207 3451
rect 1501 3349 1535 3383
rect 2237 3349 2271 3383
rect 3893 3349 3927 3383
rect 6653 3349 6687 3383
rect 10977 3349 11011 3383
rect 13277 3349 13311 3383
rect 15117 3349 15151 3383
rect 17509 3349 17543 3383
rect 18613 3349 18647 3383
rect 19625 3349 19659 3383
rect 20269 3349 20303 3383
rect 21005 3349 21039 3383
rect 22017 3349 22051 3383
rect 24317 3349 24351 3383
rect 28641 3349 28675 3383
rect 29377 3349 29411 3383
rect 34253 3349 34287 3383
rect 37197 3349 37231 3383
rect 38209 3349 38243 3383
rect 41061 3349 41095 3383
rect 42717 3349 42751 3383
rect 43177 3349 43211 3383
rect 44465 3349 44499 3383
rect 45845 3349 45879 3383
rect 46397 3349 46431 3383
rect 47317 3349 47351 3383
rect 49617 3349 49651 3383
rect 50077 3349 50111 3383
rect 52101 3349 52135 3383
rect 52561 3349 52595 3383
rect 53205 3349 53239 3383
rect 53757 3349 53791 3383
rect 55229 3349 55263 3383
rect 56333 3349 56367 3383
rect 7021 3145 7055 3179
rect 8769 3145 8803 3179
rect 9689 3145 9723 3179
rect 13737 3145 13771 3179
rect 15393 3145 15427 3179
rect 17049 3145 17083 3179
rect 19809 3145 19843 3179
rect 27813 3145 27847 3179
rect 47041 3145 47075 3179
rect 53113 3145 53147 3179
rect 57253 3145 57287 3179
rect 38393 3077 38427 3111
rect 41705 3077 41739 3111
rect 42349 3077 42383 3111
rect 43637 3077 43671 3111
rect 45477 3077 45511 3111
rect 49709 3077 49743 3111
rect 55965 3077 55999 3111
rect 3525 3009 3559 3043
rect 28365 3009 28399 3043
rect 29929 3009 29963 3043
rect 34713 3009 34747 3043
rect 36185 3009 36219 3043
rect 39313 3009 39347 3043
rect 41061 3009 41095 3043
rect 41245 3009 41279 3043
rect 44097 3009 44131 3043
rect 57805 3009 57839 3043
rect 1409 2941 1443 2975
rect 2145 2941 2179 2975
rect 2973 2941 3007 2975
rect 4353 2941 4387 2975
rect 6837 2941 6871 2975
rect 8953 2941 8987 2975
rect 9873 2941 9907 2975
rect 10333 2941 10367 2975
rect 11069 2941 11103 2975
rect 13093 2941 13127 2975
rect 15393 2941 15427 2975
rect 15577 2941 15611 2975
rect 16313 2941 16347 2975
rect 17969 2941 18003 2975
rect 19073 2941 19107 2975
rect 19625 2941 19659 2975
rect 20729 2941 20763 2975
rect 22753 2941 22787 2975
rect 23673 2941 23707 2975
rect 24409 2941 24443 2975
rect 25145 2941 25179 2975
rect 25973 2941 26007 2975
rect 26709 2941 26743 2975
rect 28181 2941 28215 2975
rect 28273 2941 28307 2975
rect 29193 2941 29227 2975
rect 29837 2941 29871 2975
rect 31125 2941 31159 2975
rect 31953 2941 31987 2975
rect 33149 2941 33183 2975
rect 33609 2941 33643 2975
rect 34621 2941 34655 2975
rect 36461 2941 36495 2975
rect 37105 2941 37139 2975
rect 38301 2941 38335 2975
rect 39957 2941 39991 2975
rect 40325 2941 40359 2975
rect 41337 2941 41371 2975
rect 45661 2941 45695 2975
rect 46305 2941 46339 2975
rect 47133 2941 47167 2975
rect 47685 2941 47719 2975
rect 47869 2941 47903 2975
rect 49893 2941 49927 2975
rect 51733 2941 51767 2975
rect 52469 2941 52503 2975
rect 52929 2941 52963 2975
rect 54033 2941 54067 2975
rect 54217 2941 54251 2975
rect 54953 2941 54987 2975
rect 55781 2941 55815 2975
rect 57529 2941 57563 2975
rect 2329 2873 2363 2907
rect 2789 2873 2823 2907
rect 4169 2873 4203 2907
rect 4905 2873 4939 2907
rect 5089 2873 5123 2907
rect 5733 2873 5767 2907
rect 12909 2873 12943 2907
rect 14289 2873 14323 2907
rect 14473 2873 14507 2907
rect 16129 2873 16163 2907
rect 24593 2873 24627 2907
rect 25329 2873 25363 2907
rect 25789 2873 25823 2907
rect 30941 2873 30975 2907
rect 31769 2873 31803 2907
rect 35265 2873 35299 2907
rect 39129 2873 39163 2907
rect 42533 2873 42567 2907
rect 44189 2873 44223 2907
rect 44741 2873 44775 2907
rect 44925 2873 44959 2907
rect 46489 2873 46523 2907
rect 48789 2873 48823 2907
rect 48973 2873 49007 2907
rect 50445 2873 50479 2907
rect 50629 2873 50663 2907
rect 51549 2873 51583 2907
rect 54769 2873 54803 2907
rect 56517 2873 56551 2907
rect 57713 2873 57747 2907
rect 1593 2805 1627 2839
rect 7757 2805 7791 2839
rect 10977 2805 11011 2839
rect 12081 2805 12115 2839
rect 19073 2805 19107 2839
rect 20913 2805 20947 2839
rect 21649 2805 21683 2839
rect 22569 2805 22603 2839
rect 23765 2805 23799 2839
rect 26801 2805 26835 2839
rect 33793 2805 33827 2839
rect 40049 2805 40083 2839
rect 44097 2805 44131 2839
rect 47777 2805 47811 2839
rect 52285 2805 52319 2839
rect 54125 2805 54159 2839
rect 56609 2805 56643 2839
rect 14933 2601 14967 2635
rect 15301 2601 15335 2635
rect 29377 2601 29411 2635
rect 33701 2601 33735 2635
rect 35081 2601 35115 2635
rect 37381 2601 37415 2635
rect 39957 2601 39991 2635
rect 43177 2601 43211 2635
rect 44005 2601 44039 2635
rect 44557 2601 44591 2635
rect 46949 2601 46983 2635
rect 52377 2601 52411 2635
rect 1685 2533 1719 2567
rect 8309 2533 8343 2567
rect 9229 2533 9263 2567
rect 9965 2533 9999 2567
rect 13829 2533 13863 2567
rect 15393 2533 15427 2567
rect 16313 2533 16347 2567
rect 18153 2533 18187 2567
rect 19073 2533 19107 2567
rect 20453 2533 20487 2567
rect 21833 2533 21867 2567
rect 23121 2533 23155 2567
rect 26985 2533 27019 2567
rect 27169 2533 27203 2567
rect 28641 2533 28675 2567
rect 30573 2533 30607 2567
rect 31493 2533 31527 2567
rect 48329 2533 48363 2567
rect 50629 2533 50663 2567
rect 55137 2533 55171 2567
rect 56609 2533 56643 2567
rect 2053 2465 2087 2499
rect 3157 2465 3191 2499
rect 4905 2465 4939 2499
rect 5641 2465 5675 2499
rect 6561 2465 6595 2499
rect 7481 2465 7515 2499
rect 10149 2465 10183 2499
rect 10701 2465 10735 2499
rect 12357 2465 12391 2499
rect 13093 2465 13127 2499
rect 16497 2465 16531 2499
rect 16681 2465 16715 2499
rect 21649 2465 21683 2499
rect 24133 2465 24167 2499
rect 25973 2465 26007 2499
rect 26341 2465 26375 2499
rect 28457 2465 28491 2499
rect 29377 2465 29411 2499
rect 29653 2465 29687 2499
rect 32505 2465 32539 2499
rect 33793 2465 33827 2499
rect 34897 2465 34931 2499
rect 35357 2465 35391 2499
rect 36277 2465 36311 2499
rect 36553 2465 36587 2499
rect 37565 2465 37599 2499
rect 37841 2465 37875 2499
rect 39129 2465 39163 2499
rect 40325 2465 40359 2499
rect 40417 2465 40451 2499
rect 41613 2465 41647 2499
rect 41797 2465 41831 2499
rect 43269 2465 43303 2499
rect 44925 2465 44959 2499
rect 45017 2465 45051 2499
rect 45753 2465 45787 2499
rect 45937 2465 45971 2499
rect 47317 2465 47351 2499
rect 3893 2397 3927 2431
rect 15577 2397 15611 2431
rect 18153 2397 18187 2431
rect 18245 2397 18279 2431
rect 21925 2397 21959 2431
rect 26065 2397 26099 2431
rect 40601 2397 40635 2431
rect 43177 2397 43211 2431
rect 45201 2397 45235 2431
rect 47409 2397 47443 2431
rect 47593 2397 47627 2431
rect 48605 2465 48639 2499
rect 50537 2465 50571 2499
rect 52469 2465 52503 2499
rect 53573 2465 53607 2499
rect 55873 2465 55907 2499
rect 57713 2465 57747 2499
rect 58081 2465 58115 2499
rect 50721 2397 50755 2431
rect 5089 2329 5123 2363
rect 8125 2329 8159 2363
rect 13277 2329 13311 2363
rect 18889 2329 18923 2363
rect 20269 2329 20303 2363
rect 22937 2329 22971 2363
rect 23949 2329 23983 2363
rect 25329 2329 25363 2363
rect 31309 2329 31343 2363
rect 32689 2329 32723 2363
rect 36553 2329 36587 2363
rect 41889 2329 41923 2363
rect 48329 2329 48363 2363
rect 54953 2329 54987 2363
rect 56425 2329 56459 2363
rect 3249 2261 3283 2295
rect 5733 2261 5767 2295
rect 7573 2261 7607 2295
rect 10793 2261 10827 2295
rect 12449 2261 12483 2295
rect 13921 2261 13955 2295
rect 17693 2261 17727 2295
rect 21373 2261 21407 2295
rect 39037 2261 39071 2295
rect 42717 2261 42751 2295
rect 48513 2261 48547 2295
rect 49341 2261 49375 2295
rect 50169 2261 50203 2295
rect 53481 2261 53515 2295
rect 55781 2261 55815 2295
rect 48329 1921 48363 1955
rect 48329 1717 48363 1751
<< metal1 >>
rect 17034 28092 17040 28144
rect 17092 28132 17098 28144
rect 18598 28132 18604 28144
rect 17092 28104 18604 28132
rect 17092 28092 17098 28104
rect 18598 28092 18604 28104
rect 18656 28092 18662 28144
rect 18966 28092 18972 28144
rect 19024 28132 19030 28144
rect 37458 28132 37464 28144
rect 19024 28104 37464 28132
rect 19024 28092 19030 28104
rect 37458 28092 37464 28104
rect 37516 28092 37522 28144
rect 16482 28024 16488 28076
rect 16540 28064 16546 28076
rect 24302 28064 24308 28076
rect 16540 28036 24308 28064
rect 16540 28024 16546 28036
rect 24302 28024 24308 28036
rect 24360 28024 24366 28076
rect 34330 28064 34336 28076
rect 30024 28036 34336 28064
rect 5718 27956 5724 28008
rect 5776 27996 5782 28008
rect 17402 27996 17408 28008
rect 5776 27968 17408 27996
rect 5776 27956 5782 27968
rect 17402 27956 17408 27968
rect 17460 27956 17466 28008
rect 20622 27956 20628 28008
rect 20680 27996 20686 28008
rect 29730 27996 29736 28008
rect 20680 27968 29736 27996
rect 20680 27956 20686 27968
rect 29730 27956 29736 27968
rect 29788 27956 29794 28008
rect 8018 27888 8024 27940
rect 8076 27928 8082 27940
rect 30024 27928 30052 28036
rect 34330 28024 34336 28036
rect 34388 28024 34394 28076
rect 33962 27956 33968 28008
rect 34020 27996 34026 28008
rect 45370 27996 45376 28008
rect 34020 27968 45376 27996
rect 34020 27956 34026 27968
rect 45370 27956 45376 27968
rect 45428 27956 45434 28008
rect 8076 27900 30052 27928
rect 8076 27888 8082 27900
rect 30190 27888 30196 27940
rect 30248 27928 30254 27940
rect 34606 27928 34612 27940
rect 30248 27900 34612 27928
rect 30248 27888 30254 27900
rect 34606 27888 34612 27900
rect 34664 27888 34670 27940
rect 9398 27820 9404 27872
rect 9456 27860 9462 27872
rect 47026 27860 47032 27872
rect 9456 27832 47032 27860
rect 9456 27820 9462 27832
rect 47026 27820 47032 27832
rect 47084 27820 47090 27872
rect 1104 27770 58880 27792
rect 1104 27718 20246 27770
rect 20298 27718 20310 27770
rect 20362 27718 20374 27770
rect 20426 27718 20438 27770
rect 20490 27718 39510 27770
rect 39562 27718 39574 27770
rect 39626 27718 39638 27770
rect 39690 27718 39702 27770
rect 39754 27718 58880 27770
rect 1104 27696 58880 27718
rect 3145 27659 3203 27665
rect 3145 27625 3157 27659
rect 3191 27656 3203 27659
rect 3234 27656 3240 27668
rect 3191 27628 3240 27656
rect 3191 27625 3203 27628
rect 3145 27619 3203 27625
rect 3234 27616 3240 27628
rect 3292 27616 3298 27668
rect 8018 27656 8024 27668
rect 7979 27628 8024 27656
rect 8018 27616 8024 27628
rect 8076 27616 8082 27668
rect 8110 27616 8116 27668
rect 8168 27656 8174 27668
rect 13814 27656 13820 27668
rect 8168 27628 10732 27656
rect 8168 27616 8174 27628
rect 2593 27591 2651 27597
rect 2593 27557 2605 27591
rect 2639 27588 2651 27591
rect 2774 27588 2780 27600
rect 2639 27560 2780 27588
rect 2639 27557 2651 27560
rect 2593 27551 2651 27557
rect 2774 27548 2780 27560
rect 2832 27548 2838 27600
rect 5534 27588 5540 27600
rect 5495 27560 5540 27588
rect 5534 27548 5540 27560
rect 5592 27548 5598 27600
rect 5718 27588 5724 27600
rect 5679 27560 5724 27588
rect 5718 27548 5724 27560
rect 5776 27548 5782 27600
rect 7834 27548 7840 27600
rect 7892 27588 7898 27600
rect 7929 27591 7987 27597
rect 7929 27588 7941 27591
rect 7892 27560 7941 27588
rect 7892 27548 7898 27560
rect 7929 27557 7941 27560
rect 7975 27588 7987 27591
rect 8573 27591 8631 27597
rect 8573 27588 8585 27591
rect 7975 27560 8585 27588
rect 7975 27557 7987 27560
rect 7929 27551 7987 27557
rect 8573 27557 8585 27560
rect 8619 27557 8631 27591
rect 9674 27588 9680 27600
rect 9635 27560 9680 27588
rect 8573 27551 8631 27557
rect 9674 27548 9680 27560
rect 9732 27548 9738 27600
rect 10594 27588 10600 27600
rect 10555 27560 10600 27588
rect 10594 27548 10600 27560
rect 10652 27548 10658 27600
rect 10704 27588 10732 27628
rect 11578 27628 12572 27656
rect 13775 27628 13820 27656
rect 11578 27588 11606 27628
rect 11974 27588 11980 27600
rect 10704 27560 11606 27588
rect 11935 27560 11980 27588
rect 11974 27548 11980 27560
rect 12032 27548 12038 27600
rect 12434 27588 12440 27600
rect 12395 27560 12440 27588
rect 12434 27548 12440 27560
rect 12492 27548 12498 27600
rect 12544 27588 12572 27628
rect 13814 27616 13820 27628
rect 13872 27616 13878 27668
rect 22005 27659 22063 27665
rect 14660 27628 21772 27656
rect 14660 27588 14688 27628
rect 12544 27560 14688 27588
rect 14734 27548 14740 27600
rect 14792 27588 14798 27600
rect 14921 27591 14979 27597
rect 14921 27588 14933 27591
rect 14792 27560 14933 27588
rect 14792 27548 14798 27560
rect 14921 27557 14933 27560
rect 14967 27557 14979 27591
rect 14921 27551 14979 27557
rect 15933 27591 15991 27597
rect 15933 27557 15945 27591
rect 15979 27588 15991 27591
rect 16114 27588 16120 27600
rect 15979 27560 16120 27588
rect 15979 27557 15991 27560
rect 15933 27551 15991 27557
rect 16114 27548 16120 27560
rect 16172 27548 16178 27600
rect 16482 27588 16488 27600
rect 16443 27560 16488 27588
rect 16482 27548 16488 27560
rect 16540 27548 16546 27600
rect 16669 27591 16727 27597
rect 16669 27557 16681 27591
rect 16715 27588 16727 27591
rect 17954 27588 17960 27600
rect 16715 27560 17960 27588
rect 16715 27557 16727 27560
rect 16669 27551 16727 27557
rect 17954 27548 17960 27560
rect 18012 27548 18018 27600
rect 19334 27588 19340 27600
rect 19295 27560 19340 27588
rect 19334 27548 19340 27560
rect 19392 27548 19398 27600
rect 20622 27548 20628 27600
rect 20680 27588 20686 27600
rect 20680 27560 20725 27588
rect 20680 27548 20686 27560
rect 934 27480 940 27532
rect 992 27520 998 27532
rect 1397 27523 1455 27529
rect 1397 27520 1409 27523
rect 992 27492 1409 27520
rect 992 27480 998 27492
rect 1397 27489 1409 27492
rect 1443 27520 1455 27523
rect 2222 27520 2228 27532
rect 1443 27492 2228 27520
rect 1443 27489 1455 27492
rect 1397 27483 1455 27489
rect 2222 27480 2228 27492
rect 2280 27480 2286 27532
rect 2409 27523 2467 27529
rect 2409 27489 2421 27523
rect 2455 27489 2467 27523
rect 3234 27520 3240 27532
rect 3195 27492 3240 27520
rect 2409 27483 2467 27489
rect 2424 27384 2452 27483
rect 3234 27480 3240 27492
rect 3292 27480 3298 27532
rect 3878 27480 3884 27532
rect 3936 27520 3942 27532
rect 4617 27523 4675 27529
rect 4617 27520 4629 27523
rect 3936 27492 4629 27520
rect 3936 27480 3942 27492
rect 4617 27489 4629 27492
rect 4663 27489 4675 27523
rect 4617 27483 4675 27489
rect 4709 27523 4767 27529
rect 4709 27489 4721 27523
rect 4755 27520 4767 27523
rect 5166 27520 5172 27532
rect 4755 27492 5172 27520
rect 4755 27489 4767 27492
rect 4709 27483 4767 27489
rect 5166 27480 5172 27492
rect 5224 27480 5230 27532
rect 7101 27523 7159 27529
rect 7101 27489 7113 27523
rect 7147 27489 7159 27523
rect 7101 27483 7159 27489
rect 9861 27523 9919 27529
rect 9861 27489 9873 27523
rect 9907 27489 9919 27523
rect 9861 27483 9919 27489
rect 4890 27452 4896 27464
rect 4851 27424 4896 27452
rect 4890 27412 4896 27424
rect 4948 27412 4954 27464
rect 6914 27384 6920 27396
rect 2424 27356 6454 27384
rect 6875 27356 6920 27384
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 1762 27316 1768 27328
rect 1627 27288 1768 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 1762 27276 1768 27288
rect 1820 27276 1826 27328
rect 4249 27319 4307 27325
rect 4249 27285 4261 27319
rect 4295 27316 4307 27319
rect 4430 27316 4436 27328
rect 4295 27288 4436 27316
rect 4295 27285 4307 27288
rect 4249 27279 4307 27285
rect 4430 27276 4436 27288
rect 4488 27276 4494 27328
rect 6426 27316 6454 27356
rect 6914 27344 6920 27356
rect 6972 27344 6978 27396
rect 7116 27384 7144 27483
rect 9876 27452 9904 27483
rect 10410 27480 10416 27532
rect 10468 27520 10474 27532
rect 10781 27523 10839 27529
rect 10781 27520 10793 27523
rect 10468 27492 10793 27520
rect 10468 27480 10474 27492
rect 10781 27489 10793 27492
rect 10827 27489 10839 27523
rect 10781 27483 10839 27489
rect 12621 27523 12679 27529
rect 12621 27489 12633 27523
rect 12667 27520 12679 27523
rect 13538 27520 13544 27532
rect 12667 27492 13544 27520
rect 12667 27489 12679 27492
rect 12621 27483 12679 27489
rect 13538 27480 13544 27492
rect 13596 27480 13602 27532
rect 13909 27523 13967 27529
rect 13909 27489 13921 27523
rect 13955 27489 13967 27523
rect 13909 27483 13967 27489
rect 13924 27452 13952 27483
rect 15010 27480 15016 27532
rect 15068 27520 15074 27532
rect 15105 27523 15163 27529
rect 15105 27520 15117 27523
rect 15068 27492 15117 27520
rect 15068 27480 15074 27492
rect 15105 27489 15117 27492
rect 15151 27489 15163 27523
rect 15105 27483 15163 27489
rect 15749 27523 15807 27529
rect 15749 27489 15761 27523
rect 15795 27520 15807 27523
rect 15838 27520 15844 27532
rect 15795 27492 15844 27520
rect 15795 27489 15807 27492
rect 15749 27483 15807 27489
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 17678 27520 17684 27532
rect 17639 27492 17684 27520
rect 17678 27480 17684 27492
rect 17736 27480 17742 27532
rect 17862 27520 17868 27532
rect 17823 27492 17868 27520
rect 17862 27480 17868 27492
rect 17920 27480 17926 27532
rect 18598 27520 18604 27532
rect 18559 27492 18604 27520
rect 18598 27480 18604 27492
rect 18656 27480 18662 27532
rect 19153 27523 19211 27529
rect 19153 27489 19165 27523
rect 19199 27520 19211 27523
rect 19794 27520 19800 27532
rect 19199 27492 19800 27520
rect 19199 27489 19211 27492
rect 19153 27483 19211 27489
rect 19794 27480 19800 27492
rect 19852 27480 19858 27532
rect 20254 27520 20260 27532
rect 20215 27492 20260 27520
rect 20254 27480 20260 27492
rect 20312 27480 20318 27532
rect 20438 27520 20444 27532
rect 20399 27492 20444 27520
rect 20438 27480 20444 27492
rect 20496 27480 20502 27532
rect 20530 27480 20536 27532
rect 20588 27520 20594 27532
rect 21269 27523 21327 27529
rect 21269 27520 21281 27523
rect 20588 27492 21281 27520
rect 20588 27480 20594 27492
rect 21269 27489 21281 27492
rect 21315 27489 21327 27523
rect 21269 27483 21327 27489
rect 17034 27452 17040 27464
rect 9876 27424 13308 27452
rect 13924 27424 17040 27452
rect 13280 27393 13308 27424
rect 17034 27412 17040 27424
rect 17092 27412 17098 27464
rect 17402 27412 17408 27464
rect 17460 27452 17466 27464
rect 17589 27455 17647 27461
rect 17589 27452 17601 27455
rect 17460 27424 17601 27452
rect 17460 27412 17466 27424
rect 17589 27421 17601 27424
rect 17635 27421 17647 27455
rect 17589 27415 17647 27421
rect 20714 27412 20720 27464
rect 20772 27452 20778 27464
rect 21085 27455 21143 27461
rect 21085 27452 21097 27455
rect 20772 27424 21097 27452
rect 20772 27412 20778 27424
rect 21085 27421 21097 27424
rect 21131 27421 21143 27455
rect 21744 27452 21772 27628
rect 22005 27625 22017 27659
rect 22051 27656 22063 27659
rect 25866 27656 25872 27668
rect 22051 27628 25872 27656
rect 22051 27625 22063 27628
rect 22005 27619 22063 27625
rect 25866 27616 25872 27628
rect 25924 27616 25930 27668
rect 29914 27656 29920 27668
rect 29875 27628 29920 27656
rect 29914 27616 29920 27628
rect 29972 27616 29978 27668
rect 31478 27616 31484 27668
rect 31536 27656 31542 27668
rect 37369 27659 37427 27665
rect 37369 27656 37381 27659
rect 31536 27628 37381 27656
rect 31536 27616 31542 27628
rect 37369 27625 37381 27628
rect 37415 27625 37427 27659
rect 37369 27619 37427 27625
rect 37826 27616 37832 27668
rect 37884 27656 37890 27668
rect 43165 27659 43223 27665
rect 37884 27628 42472 27656
rect 37884 27616 37890 27628
rect 23934 27588 23940 27600
rect 23895 27560 23940 27588
rect 23934 27548 23940 27560
rect 23992 27548 23998 27600
rect 24486 27548 24492 27600
rect 24544 27588 24550 27600
rect 25593 27591 25651 27597
rect 25593 27588 25605 27591
rect 24544 27560 25605 27588
rect 24544 27548 24550 27560
rect 25593 27557 25605 27560
rect 25639 27557 25651 27591
rect 25593 27551 25651 27557
rect 25777 27591 25835 27597
rect 25777 27557 25789 27591
rect 25823 27588 25835 27591
rect 28077 27591 28135 27597
rect 25823 27560 28028 27588
rect 25823 27557 25835 27560
rect 25777 27551 25835 27557
rect 21821 27523 21879 27529
rect 21821 27489 21833 27523
rect 21867 27520 21879 27523
rect 22094 27520 22100 27532
rect 21867 27492 22100 27520
rect 21867 27489 21879 27492
rect 21821 27483 21879 27489
rect 22094 27480 22100 27492
rect 22152 27520 22158 27532
rect 22557 27523 22615 27529
rect 22557 27520 22569 27523
rect 22152 27492 22569 27520
rect 22152 27480 22158 27492
rect 22557 27489 22569 27492
rect 22603 27489 22615 27523
rect 22557 27483 22615 27489
rect 23293 27523 23351 27529
rect 23293 27489 23305 27523
rect 23339 27520 23351 27523
rect 23750 27520 23756 27532
rect 23339 27492 23756 27520
rect 23339 27489 23351 27492
rect 23293 27483 23351 27489
rect 23750 27480 23756 27492
rect 23808 27480 23814 27532
rect 24118 27520 24124 27532
rect 24079 27492 24124 27520
rect 24118 27480 24124 27492
rect 24176 27480 24182 27532
rect 26789 27523 26847 27529
rect 26789 27520 26801 27523
rect 24228 27492 26801 27520
rect 24228 27452 24256 27492
rect 26789 27489 26801 27492
rect 26835 27489 26847 27523
rect 26789 27483 26847 27489
rect 26881 27523 26939 27529
rect 26881 27489 26893 27523
rect 26927 27489 26939 27523
rect 26881 27483 26939 27489
rect 21744 27424 24256 27452
rect 26896 27452 26924 27483
rect 26970 27480 26976 27532
rect 27028 27520 27034 27532
rect 27065 27523 27123 27529
rect 27065 27520 27077 27523
rect 27028 27492 27077 27520
rect 27028 27480 27034 27492
rect 27065 27489 27077 27492
rect 27111 27489 27123 27523
rect 27065 27483 27123 27489
rect 27246 27452 27252 27464
rect 26896 27424 27252 27452
rect 21085 27415 21143 27421
rect 27246 27412 27252 27424
rect 27304 27412 27310 27464
rect 28000 27452 28028 27560
rect 28077 27557 28089 27591
rect 28123 27588 28135 27591
rect 28534 27588 28540 27600
rect 28123 27560 28540 27588
rect 28123 27557 28135 27560
rect 28077 27551 28135 27557
rect 28534 27548 28540 27560
rect 28592 27588 28598 27600
rect 28629 27591 28687 27597
rect 28629 27588 28641 27591
rect 28592 27560 28641 27588
rect 28592 27548 28598 27560
rect 28629 27557 28641 27560
rect 28675 27557 28687 27591
rect 28629 27551 28687 27557
rect 29730 27548 29736 27600
rect 29788 27588 29794 27600
rect 32214 27588 32220 27600
rect 29788 27560 29960 27588
rect 29788 27548 29794 27560
rect 29362 27480 29368 27532
rect 29420 27520 29426 27532
rect 29825 27523 29883 27529
rect 29825 27520 29837 27523
rect 29420 27492 29837 27520
rect 29420 27480 29426 27492
rect 29825 27489 29837 27492
rect 29871 27489 29883 27523
rect 29932 27520 29960 27560
rect 31404 27560 31708 27588
rect 32175 27560 32220 27588
rect 31404 27520 31432 27560
rect 29932 27492 31432 27520
rect 31573 27523 31631 27529
rect 29825 27483 29883 27489
rect 31573 27489 31585 27523
rect 31619 27489 31631 27523
rect 31680 27520 31708 27560
rect 32214 27548 32220 27560
rect 32272 27548 32278 27600
rect 33962 27588 33968 27600
rect 33923 27560 33968 27588
rect 33962 27548 33968 27560
rect 34020 27548 34026 27600
rect 34146 27588 34152 27600
rect 34107 27560 34152 27588
rect 34146 27548 34152 27560
rect 34204 27548 34210 27600
rect 35434 27548 35440 27600
rect 35492 27588 35498 27600
rect 36265 27591 36323 27597
rect 36265 27588 36277 27591
rect 35492 27560 36277 27588
rect 35492 27548 35498 27560
rect 36265 27557 36277 27560
rect 36311 27557 36323 27591
rect 36265 27551 36323 27557
rect 37274 27548 37280 27600
rect 37332 27548 37338 27600
rect 37550 27597 37556 27600
rect 37532 27591 37556 27597
rect 37532 27557 37544 27591
rect 37532 27551 37556 27557
rect 37550 27548 37556 27551
rect 37608 27548 37614 27600
rect 37737 27591 37795 27597
rect 37737 27557 37749 27591
rect 37783 27588 37795 27591
rect 38010 27588 38016 27600
rect 37783 27560 38016 27588
rect 37783 27557 37795 27560
rect 37737 27551 37795 27557
rect 38010 27548 38016 27560
rect 38068 27548 38074 27600
rect 39485 27591 39543 27597
rect 39485 27557 39497 27591
rect 39531 27588 39543 27591
rect 40126 27588 40132 27600
rect 39531 27560 40132 27588
rect 39531 27557 39543 27560
rect 39485 27551 39543 27557
rect 40126 27548 40132 27560
rect 40184 27548 40190 27600
rect 42444 27597 42472 27628
rect 43165 27625 43177 27659
rect 43211 27656 43223 27659
rect 43254 27656 43260 27668
rect 43211 27628 43260 27656
rect 43211 27625 43223 27628
rect 43165 27619 43223 27625
rect 43254 27616 43260 27628
rect 43312 27616 43318 27668
rect 47026 27656 47032 27668
rect 46987 27628 47032 27656
rect 47026 27616 47032 27628
rect 47084 27616 47090 27668
rect 50525 27659 50583 27665
rect 50525 27625 50537 27659
rect 50571 27656 50583 27659
rect 52914 27656 52920 27668
rect 50571 27628 52920 27656
rect 50571 27625 50583 27628
rect 50525 27619 50583 27625
rect 52914 27616 52920 27628
rect 52972 27616 52978 27668
rect 54754 27616 54760 27668
rect 54812 27656 54818 27668
rect 56505 27659 56563 27665
rect 56505 27656 56517 27659
rect 54812 27628 56517 27656
rect 54812 27616 54818 27628
rect 56505 27625 56517 27628
rect 56551 27625 56563 27659
rect 56505 27619 56563 27625
rect 42429 27591 42487 27597
rect 42429 27557 42441 27591
rect 42475 27557 42487 27591
rect 42429 27551 42487 27557
rect 42613 27591 42671 27597
rect 42613 27557 42625 27591
rect 42659 27588 42671 27591
rect 42794 27588 42800 27600
rect 42659 27560 42800 27588
rect 42659 27557 42671 27560
rect 42613 27551 42671 27557
rect 42794 27548 42800 27560
rect 42852 27548 42858 27600
rect 43806 27548 43812 27600
rect 43864 27588 43870 27600
rect 44269 27591 44327 27597
rect 44269 27588 44281 27591
rect 43864 27560 44281 27588
rect 43864 27548 43870 27560
rect 44269 27557 44281 27560
rect 44315 27557 44327 27591
rect 44269 27551 44327 27557
rect 45281 27591 45339 27597
rect 45281 27557 45293 27591
rect 45327 27588 45339 27591
rect 45554 27588 45560 27600
rect 45327 27560 45560 27588
rect 45327 27557 45339 27560
rect 45281 27551 45339 27557
rect 45554 27548 45560 27560
rect 45612 27548 45618 27600
rect 46017 27591 46075 27597
rect 46017 27557 46029 27591
rect 46063 27588 46075 27591
rect 46474 27588 46480 27600
rect 46063 27560 46480 27588
rect 46063 27557 46075 27560
rect 46017 27551 46075 27557
rect 46474 27548 46480 27560
rect 46532 27548 46538 27600
rect 46934 27548 46940 27600
rect 46992 27588 46998 27600
rect 47121 27591 47179 27597
rect 47121 27588 47133 27591
rect 46992 27560 47133 27588
rect 46992 27548 46998 27560
rect 47121 27557 47133 27560
rect 47167 27588 47179 27591
rect 47673 27591 47731 27597
rect 47673 27588 47685 27591
rect 47167 27560 47685 27588
rect 47167 27557 47179 27560
rect 47121 27551 47179 27557
rect 47673 27557 47685 27560
rect 47719 27557 47731 27591
rect 47673 27551 47731 27557
rect 48314 27548 48320 27600
rect 48372 27588 48378 27600
rect 48501 27591 48559 27597
rect 48501 27588 48513 27591
rect 48372 27560 48513 27588
rect 48372 27548 48378 27560
rect 48501 27557 48513 27560
rect 48547 27557 48559 27591
rect 48501 27551 48559 27557
rect 48958 27548 48964 27600
rect 49016 27588 49022 27600
rect 49605 27591 49663 27597
rect 49605 27588 49617 27591
rect 49016 27560 49617 27588
rect 49016 27548 49022 27560
rect 49605 27557 49617 27560
rect 49651 27557 49663 27591
rect 49605 27551 49663 27557
rect 51261 27591 51319 27597
rect 51261 27557 51273 27591
rect 51307 27588 51319 27591
rect 51534 27588 51540 27600
rect 51307 27560 51540 27588
rect 51307 27557 51319 27560
rect 51261 27551 51319 27557
rect 51534 27548 51540 27560
rect 51592 27548 51598 27600
rect 51994 27548 52000 27600
rect 52052 27588 52058 27600
rect 52457 27591 52515 27597
rect 52457 27588 52469 27591
rect 52052 27560 52469 27588
rect 52052 27548 52058 27560
rect 52457 27557 52469 27560
rect 52503 27557 52515 27591
rect 52457 27551 52515 27557
rect 53374 27548 53380 27600
rect 53432 27588 53438 27600
rect 53561 27591 53619 27597
rect 53561 27588 53573 27591
rect 53432 27560 53573 27588
rect 53432 27548 53438 27560
rect 53561 27557 53573 27560
rect 53607 27557 53619 27591
rect 53561 27551 53619 27557
rect 54294 27548 54300 27600
rect 54352 27588 54358 27600
rect 54941 27591 54999 27597
rect 54941 27588 54953 27591
rect 54352 27560 54953 27588
rect 54352 27548 54358 27560
rect 54941 27557 54953 27560
rect 54987 27557 54999 27591
rect 54941 27551 54999 27557
rect 55214 27548 55220 27600
rect 55272 27588 55278 27600
rect 55677 27591 55735 27597
rect 55677 27588 55689 27591
rect 55272 27560 55689 27588
rect 55272 27548 55278 27560
rect 55677 27557 55689 27560
rect 55723 27557 55735 27591
rect 55677 27551 55735 27557
rect 57974 27548 57980 27600
rect 58032 27588 58038 27600
rect 58069 27591 58127 27597
rect 58069 27588 58081 27591
rect 58032 27560 58081 27588
rect 58032 27548 58038 27560
rect 58069 27557 58081 27560
rect 58115 27557 58127 27591
rect 58069 27551 58127 27557
rect 32401 27523 32459 27529
rect 32401 27520 32413 27523
rect 31680 27492 32413 27520
rect 31573 27483 31631 27489
rect 32401 27489 32413 27492
rect 32447 27489 32459 27523
rect 32401 27483 32459 27489
rect 31478 27452 31484 27464
rect 28000 27424 31484 27452
rect 31478 27412 31484 27424
rect 31536 27412 31542 27464
rect 13265 27387 13323 27393
rect 7116 27356 11606 27384
rect 9858 27316 9864 27328
rect 6426 27288 9864 27316
rect 9858 27276 9864 27288
rect 9916 27276 9922 27328
rect 11578 27316 11606 27356
rect 13265 27353 13277 27387
rect 13311 27384 13323 27387
rect 30282 27384 30288 27396
rect 13311 27356 25912 27384
rect 13311 27353 13323 27356
rect 13265 27347 13323 27353
rect 17126 27316 17132 27328
rect 11578 27288 17132 27316
rect 17126 27276 17132 27288
rect 17184 27276 17190 27328
rect 17494 27276 17500 27328
rect 17552 27316 17558 27328
rect 18417 27319 18475 27325
rect 18417 27316 18429 27319
rect 17552 27288 18429 27316
rect 17552 27276 17558 27288
rect 18417 27285 18429 27288
rect 18463 27285 18475 27319
rect 18417 27279 18475 27285
rect 23385 27319 23443 27325
rect 23385 27285 23397 27319
rect 23431 27316 23443 27319
rect 25774 27316 25780 27328
rect 23431 27288 25780 27316
rect 23431 27285 23443 27288
rect 23385 27279 23443 27285
rect 25774 27276 25780 27288
rect 25832 27276 25838 27328
rect 25884 27316 25912 27356
rect 26988 27356 30288 27384
rect 26988 27316 27016 27356
rect 30282 27344 30288 27356
rect 30340 27344 30346 27396
rect 31588 27384 31616 27483
rect 33594 27480 33600 27532
rect 33652 27520 33658 27532
rect 34422 27520 34428 27532
rect 33652 27492 34428 27520
rect 33652 27480 33658 27492
rect 34422 27480 34428 27492
rect 34480 27520 34486 27532
rect 34977 27523 35035 27529
rect 34977 27520 34989 27523
rect 34480 27492 34989 27520
rect 34480 27480 34486 27492
rect 34977 27489 34989 27492
rect 35023 27489 35035 27523
rect 34977 27483 35035 27489
rect 36449 27523 36507 27529
rect 36449 27489 36461 27523
rect 36495 27520 36507 27523
rect 36630 27520 36636 27532
rect 36495 27492 36636 27520
rect 36495 27489 36507 27492
rect 36449 27483 36507 27489
rect 36630 27480 36636 27492
rect 36688 27480 36694 27532
rect 33502 27412 33508 27464
rect 33560 27452 33566 27464
rect 34241 27455 34299 27461
rect 34241 27452 34253 27455
rect 33560 27424 34253 27452
rect 33560 27412 33566 27424
rect 34241 27421 34253 27424
rect 34287 27421 34299 27455
rect 37292 27452 37320 27548
rect 39298 27520 39304 27532
rect 39259 27492 39304 27520
rect 39298 27480 39304 27492
rect 39356 27480 39362 27532
rect 40218 27480 40224 27532
rect 40276 27520 40282 27532
rect 40313 27523 40371 27529
rect 40313 27520 40325 27523
rect 40276 27492 40325 27520
rect 40276 27480 40282 27492
rect 40313 27489 40325 27492
rect 40359 27489 40371 27523
rect 40313 27483 40371 27489
rect 41414 27480 41420 27532
rect 41472 27520 41478 27532
rect 41601 27523 41659 27529
rect 41601 27520 41613 27523
rect 41472 27492 41613 27520
rect 41472 27480 41478 27492
rect 41601 27489 41613 27492
rect 41647 27489 41659 27523
rect 41601 27483 41659 27489
rect 43257 27523 43315 27529
rect 43257 27489 43269 27523
rect 43303 27520 43315 27523
rect 43530 27520 43536 27532
rect 43303 27492 43536 27520
rect 43303 27489 43315 27492
rect 43257 27483 43315 27489
rect 43530 27480 43536 27492
rect 43588 27480 43594 27532
rect 44082 27480 44088 27532
rect 44140 27520 44146 27532
rect 44453 27523 44511 27529
rect 44453 27520 44465 27523
rect 44140 27492 44465 27520
rect 44140 27480 44146 27492
rect 44453 27489 44465 27492
rect 44499 27489 44511 27523
rect 44453 27483 44511 27489
rect 45097 27523 45155 27529
rect 45097 27489 45109 27523
rect 45143 27489 45155 27523
rect 45830 27520 45836 27532
rect 45791 27492 45836 27520
rect 45097 27483 45155 27489
rect 39577 27455 39635 27461
rect 37292 27424 39160 27452
rect 34241 27415 34299 27421
rect 30392 27356 31616 27384
rect 31757 27387 31815 27393
rect 28718 27316 28724 27328
rect 25884 27288 27016 27316
rect 28679 27288 28724 27316
rect 28718 27276 28724 27288
rect 28776 27276 28782 27328
rect 29178 27276 29184 27328
rect 29236 27316 29242 27328
rect 30392 27316 30420 27356
rect 31757 27353 31769 27387
rect 31803 27384 31815 27387
rect 36814 27384 36820 27396
rect 31803 27356 36820 27384
rect 31803 27353 31815 27356
rect 31757 27347 31815 27353
rect 36814 27344 36820 27356
rect 36872 27344 36878 27396
rect 39022 27384 39028 27396
rect 38983 27356 39028 27384
rect 39022 27344 39028 27356
rect 39080 27344 39086 27396
rect 39132 27384 39160 27424
rect 39577 27421 39589 27455
rect 39623 27452 39635 27455
rect 39758 27452 39764 27464
rect 39623 27424 39764 27452
rect 39623 27421 39635 27424
rect 39577 27415 39635 27421
rect 39758 27412 39764 27424
rect 39816 27412 39822 27464
rect 40129 27387 40187 27393
rect 40129 27384 40141 27387
rect 39132 27356 40141 27384
rect 40129 27353 40141 27356
rect 40175 27353 40187 27387
rect 45112 27384 45140 27483
rect 45830 27480 45836 27492
rect 45888 27480 45894 27532
rect 49510 27480 49516 27532
rect 49568 27520 49574 27532
rect 49789 27523 49847 27529
rect 49789 27520 49801 27523
rect 49568 27492 49801 27520
rect 49568 27480 49574 27492
rect 49789 27489 49801 27492
rect 49835 27489 49847 27523
rect 50430 27520 50436 27532
rect 50391 27492 50436 27520
rect 49789 27483 49847 27489
rect 50430 27480 50436 27492
rect 50488 27480 50494 27532
rect 54386 27480 54392 27532
rect 54444 27520 54450 27532
rect 55125 27523 55183 27529
rect 55125 27520 55137 27523
rect 54444 27492 55137 27520
rect 54444 27480 54450 27492
rect 55125 27489 55137 27492
rect 55171 27489 55183 27523
rect 55125 27483 55183 27489
rect 55861 27523 55919 27529
rect 55861 27489 55873 27523
rect 55907 27489 55919 27523
rect 55861 27483 55919 27489
rect 55876 27452 55904 27483
rect 56042 27480 56048 27532
rect 56100 27520 56106 27532
rect 56597 27523 56655 27529
rect 56597 27520 56609 27523
rect 56100 27492 56609 27520
rect 56100 27480 56106 27492
rect 56597 27489 56609 27492
rect 56643 27489 56655 27523
rect 56597 27483 56655 27489
rect 55140 27424 55904 27452
rect 55140 27396 55168 27424
rect 40129 27347 40187 27353
rect 40328 27356 45140 27384
rect 29236 27288 30420 27316
rect 29236 27276 29242 27288
rect 30466 27276 30472 27328
rect 30524 27316 30530 27328
rect 30561 27319 30619 27325
rect 30561 27316 30573 27319
rect 30524 27288 30573 27316
rect 30524 27276 30530 27288
rect 30561 27285 30573 27288
rect 30607 27285 30619 27319
rect 30561 27279 30619 27285
rect 31202 27276 31208 27328
rect 31260 27316 31266 27328
rect 33689 27319 33747 27325
rect 33689 27316 33701 27319
rect 31260 27288 33701 27316
rect 31260 27276 31266 27288
rect 33689 27285 33701 27288
rect 33735 27285 33747 27319
rect 34882 27316 34888 27328
rect 34843 27288 34888 27316
rect 33689 27279 33747 27285
rect 34882 27276 34888 27288
rect 34940 27276 34946 27328
rect 37553 27319 37611 27325
rect 37553 27285 37565 27319
rect 37599 27316 37611 27319
rect 38470 27316 38476 27328
rect 37599 27288 38476 27316
rect 37599 27285 37611 27288
rect 37553 27279 37611 27285
rect 38470 27276 38476 27288
rect 38528 27276 38534 27328
rect 39114 27276 39120 27328
rect 39172 27316 39178 27328
rect 40328 27316 40356 27356
rect 55122 27344 55128 27396
rect 55180 27344 55186 27396
rect 41782 27316 41788 27328
rect 39172 27288 40356 27316
rect 41743 27288 41788 27316
rect 39172 27276 39178 27288
rect 41782 27276 41788 27288
rect 41840 27276 41846 27328
rect 48406 27316 48412 27328
rect 48367 27288 48412 27316
rect 48406 27276 48412 27288
rect 48464 27276 48470 27328
rect 51166 27316 51172 27328
rect 51127 27288 51172 27316
rect 51166 27276 51172 27288
rect 51224 27276 51230 27328
rect 52362 27316 52368 27328
rect 52323 27288 52368 27316
rect 52362 27276 52368 27288
rect 52420 27276 52426 27328
rect 53466 27316 53472 27328
rect 53427 27288 53472 27316
rect 53466 27276 53472 27288
rect 53524 27276 53530 27328
rect 57606 27276 57612 27328
rect 57664 27316 57670 27328
rect 57793 27319 57851 27325
rect 57793 27316 57805 27319
rect 57664 27288 57805 27316
rect 57664 27276 57670 27288
rect 57793 27285 57805 27288
rect 57839 27285 57851 27319
rect 57793 27279 57851 27285
rect 1104 27226 58880 27248
rect 1104 27174 10614 27226
rect 10666 27174 10678 27226
rect 10730 27174 10742 27226
rect 10794 27174 10806 27226
rect 10858 27174 29878 27226
rect 29930 27174 29942 27226
rect 29994 27174 30006 27226
rect 30058 27174 30070 27226
rect 30122 27174 49142 27226
rect 49194 27174 49206 27226
rect 49258 27174 49270 27226
rect 49322 27174 49334 27226
rect 49386 27174 58880 27226
rect 1104 27152 58880 27174
rect 19978 27072 19984 27124
rect 20036 27112 20042 27124
rect 20530 27112 20536 27124
rect 20036 27084 20536 27112
rect 20036 27072 20042 27084
rect 20530 27072 20536 27084
rect 20588 27072 20594 27124
rect 23293 27115 23351 27121
rect 23293 27081 23305 27115
rect 23339 27112 23351 27115
rect 24118 27112 24124 27124
rect 23339 27084 24124 27112
rect 23339 27081 23351 27084
rect 23293 27075 23351 27081
rect 24118 27072 24124 27084
rect 24176 27072 24182 27124
rect 25866 27072 25872 27124
rect 25924 27112 25930 27124
rect 30190 27112 30196 27124
rect 25924 27084 30196 27112
rect 25924 27072 25930 27084
rect 30190 27072 30196 27084
rect 30248 27072 30254 27124
rect 30282 27072 30288 27124
rect 30340 27112 30346 27124
rect 30340 27084 35756 27112
rect 30340 27072 30346 27084
rect 1394 27004 1400 27056
rect 1452 27044 1458 27056
rect 2133 27047 2191 27053
rect 2133 27044 2145 27047
rect 1452 27016 2145 27044
rect 1452 27004 1458 27016
rect 2133 27013 2145 27016
rect 2179 27013 2191 27047
rect 2133 27007 2191 27013
rect 3053 27047 3111 27053
rect 3053 27013 3065 27047
rect 3099 27044 3111 27047
rect 3878 27044 3884 27056
rect 3099 27016 3884 27044
rect 3099 27013 3111 27016
rect 3053 27007 3111 27013
rect 3878 27004 3884 27016
rect 3936 27004 3942 27056
rect 4246 27044 4252 27056
rect 4207 27016 4252 27044
rect 4246 27004 4252 27016
rect 4304 27004 4310 27056
rect 5994 27004 6000 27056
rect 6052 27044 6058 27056
rect 6914 27044 6920 27056
rect 6052 27016 6920 27044
rect 6052 27004 6058 27016
rect 6914 27004 6920 27016
rect 6972 27004 6978 27056
rect 8665 27047 8723 27053
rect 8665 27013 8677 27047
rect 8711 27044 8723 27047
rect 16301 27047 16359 27053
rect 8711 27016 11606 27044
rect 8711 27013 8723 27016
rect 8665 27007 8723 27013
rect 4709 26979 4767 26985
rect 4709 26945 4721 26979
rect 4755 26976 4767 26979
rect 5718 26976 5724 26988
rect 4755 26948 5724 26976
rect 4755 26945 4767 26948
rect 4709 26939 4767 26945
rect 5718 26936 5724 26948
rect 5776 26936 5782 26988
rect 6454 26936 6460 26988
rect 6512 26976 6518 26988
rect 6825 26979 6883 26985
rect 6825 26976 6837 26979
rect 6512 26948 6837 26976
rect 6512 26936 6518 26948
rect 6825 26945 6837 26948
rect 6871 26945 6883 26979
rect 8110 26976 8116 26988
rect 6825 26939 6883 26945
rect 7024 26948 8116 26976
rect 1486 26908 1492 26920
rect 1447 26880 1492 26908
rect 1486 26868 1492 26880
rect 1544 26868 1550 26920
rect 2866 26908 2872 26920
rect 2827 26880 2872 26908
rect 2866 26868 2872 26880
rect 2924 26908 2930 26920
rect 3513 26911 3571 26917
rect 3513 26908 3525 26911
rect 2924 26880 3525 26908
rect 2924 26868 2930 26880
rect 3513 26877 3525 26880
rect 3559 26877 3571 26911
rect 3513 26871 3571 26877
rect 4614 26868 4620 26920
rect 4672 26908 4678 26920
rect 7024 26917 7052 26948
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 8846 26936 8852 26988
rect 8904 26976 8910 26988
rect 9309 26979 9367 26985
rect 9309 26976 9321 26979
rect 8904 26948 9321 26976
rect 8904 26936 8910 26948
rect 9309 26945 9321 26948
rect 9355 26976 9367 26979
rect 11238 26976 11244 26988
rect 9355 26948 11244 26976
rect 9355 26945 9367 26948
rect 9309 26939 9367 26945
rect 11238 26936 11244 26948
rect 11296 26936 11302 26988
rect 11578 26976 11606 27016
rect 16301 27013 16313 27047
rect 16347 27044 16359 27047
rect 16942 27044 16948 27056
rect 16347 27016 16948 27044
rect 16347 27013 16359 27016
rect 16301 27007 16359 27013
rect 16942 27004 16948 27016
rect 17000 27044 17006 27056
rect 17678 27044 17684 27056
rect 17000 27016 17684 27044
rect 17000 27004 17006 27016
rect 17678 27004 17684 27016
rect 17736 27004 17742 27056
rect 17954 27044 17960 27056
rect 17915 27016 17960 27044
rect 17954 27004 17960 27016
rect 18012 27004 18018 27056
rect 22278 27044 22284 27056
rect 18064 27016 22284 27044
rect 18064 26976 18092 27016
rect 22278 27004 22284 27016
rect 22336 27004 22342 27056
rect 22554 27044 22560 27056
rect 22515 27016 22560 27044
rect 22554 27004 22560 27016
rect 22612 27004 22618 27056
rect 26881 27047 26939 27053
rect 24228 27016 26832 27044
rect 11578 26948 18092 26976
rect 19061 26979 19119 26985
rect 19061 26945 19073 26979
rect 19107 26976 19119 26979
rect 24228 26976 24256 27016
rect 19107 26948 24256 26976
rect 19107 26945 19119 26948
rect 19061 26939 19119 26945
rect 5537 26911 5595 26917
rect 5537 26908 5549 26911
rect 4672 26880 5549 26908
rect 4672 26868 4678 26880
rect 5537 26877 5549 26880
rect 5583 26877 5595 26911
rect 5537 26871 5595 26877
rect 7009 26911 7067 26917
rect 7009 26877 7021 26911
rect 7055 26877 7067 26911
rect 7009 26871 7067 26877
rect 7374 26868 7380 26920
rect 7432 26908 7438 26920
rect 7561 26911 7619 26917
rect 7561 26908 7573 26911
rect 7432 26880 7573 26908
rect 7432 26868 7438 26880
rect 7561 26877 7573 26880
rect 7607 26877 7619 26911
rect 7561 26871 7619 26877
rect 8481 26911 8539 26917
rect 8481 26877 8493 26911
rect 8527 26908 8539 26911
rect 8754 26908 8760 26920
rect 8527 26880 8760 26908
rect 8527 26877 8539 26880
rect 8481 26871 8539 26877
rect 8754 26868 8760 26880
rect 8812 26868 8818 26920
rect 9398 26908 9404 26920
rect 9359 26880 9404 26908
rect 9398 26868 9404 26880
rect 9456 26868 9462 26920
rect 10318 26868 10324 26920
rect 10376 26908 10382 26920
rect 10597 26911 10655 26917
rect 10597 26908 10609 26911
rect 10376 26880 10609 26908
rect 10376 26868 10382 26880
rect 10597 26877 10609 26880
rect 10643 26877 10655 26911
rect 10597 26871 10655 26877
rect 11149 26911 11207 26917
rect 11149 26877 11161 26911
rect 11195 26877 11207 26911
rect 11149 26871 11207 26877
rect 1670 26840 1676 26852
rect 1631 26812 1676 26840
rect 1670 26800 1676 26812
rect 1728 26800 1734 26852
rect 2317 26843 2375 26849
rect 2317 26809 2329 26843
rect 2363 26840 2375 26843
rect 3326 26840 3332 26852
rect 2363 26812 3332 26840
rect 2363 26809 2375 26812
rect 2317 26803 2375 26809
rect 3326 26800 3332 26812
rect 3384 26800 3390 26852
rect 4801 26843 4859 26849
rect 4801 26809 4813 26843
rect 4847 26840 4859 26843
rect 4890 26840 4896 26852
rect 4847 26812 4896 26840
rect 4847 26809 4859 26812
rect 4801 26803 4859 26809
rect 4890 26800 4896 26812
rect 4948 26800 4954 26852
rect 7926 26800 7932 26852
rect 7984 26840 7990 26852
rect 9493 26843 9551 26849
rect 9493 26840 9505 26843
rect 7984 26812 9505 26840
rect 7984 26800 7990 26812
rect 9493 26809 9505 26812
rect 9539 26809 9551 26843
rect 11164 26840 11192 26871
rect 11974 26868 11980 26920
rect 12032 26908 12038 26920
rect 12069 26911 12127 26917
rect 12069 26908 12081 26911
rect 12032 26880 12081 26908
rect 12032 26868 12038 26880
rect 12069 26877 12081 26880
rect 12115 26877 12127 26911
rect 12894 26908 12900 26920
rect 12855 26880 12900 26908
rect 12069 26871 12127 26877
rect 12894 26868 12900 26880
rect 12952 26908 12958 26920
rect 13541 26911 13599 26917
rect 13541 26908 13553 26911
rect 12952 26880 13553 26908
rect 12952 26868 12958 26880
rect 13541 26877 13553 26880
rect 13587 26877 13599 26911
rect 14274 26908 14280 26920
rect 14235 26880 14280 26908
rect 13541 26871 13599 26877
rect 14274 26868 14280 26880
rect 14332 26908 14338 26920
rect 14921 26911 14979 26917
rect 14921 26908 14933 26911
rect 14332 26880 14933 26908
rect 14332 26868 14338 26880
rect 14921 26877 14933 26880
rect 14967 26877 14979 26911
rect 14921 26871 14979 26877
rect 15654 26868 15660 26920
rect 15712 26908 15718 26920
rect 15749 26911 15807 26917
rect 15749 26908 15761 26911
rect 15712 26880 15761 26908
rect 15712 26868 15718 26880
rect 15749 26877 15761 26880
rect 15795 26877 15807 26911
rect 16390 26908 16396 26920
rect 16351 26880 16396 26908
rect 15749 26871 15807 26877
rect 16390 26868 16396 26880
rect 16448 26868 16454 26920
rect 16758 26868 16764 26920
rect 16816 26908 16822 26920
rect 17405 26911 17463 26917
rect 17405 26908 17417 26911
rect 16816 26880 17417 26908
rect 16816 26868 16822 26880
rect 17405 26877 17417 26880
rect 17451 26908 17463 26911
rect 19076 26908 19104 26939
rect 24302 26936 24308 26988
rect 24360 26976 24366 26988
rect 26053 26979 26111 26985
rect 26053 26976 26065 26979
rect 24360 26948 26065 26976
rect 24360 26936 24366 26948
rect 26053 26945 26065 26948
rect 26099 26945 26111 26979
rect 26804 26976 26832 27016
rect 26881 27013 26893 27047
rect 26927 27044 26939 27047
rect 27154 27044 27160 27056
rect 26927 27016 27160 27044
rect 26927 27013 26939 27016
rect 26881 27007 26939 27013
rect 27154 27004 27160 27016
rect 27212 27004 27218 27056
rect 28994 27044 29000 27056
rect 28955 27016 29000 27044
rect 28994 27004 29000 27016
rect 29052 27004 29058 27056
rect 29546 27044 29552 27056
rect 29507 27016 29552 27044
rect 29546 27004 29552 27016
rect 29604 27004 29610 27056
rect 30834 27044 30840 27056
rect 30795 27016 30840 27044
rect 30834 27004 30840 27016
rect 30892 27004 30898 27056
rect 33336 27016 35664 27044
rect 29454 26976 29460 26988
rect 26804 26948 29460 26976
rect 26053 26939 26111 26945
rect 29454 26936 29460 26948
rect 29512 26976 29518 26988
rect 30009 26979 30067 26985
rect 29512 26948 29638 26976
rect 29512 26936 29518 26948
rect 17451 26880 19104 26908
rect 19260 26880 20024 26908
rect 17451 26877 17463 26880
rect 17405 26871 17463 26877
rect 17494 26840 17500 26852
rect 11164 26812 12940 26840
rect 9493 26803 9551 26809
rect 12912 26784 12940 26812
rect 13096 26812 16436 26840
rect 17455 26812 17500 26840
rect 4709 26775 4767 26781
rect 4709 26741 4721 26775
rect 4755 26772 4767 26775
rect 5353 26775 5411 26781
rect 5353 26772 5365 26775
rect 4755 26744 5365 26772
rect 4755 26741 4767 26744
rect 4709 26735 4767 26741
rect 5353 26741 5365 26744
rect 5399 26741 5411 26775
rect 5353 26735 5411 26741
rect 7745 26775 7803 26781
rect 7745 26741 7757 26775
rect 7791 26772 7803 26775
rect 8018 26772 8024 26784
rect 7791 26744 8024 26772
rect 7791 26741 7803 26744
rect 7745 26735 7803 26741
rect 8018 26732 8024 26744
rect 8076 26732 8082 26784
rect 9674 26732 9680 26784
rect 9732 26772 9738 26784
rect 9861 26775 9919 26781
rect 9861 26772 9873 26775
rect 9732 26744 9873 26772
rect 9732 26732 9738 26744
rect 9861 26741 9873 26744
rect 9907 26741 9919 26775
rect 11054 26772 11060 26784
rect 11015 26744 11060 26772
rect 9861 26735 9919 26741
rect 11054 26732 11060 26744
rect 11112 26732 11118 26784
rect 12250 26772 12256 26784
rect 12211 26744 12256 26772
rect 12250 26732 12256 26744
rect 12308 26732 12314 26784
rect 12894 26732 12900 26784
rect 12952 26732 12958 26784
rect 13096 26781 13124 26812
rect 13081 26775 13139 26781
rect 13081 26741 13093 26775
rect 13127 26741 13139 26775
rect 14458 26772 14464 26784
rect 14419 26744 14464 26772
rect 13081 26735 13139 26741
rect 14458 26732 14464 26744
rect 14516 26732 14522 26784
rect 15562 26772 15568 26784
rect 15523 26744 15568 26772
rect 15562 26732 15568 26744
rect 15620 26732 15626 26784
rect 16408 26772 16436 26812
rect 17494 26800 17500 26812
rect 17552 26800 17558 26852
rect 17678 26840 17684 26852
rect 17639 26812 17684 26840
rect 17678 26800 17684 26812
rect 17736 26800 17742 26852
rect 18046 26800 18052 26852
rect 18104 26840 18110 26852
rect 19058 26840 19064 26852
rect 18104 26812 19064 26840
rect 18104 26800 18110 26812
rect 19058 26800 19064 26812
rect 19116 26840 19122 26852
rect 19260 26840 19288 26880
rect 19116 26812 19288 26840
rect 19996 26840 20024 26880
rect 20438 26868 20444 26920
rect 20496 26908 20502 26920
rect 20533 26911 20591 26917
rect 20533 26908 20545 26911
rect 20496 26880 20545 26908
rect 20496 26868 20502 26880
rect 20533 26877 20545 26880
rect 20579 26877 20591 26911
rect 21082 26908 21088 26920
rect 21043 26880 21088 26908
rect 20533 26871 20591 26877
rect 21082 26868 21088 26880
rect 21140 26868 21146 26920
rect 22830 26868 22836 26920
rect 22888 26908 22894 26920
rect 23293 26911 23351 26917
rect 23293 26908 23305 26911
rect 22888 26880 23305 26908
rect 22888 26868 22894 26880
rect 23293 26877 23305 26880
rect 23339 26877 23351 26911
rect 23293 26871 23351 26877
rect 23477 26911 23535 26917
rect 23477 26877 23489 26911
rect 23523 26877 23535 26911
rect 23477 26871 23535 26877
rect 20254 26840 20260 26852
rect 19996 26812 20260 26840
rect 19116 26800 19122 26812
rect 20254 26800 20260 26812
rect 20312 26840 20318 26852
rect 21545 26843 21603 26849
rect 21545 26840 21557 26843
rect 20312 26812 21557 26840
rect 20312 26800 20318 26812
rect 21545 26809 21557 26812
rect 21591 26809 21603 26843
rect 22738 26840 22744 26852
rect 22699 26812 22744 26840
rect 21545 26803 21603 26809
rect 22738 26800 22744 26812
rect 22796 26800 22802 26852
rect 23198 26800 23204 26852
rect 23256 26840 23262 26852
rect 23492 26840 23520 26871
rect 23566 26868 23572 26920
rect 23624 26908 23630 26920
rect 24121 26911 24179 26917
rect 24121 26908 24133 26911
rect 23624 26880 24133 26908
rect 23624 26868 23630 26880
rect 24121 26877 24133 26880
rect 24167 26877 24179 26911
rect 24121 26871 24179 26877
rect 24857 26911 24915 26917
rect 24857 26877 24869 26911
rect 24903 26908 24915 26911
rect 25314 26908 25320 26920
rect 24903 26880 25320 26908
rect 24903 26877 24915 26880
rect 24857 26871 24915 26877
rect 25314 26868 25320 26880
rect 25372 26868 25378 26920
rect 25961 26911 26019 26917
rect 25961 26877 25973 26911
rect 26007 26877 26019 26911
rect 25961 26871 26019 26877
rect 26145 26911 26203 26917
rect 26145 26877 26157 26911
rect 26191 26908 26203 26911
rect 26326 26908 26332 26920
rect 26191 26880 26332 26908
rect 26191 26877 26203 26880
rect 26145 26871 26203 26877
rect 23256 26812 23520 26840
rect 25976 26840 26004 26871
rect 26326 26868 26332 26880
rect 26384 26868 26390 26920
rect 26878 26908 26884 26920
rect 26436 26880 26884 26908
rect 26436 26840 26464 26880
rect 26878 26868 26884 26880
rect 26936 26908 26942 26920
rect 27801 26911 27859 26917
rect 27801 26908 27813 26911
rect 26936 26880 27813 26908
rect 26936 26868 26942 26880
rect 27801 26877 27813 26880
rect 27847 26877 27859 26911
rect 28074 26908 28080 26920
rect 27801 26871 27859 26877
rect 27908 26880 28080 26908
rect 25976 26812 26464 26840
rect 23256 26800 23262 26812
rect 26602 26800 26608 26852
rect 26660 26840 26666 26852
rect 26697 26843 26755 26849
rect 26697 26840 26709 26843
rect 26660 26812 26709 26840
rect 26660 26800 26666 26812
rect 26697 26809 26709 26812
rect 26743 26809 26755 26843
rect 26697 26803 26755 26809
rect 27246 26800 27252 26852
rect 27304 26840 27310 26852
rect 27908 26840 27936 26880
rect 28074 26868 28080 26880
rect 28132 26868 28138 26920
rect 29610 26908 29638 26948
rect 30009 26945 30021 26979
rect 30055 26976 30067 26979
rect 30466 26976 30472 26988
rect 30055 26948 30472 26976
rect 30055 26945 30067 26948
rect 30009 26939 30067 26945
rect 30466 26936 30472 26948
rect 30524 26936 30530 26988
rect 33336 26976 33364 27016
rect 30852 26948 33364 26976
rect 30101 26911 30159 26917
rect 30101 26908 30113 26911
rect 29610 26880 30113 26908
rect 30101 26877 30113 26880
rect 30147 26877 30159 26911
rect 30101 26871 30159 26877
rect 28166 26840 28172 26852
rect 27304 26812 27936 26840
rect 28127 26812 28172 26840
rect 27304 26800 27310 26812
rect 28166 26800 28172 26812
rect 28224 26800 28230 26852
rect 28350 26800 28356 26852
rect 28408 26840 28414 26852
rect 28813 26843 28871 26849
rect 28813 26840 28825 26843
rect 28408 26812 28825 26840
rect 28408 26800 28414 26812
rect 28813 26809 28825 26812
rect 28859 26809 28871 26843
rect 28813 26803 28871 26809
rect 30009 26843 30067 26849
rect 30009 26809 30021 26843
rect 30055 26840 30067 26843
rect 30852 26840 30880 26948
rect 33410 26936 33416 26988
rect 33468 26976 33474 26988
rect 33505 26979 33563 26985
rect 33505 26976 33517 26979
rect 33468 26948 33517 26976
rect 33468 26936 33474 26948
rect 33505 26945 33517 26948
rect 33551 26945 33563 26979
rect 33505 26939 33563 26945
rect 33597 26979 33655 26985
rect 33597 26945 33609 26979
rect 33643 26945 33655 26979
rect 33597 26939 33655 26945
rect 31754 26868 31760 26920
rect 31812 26908 31818 26920
rect 31941 26911 31999 26917
rect 31941 26908 31953 26911
rect 31812 26880 31953 26908
rect 31812 26868 31818 26880
rect 31941 26877 31953 26880
rect 31987 26877 31999 26911
rect 31941 26871 31999 26877
rect 31018 26840 31024 26852
rect 30055 26812 30880 26840
rect 30979 26812 31024 26840
rect 30055 26809 30067 26812
rect 30009 26803 30067 26809
rect 31018 26800 31024 26812
rect 31076 26800 31082 26852
rect 32582 26800 32588 26852
rect 32640 26840 32646 26852
rect 33413 26843 33471 26849
rect 33413 26840 33425 26843
rect 32640 26812 33425 26840
rect 32640 26800 32646 26812
rect 33413 26809 33425 26812
rect 33459 26809 33471 26843
rect 33612 26840 33640 26939
rect 33870 26868 33876 26920
rect 33928 26908 33934 26920
rect 34425 26911 34483 26917
rect 34425 26908 34437 26911
rect 33928 26880 34437 26908
rect 33928 26868 33934 26880
rect 34425 26877 34437 26880
rect 34471 26877 34483 26911
rect 34698 26908 34704 26920
rect 34659 26880 34704 26908
rect 34425 26871 34483 26877
rect 34698 26868 34704 26880
rect 34756 26868 34762 26920
rect 35529 26911 35587 26917
rect 35529 26877 35541 26911
rect 35575 26877 35587 26911
rect 35529 26871 35587 26877
rect 33413 26803 33471 26809
rect 33520 26812 33640 26840
rect 33520 26784 33548 26812
rect 19245 26775 19303 26781
rect 19245 26772 19257 26775
rect 16408 26744 19257 26772
rect 19245 26741 19257 26744
rect 19291 26741 19303 26775
rect 19245 26735 19303 26741
rect 19337 26775 19395 26781
rect 19337 26741 19349 26775
rect 19383 26772 19395 26775
rect 19610 26772 19616 26784
rect 19383 26744 19616 26772
rect 19383 26741 19395 26744
rect 19337 26735 19395 26741
rect 19610 26732 19616 26744
rect 19668 26732 19674 26784
rect 19705 26775 19763 26781
rect 19705 26741 19717 26775
rect 19751 26772 19763 26775
rect 20714 26772 20720 26784
rect 19751 26744 20720 26772
rect 19751 26741 19763 26744
rect 19705 26735 19763 26741
rect 20714 26732 20720 26744
rect 20772 26732 20778 26784
rect 20990 26772 20996 26784
rect 20951 26744 20996 26772
rect 20990 26732 20996 26744
rect 21048 26732 21054 26784
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 23937 26775 23995 26781
rect 23937 26772 23949 26775
rect 23624 26744 23949 26772
rect 23624 26732 23630 26744
rect 23937 26741 23949 26744
rect 23983 26741 23995 26775
rect 23937 26735 23995 26741
rect 25501 26775 25559 26781
rect 25501 26741 25513 26775
rect 25547 26772 25559 26775
rect 25958 26772 25964 26784
rect 25547 26744 25964 26772
rect 25547 26741 25559 26744
rect 25501 26735 25559 26741
rect 25958 26732 25964 26744
rect 26016 26732 26022 26784
rect 30926 26732 30932 26784
rect 30984 26772 30990 26784
rect 31757 26775 31815 26781
rect 31757 26772 31769 26775
rect 30984 26744 31769 26772
rect 30984 26732 30990 26744
rect 31757 26741 31769 26744
rect 31803 26741 31815 26775
rect 31757 26735 31815 26741
rect 33045 26775 33103 26781
rect 33045 26741 33057 26775
rect 33091 26772 33103 26775
rect 33318 26772 33324 26784
rect 33091 26744 33324 26772
rect 33091 26741 33103 26744
rect 33045 26735 33103 26741
rect 33318 26732 33324 26744
rect 33376 26732 33382 26784
rect 33502 26732 33508 26784
rect 33560 26732 33566 26784
rect 34514 26772 34520 26784
rect 34475 26744 34520 26772
rect 34514 26732 34520 26744
rect 34572 26732 34578 26784
rect 35544 26772 35572 26871
rect 35636 26840 35664 27016
rect 35728 26985 35756 27084
rect 48314 27072 48320 27124
rect 48372 27112 48378 27124
rect 48685 27115 48743 27121
rect 48685 27112 48697 27115
rect 48372 27084 48697 27112
rect 48372 27072 48378 27084
rect 48685 27081 48697 27084
rect 48731 27081 48743 27115
rect 48685 27075 48743 27081
rect 51994 27072 52000 27124
rect 52052 27112 52058 27124
rect 52089 27115 52147 27121
rect 52089 27112 52101 27115
rect 52052 27084 52101 27112
rect 52052 27072 52058 27084
rect 52089 27081 52101 27084
rect 52135 27081 52147 27115
rect 52089 27075 52147 27081
rect 53374 27072 53380 27124
rect 53432 27112 53438 27124
rect 53745 27115 53803 27121
rect 53745 27112 53757 27115
rect 53432 27084 53757 27112
rect 53432 27072 53438 27084
rect 53745 27081 53757 27084
rect 53791 27081 53803 27115
rect 53745 27075 53803 27081
rect 38473 27047 38531 27053
rect 38473 27013 38485 27047
rect 38519 27044 38531 27047
rect 39298 27044 39304 27056
rect 38519 27016 39304 27044
rect 38519 27013 38531 27016
rect 38473 27007 38531 27013
rect 39298 27004 39304 27016
rect 39356 27004 39362 27056
rect 39850 27004 39856 27056
rect 39908 27044 39914 27056
rect 40405 27047 40463 27053
rect 40405 27044 40417 27047
rect 39908 27016 40417 27044
rect 39908 27004 39914 27016
rect 40405 27013 40417 27016
rect 40451 27013 40463 27047
rect 41874 27044 41880 27056
rect 41835 27016 41880 27044
rect 40405 27007 40463 27013
rect 41874 27004 41880 27016
rect 41932 27004 41938 27056
rect 44082 27044 44088 27056
rect 44043 27016 44088 27044
rect 44082 27004 44088 27016
rect 44140 27004 44146 27056
rect 44634 27044 44640 27056
rect 44595 27016 44640 27044
rect 44634 27004 44640 27016
rect 44692 27004 44698 27056
rect 45370 27044 45376 27056
rect 45331 27016 45376 27044
rect 45370 27004 45376 27016
rect 45428 27004 45434 27056
rect 47854 27044 47860 27056
rect 47815 27016 47860 27044
rect 47854 27004 47860 27016
rect 47912 27004 47918 27056
rect 49694 27044 49700 27056
rect 49655 27016 49700 27044
rect 49694 27004 49700 27016
rect 49752 27004 49758 27056
rect 50154 27044 50160 27056
rect 50115 27016 50160 27044
rect 50154 27004 50160 27016
rect 50212 27004 50218 27056
rect 51074 27044 51080 27056
rect 51035 27016 51080 27044
rect 51074 27004 51080 27016
rect 51132 27004 51138 27056
rect 56134 27044 56140 27056
rect 56095 27016 56140 27044
rect 56134 27004 56140 27016
rect 56192 27004 56198 27056
rect 57425 27047 57483 27053
rect 57425 27013 57437 27047
rect 57471 27044 57483 27047
rect 57514 27044 57520 27056
rect 57471 27016 57520 27044
rect 57471 27013 57483 27016
rect 57425 27007 57483 27013
rect 57514 27004 57520 27016
rect 57572 27004 57578 27056
rect 35713 26979 35771 26985
rect 35713 26945 35725 26979
rect 35759 26945 35771 26979
rect 35713 26939 35771 26945
rect 39577 26979 39635 26985
rect 39577 26945 39589 26979
rect 39623 26976 39635 26979
rect 41690 26976 41696 26988
rect 39623 26948 41696 26976
rect 39623 26945 39635 26948
rect 39577 26939 39635 26945
rect 41690 26936 41696 26948
rect 41748 26936 41754 26988
rect 55033 26979 55091 26985
rect 41800 26948 50384 26976
rect 35802 26908 35808 26920
rect 35715 26880 35808 26908
rect 35802 26868 35808 26880
rect 35860 26908 35866 26920
rect 36541 26911 36599 26917
rect 36541 26908 36553 26911
rect 35860 26880 36553 26908
rect 35860 26868 35866 26880
rect 36541 26877 36553 26880
rect 36587 26877 36599 26911
rect 36722 26908 36728 26920
rect 36683 26880 36728 26908
rect 36541 26871 36599 26877
rect 36722 26868 36728 26880
rect 36780 26868 36786 26920
rect 37369 26911 37427 26917
rect 37369 26877 37381 26911
rect 37415 26908 37427 26911
rect 38289 26911 38347 26917
rect 38289 26908 38301 26911
rect 37415 26880 38301 26908
rect 37415 26877 37427 26880
rect 37369 26871 37427 26877
rect 38289 26877 38301 26880
rect 38335 26908 38347 26911
rect 38654 26908 38660 26920
rect 38335 26880 38660 26908
rect 38335 26877 38347 26880
rect 38289 26871 38347 26877
rect 38654 26868 38660 26880
rect 38712 26868 38718 26920
rect 39850 26908 39856 26920
rect 39811 26880 39856 26908
rect 39850 26868 39856 26880
rect 39908 26868 39914 26920
rect 40034 26868 40040 26920
rect 40092 26908 40098 26920
rect 40954 26908 40960 26920
rect 40092 26880 40960 26908
rect 40092 26868 40098 26880
rect 40954 26868 40960 26880
rect 41012 26908 41018 26920
rect 41141 26911 41199 26917
rect 41141 26908 41153 26911
rect 41012 26880 41153 26908
rect 41012 26868 41018 26880
rect 41141 26877 41153 26880
rect 41187 26877 41199 26911
rect 41141 26871 41199 26877
rect 36262 26840 36268 26852
rect 35636 26812 36268 26840
rect 36262 26800 36268 26812
rect 36320 26800 36326 26852
rect 40586 26840 40592 26852
rect 36740 26812 38654 26840
rect 40547 26812 40592 26840
rect 36170 26772 36176 26784
rect 35544 26744 36176 26772
rect 36170 26732 36176 26744
rect 36228 26732 36234 26784
rect 36740 26781 36768 26812
rect 36725 26775 36783 26781
rect 36725 26741 36737 26775
rect 36771 26741 36783 26775
rect 38626 26772 38654 26812
rect 40586 26800 40592 26812
rect 40644 26800 40650 26852
rect 41800 26840 41828 26948
rect 41874 26868 41880 26920
rect 41932 26908 41938 26920
rect 43165 26911 43223 26917
rect 43165 26908 43177 26911
rect 41932 26880 43177 26908
rect 41932 26868 41938 26880
rect 43165 26877 43177 26880
rect 43211 26877 43223 26911
rect 43165 26871 43223 26877
rect 45094 26868 45100 26920
rect 45152 26908 45158 26920
rect 50356 26917 50384 26948
rect 55033 26945 55045 26979
rect 55079 26976 55091 26979
rect 59354 26976 59360 26988
rect 55079 26948 59360 26976
rect 55079 26945 55091 26948
rect 55033 26939 55091 26945
rect 45557 26911 45615 26917
rect 45557 26908 45569 26911
rect 45152 26880 45569 26908
rect 45152 26868 45158 26880
rect 45557 26877 45569 26880
rect 45603 26908 45615 26911
rect 46017 26911 46075 26917
rect 46017 26908 46029 26911
rect 45603 26880 46029 26908
rect 45603 26877 45615 26880
rect 45557 26871 45615 26877
rect 46017 26877 46029 26880
rect 46063 26877 46075 26911
rect 46017 26871 46075 26877
rect 50341 26911 50399 26917
rect 50341 26877 50353 26911
rect 50387 26877 50399 26911
rect 54386 26908 54392 26920
rect 54347 26880 54392 26908
rect 50341 26871 50399 26877
rect 54386 26868 54392 26880
rect 54444 26868 54450 26920
rect 55692 26917 55720 26948
rect 59354 26936 59360 26948
rect 59412 26936 59418 26988
rect 55677 26911 55735 26917
rect 55677 26877 55689 26911
rect 55723 26877 55735 26911
rect 57241 26911 57299 26917
rect 57241 26908 57253 26911
rect 55677 26871 55735 26877
rect 55784 26880 57253 26908
rect 41156 26812 41828 26840
rect 42061 26843 42119 26849
rect 41156 26772 41184 26812
rect 42061 26809 42073 26843
rect 42107 26840 42119 26843
rect 42334 26840 42340 26852
rect 42107 26812 42340 26840
rect 42107 26809 42119 26812
rect 42061 26803 42119 26809
rect 42334 26800 42340 26812
rect 42392 26800 42398 26852
rect 44450 26800 44456 26852
rect 44508 26840 44514 26852
rect 44821 26843 44879 26849
rect 44821 26840 44833 26843
rect 44508 26812 44833 26840
rect 44508 26800 44514 26812
rect 44821 26809 44833 26812
rect 44867 26809 44879 26843
rect 44821 26803 44879 26809
rect 47673 26843 47731 26849
rect 47673 26809 47685 26843
rect 47719 26840 47731 26843
rect 47762 26840 47768 26852
rect 47719 26812 47768 26840
rect 47719 26809 47731 26812
rect 47673 26803 47731 26809
rect 47762 26800 47768 26812
rect 47820 26800 47826 26852
rect 49513 26843 49571 26849
rect 49513 26809 49525 26843
rect 49559 26840 49571 26843
rect 49970 26840 49976 26852
rect 49559 26812 49976 26840
rect 49559 26809 49571 26812
rect 49513 26803 49571 26809
rect 49970 26800 49976 26812
rect 50028 26800 50034 26852
rect 51261 26843 51319 26849
rect 51261 26809 51273 26843
rect 51307 26809 51319 26843
rect 51261 26803 51319 26809
rect 41322 26772 41328 26784
rect 38626 26744 41184 26772
rect 41283 26744 41328 26772
rect 36725 26735 36783 26741
rect 41322 26732 41328 26744
rect 41380 26732 41386 26784
rect 47854 26732 47860 26784
rect 47912 26772 47918 26784
rect 51276 26772 51304 26803
rect 54662 26800 54668 26852
rect 54720 26840 54726 26852
rect 55784 26840 55812 26880
rect 57241 26877 57253 26880
rect 57287 26877 57299 26911
rect 58066 26908 58072 26920
rect 58027 26880 58072 26908
rect 57241 26871 57299 26877
rect 58066 26868 58072 26880
rect 58124 26868 58130 26920
rect 54720 26812 55812 26840
rect 56321 26843 56379 26849
rect 54720 26800 54726 26812
rect 56321 26809 56333 26843
rect 56367 26809 56379 26843
rect 56321 26803 56379 26809
rect 55490 26772 55496 26784
rect 47912 26744 51304 26772
rect 55451 26744 55496 26772
rect 47912 26732 47918 26744
rect 55490 26732 55496 26744
rect 55548 26732 55554 26784
rect 55674 26732 55680 26784
rect 55732 26772 55738 26784
rect 56336 26772 56364 26803
rect 57698 26800 57704 26852
rect 57756 26840 57762 26852
rect 57885 26843 57943 26849
rect 57885 26840 57897 26843
rect 57756 26812 57897 26840
rect 57756 26800 57762 26812
rect 57885 26809 57897 26812
rect 57931 26809 57943 26843
rect 57885 26803 57943 26809
rect 55732 26744 56364 26772
rect 55732 26732 55738 26744
rect 1104 26682 58880 26704
rect 1104 26630 20246 26682
rect 20298 26630 20310 26682
rect 20362 26630 20374 26682
rect 20426 26630 20438 26682
rect 20490 26630 39510 26682
rect 39562 26630 39574 26682
rect 39626 26630 39638 26682
rect 39690 26630 39702 26682
rect 39754 26630 58880 26682
rect 1104 26608 58880 26630
rect 1489 26571 1547 26577
rect 1489 26537 1501 26571
rect 1535 26568 1547 26571
rect 2590 26568 2596 26580
rect 1535 26540 2596 26568
rect 1535 26537 1547 26540
rect 1489 26531 1547 26537
rect 2590 26528 2596 26540
rect 2648 26528 2654 26580
rect 4614 26528 4620 26580
rect 4672 26568 4678 26580
rect 5169 26571 5227 26577
rect 5169 26568 5181 26571
rect 4672 26540 5181 26568
rect 4672 26528 4678 26540
rect 5169 26537 5181 26540
rect 5215 26537 5227 26571
rect 5718 26568 5724 26580
rect 5679 26540 5724 26568
rect 5169 26531 5227 26537
rect 5718 26528 5724 26540
rect 5776 26528 5782 26580
rect 7374 26568 7380 26580
rect 7335 26540 7380 26568
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 8021 26571 8079 26577
rect 8021 26537 8033 26571
rect 8067 26568 8079 26571
rect 8110 26568 8116 26580
rect 8067 26540 8116 26568
rect 8067 26537 8079 26540
rect 8021 26531 8079 26537
rect 8110 26528 8116 26540
rect 8168 26528 8174 26580
rect 8573 26571 8631 26577
rect 8573 26537 8585 26571
rect 8619 26568 8631 26571
rect 8754 26568 8760 26580
rect 8619 26540 8760 26568
rect 8619 26537 8631 26540
rect 8573 26531 8631 26537
rect 8754 26528 8760 26540
rect 8812 26528 8818 26580
rect 9766 26528 9772 26580
rect 9824 26568 9830 26580
rect 10318 26568 10324 26580
rect 9824 26540 10324 26568
rect 9824 26528 9830 26540
rect 10318 26528 10324 26540
rect 10376 26528 10382 26580
rect 11701 26571 11759 26577
rect 11701 26537 11713 26571
rect 11747 26568 11759 26571
rect 12345 26571 12403 26577
rect 12345 26568 12357 26571
rect 11747 26540 12357 26568
rect 11747 26537 11759 26540
rect 11701 26531 11759 26537
rect 12345 26537 12357 26540
rect 12391 26537 12403 26571
rect 12345 26531 12403 26537
rect 15654 26528 15660 26580
rect 15712 26568 15718 26580
rect 15841 26571 15899 26577
rect 15841 26568 15853 26571
rect 15712 26540 15853 26568
rect 15712 26528 15718 26540
rect 15841 26537 15853 26540
rect 15887 26537 15899 26571
rect 17034 26568 17040 26580
rect 16995 26540 17040 26568
rect 15841 26531 15899 26537
rect 17034 26528 17040 26540
rect 17092 26528 17098 26580
rect 17126 26528 17132 26580
rect 17184 26568 17190 26580
rect 17681 26571 17739 26577
rect 17681 26568 17693 26571
rect 17184 26540 17693 26568
rect 17184 26528 17190 26540
rect 17681 26537 17693 26540
rect 17727 26537 17739 26571
rect 17681 26531 17739 26537
rect 17770 26528 17776 26580
rect 17828 26568 17834 26580
rect 18966 26568 18972 26580
rect 17828 26540 18972 26568
rect 17828 26528 17834 26540
rect 18966 26528 18972 26540
rect 19024 26528 19030 26580
rect 19996 26540 20622 26568
rect 1578 26500 1584 26512
rect 1539 26472 1584 26500
rect 1578 26460 1584 26472
rect 1636 26460 1642 26512
rect 2222 26460 2228 26512
rect 2280 26500 2286 26512
rect 2961 26503 3019 26509
rect 2961 26500 2973 26503
rect 2280 26472 2973 26500
rect 2280 26460 2286 26472
rect 2961 26469 2973 26472
rect 3007 26469 3019 26503
rect 2961 26463 3019 26469
rect 4154 26460 4160 26512
rect 4212 26500 4218 26512
rect 4249 26503 4307 26509
rect 4249 26500 4261 26503
rect 4212 26472 4261 26500
rect 4212 26460 4218 26472
rect 4249 26469 4261 26472
rect 4295 26469 4307 26503
rect 4430 26500 4436 26512
rect 4391 26472 4436 26500
rect 4249 26463 4307 26469
rect 4430 26460 4436 26472
rect 4488 26460 4494 26512
rect 4522 26460 4528 26512
rect 4580 26500 4586 26512
rect 7926 26500 7932 26512
rect 4580 26472 7932 26500
rect 4580 26460 4586 26472
rect 7926 26460 7932 26472
rect 7984 26460 7990 26512
rect 9214 26460 9220 26512
rect 9272 26500 9278 26512
rect 9493 26503 9551 26509
rect 9493 26500 9505 26503
rect 9272 26472 9505 26500
rect 9272 26460 9278 26472
rect 9493 26469 9505 26472
rect 9539 26469 9551 26503
rect 9674 26500 9680 26512
rect 9635 26472 9680 26500
rect 9493 26463 9551 26469
rect 9674 26460 9680 26472
rect 9732 26460 9738 26512
rect 11238 26460 11244 26512
rect 11296 26500 11302 26512
rect 11793 26503 11851 26509
rect 11793 26500 11805 26503
rect 11296 26472 11805 26500
rect 11296 26460 11302 26472
rect 11793 26469 11805 26472
rect 11839 26500 11851 26503
rect 11839 26472 14412 26500
rect 11839 26469 11851 26472
rect 11793 26463 11851 26469
rect 2314 26432 2320 26444
rect 2275 26404 2320 26432
rect 2314 26392 2320 26404
rect 2372 26392 2378 26444
rect 10226 26432 10232 26444
rect 10187 26404 10232 26432
rect 10226 26392 10232 26404
rect 10284 26392 10290 26444
rect 11146 26392 11152 26444
rect 11204 26432 11210 26444
rect 12529 26435 12587 26441
rect 12529 26432 12541 26435
rect 11204 26404 12541 26432
rect 11204 26392 11210 26404
rect 12529 26401 12541 26404
rect 12575 26432 12587 26435
rect 12989 26435 13047 26441
rect 12989 26432 13001 26435
rect 12575 26404 13001 26432
rect 12575 26401 12587 26404
rect 12529 26395 12587 26401
rect 12989 26401 13001 26404
rect 13035 26401 13047 26435
rect 14384 26432 14412 26472
rect 14458 26460 14464 26512
rect 14516 26500 14522 26512
rect 19996 26500 20024 26540
rect 14516 26472 20024 26500
rect 14516 26460 14522 26472
rect 20070 26460 20076 26512
rect 20128 26500 20134 26512
rect 20257 26503 20315 26509
rect 20257 26500 20269 26503
rect 20128 26472 20269 26500
rect 20128 26460 20134 26472
rect 20257 26469 20269 26472
rect 20303 26469 20315 26503
rect 20594 26500 20622 26540
rect 20714 26528 20720 26580
rect 20772 26568 20778 26580
rect 20772 26540 21404 26568
rect 20772 26528 20778 26540
rect 21174 26500 21180 26512
rect 20594 26472 20760 26500
rect 21135 26472 21180 26500
rect 20257 26463 20315 26469
rect 16758 26432 16764 26444
rect 14384 26404 16764 26432
rect 12989 26395 13047 26401
rect 16758 26392 16764 26404
rect 16816 26392 16822 26444
rect 16942 26432 16948 26444
rect 16903 26404 16948 26432
rect 16942 26392 16948 26404
rect 17000 26392 17006 26444
rect 17129 26435 17187 26441
rect 17129 26401 17141 26435
rect 17175 26401 17187 26435
rect 17129 26395 17187 26401
rect 17681 26435 17739 26441
rect 17681 26401 17693 26435
rect 17727 26432 17739 26435
rect 17770 26432 17776 26444
rect 17727 26404 17776 26432
rect 17727 26401 17739 26404
rect 17681 26395 17739 26401
rect 11701 26367 11759 26373
rect 11701 26333 11713 26367
rect 11747 26333 11759 26367
rect 11701 26327 11759 26333
rect 2501 26299 2559 26305
rect 2501 26265 2513 26299
rect 2547 26296 2559 26299
rect 4430 26296 4436 26308
rect 2547 26268 4436 26296
rect 2547 26265 2559 26268
rect 2501 26259 2559 26265
rect 4430 26256 4436 26268
rect 4488 26256 4494 26308
rect 11716 26296 11744 26327
rect 14182 26296 14188 26308
rect 11716 26268 14188 26296
rect 14182 26256 14188 26268
rect 14240 26256 14246 26308
rect 16485 26299 16543 26305
rect 16485 26265 16497 26299
rect 16531 26296 16543 26299
rect 17144 26296 17172 26395
rect 17770 26392 17776 26404
rect 17828 26392 17834 26444
rect 17957 26435 18015 26441
rect 17957 26401 17969 26435
rect 18003 26401 18015 26435
rect 18874 26432 18880 26444
rect 18835 26404 18880 26432
rect 17957 26395 18015 26401
rect 17862 26324 17868 26376
rect 17920 26364 17926 26376
rect 17972 26364 18000 26395
rect 18874 26392 18880 26404
rect 18932 26432 18938 26444
rect 19613 26435 19671 26441
rect 19613 26432 19625 26435
rect 18932 26404 19625 26432
rect 18932 26392 18938 26404
rect 19613 26401 19625 26404
rect 19659 26401 19671 26435
rect 19613 26395 19671 26401
rect 20441 26435 20499 26441
rect 20441 26401 20453 26435
rect 20487 26432 20499 26435
rect 20732 26432 20760 26472
rect 21174 26460 21180 26472
rect 21232 26460 21238 26512
rect 21376 26509 21404 26540
rect 23474 26528 23480 26580
rect 23532 26568 23538 26580
rect 23753 26571 23811 26577
rect 23753 26568 23765 26571
rect 23532 26540 23765 26568
rect 23532 26528 23538 26540
rect 23753 26537 23765 26540
rect 23799 26537 23811 26571
rect 27982 26568 27988 26580
rect 23753 26531 23811 26537
rect 23860 26540 27988 26568
rect 21361 26503 21419 26509
rect 21361 26469 21373 26503
rect 21407 26469 21419 26503
rect 23860 26500 23888 26540
rect 27982 26528 27988 26540
rect 28040 26528 28046 26580
rect 28074 26528 28080 26580
rect 28132 26568 28138 26580
rect 29457 26571 29515 26577
rect 29457 26568 29469 26571
rect 28132 26540 29469 26568
rect 28132 26528 28138 26540
rect 29457 26537 29469 26540
rect 29503 26537 29515 26571
rect 29457 26531 29515 26537
rect 31754 26528 31760 26580
rect 31812 26568 31818 26580
rect 32033 26571 32091 26577
rect 32033 26568 32045 26571
rect 31812 26540 32045 26568
rect 31812 26528 31818 26540
rect 32033 26537 32045 26540
rect 32079 26537 32091 26571
rect 34146 26568 34152 26580
rect 34107 26540 34152 26568
rect 32033 26531 32091 26537
rect 34146 26528 34152 26540
rect 34204 26528 34210 26580
rect 35802 26568 35808 26580
rect 35763 26540 35808 26568
rect 35802 26528 35808 26540
rect 35860 26528 35866 26580
rect 36262 26528 36268 26580
rect 36320 26568 36326 26580
rect 36357 26571 36415 26577
rect 36357 26568 36369 26571
rect 36320 26540 36369 26568
rect 36320 26528 36326 26540
rect 36357 26537 36369 26540
rect 36403 26537 36415 26571
rect 36357 26531 36415 26537
rect 41414 26528 41420 26580
rect 41472 26568 41478 26580
rect 41601 26571 41659 26577
rect 41601 26568 41613 26571
rect 41472 26540 41613 26568
rect 41472 26528 41478 26540
rect 41601 26537 41613 26540
rect 41647 26537 41659 26571
rect 41601 26531 41659 26537
rect 41690 26528 41696 26580
rect 41748 26568 41754 26580
rect 47394 26568 47400 26580
rect 41748 26540 47400 26568
rect 41748 26528 41754 26540
rect 47394 26528 47400 26540
rect 47452 26528 47458 26580
rect 51534 26528 51540 26580
rect 51592 26568 51598 26580
rect 54662 26568 54668 26580
rect 51592 26540 51637 26568
rect 54623 26540 54668 26568
rect 51592 26528 51598 26540
rect 54662 26528 54668 26540
rect 54720 26528 54726 26580
rect 55769 26571 55827 26577
rect 55769 26537 55781 26571
rect 55815 26568 55827 26571
rect 58066 26568 58072 26580
rect 55815 26540 58072 26568
rect 55815 26537 55827 26540
rect 55769 26531 55827 26537
rect 58066 26528 58072 26540
rect 58124 26528 58130 26580
rect 21361 26463 21419 26469
rect 21468 26472 23888 26500
rect 21468 26432 21496 26472
rect 26326 26460 26332 26512
rect 26384 26500 26390 26512
rect 27065 26503 27123 26509
rect 27065 26500 27077 26503
rect 26384 26472 27077 26500
rect 26384 26460 26390 26472
rect 27065 26469 27077 26472
rect 27111 26469 27123 26503
rect 27614 26500 27620 26512
rect 27575 26472 27620 26500
rect 27065 26463 27123 26469
rect 27614 26460 27620 26472
rect 27672 26460 27678 26512
rect 33134 26500 33140 26512
rect 33095 26472 33140 26500
rect 33134 26460 33140 26472
rect 33192 26460 33198 26512
rect 33318 26500 33324 26512
rect 33279 26472 33324 26500
rect 33318 26460 33324 26472
rect 33376 26460 33382 26512
rect 38746 26500 38752 26512
rect 38707 26472 38752 26500
rect 38746 26460 38752 26472
rect 38804 26460 38810 26512
rect 38841 26503 38899 26509
rect 38841 26469 38853 26503
rect 38887 26500 38899 26503
rect 39390 26500 39396 26512
rect 38887 26472 39396 26500
rect 38887 26469 38899 26472
rect 38841 26463 38899 26469
rect 39390 26460 39396 26472
rect 39448 26500 39454 26512
rect 39850 26500 39856 26512
rect 39448 26472 39856 26500
rect 39448 26460 39454 26472
rect 39850 26460 39856 26472
rect 39908 26500 39914 26512
rect 41874 26500 41880 26512
rect 39908 26472 41880 26500
rect 39908 26460 39914 26472
rect 41874 26460 41880 26472
rect 41932 26460 41938 26512
rect 55122 26500 55128 26512
rect 55083 26472 55128 26500
rect 55122 26460 55128 26472
rect 55180 26460 55186 26512
rect 56594 26460 56600 26512
rect 56652 26500 56658 26512
rect 56689 26503 56747 26509
rect 56689 26500 56701 26503
rect 56652 26472 56701 26500
rect 56652 26460 56658 26472
rect 56689 26469 56701 26472
rect 56735 26469 56747 26503
rect 58158 26500 58164 26512
rect 58119 26472 58164 26500
rect 56689 26463 56747 26469
rect 58158 26460 58164 26472
rect 58216 26460 58222 26512
rect 22278 26432 22284 26444
rect 20487 26404 20622 26432
rect 20732 26404 21496 26432
rect 22239 26404 22284 26432
rect 20487 26401 20499 26404
rect 20441 26395 20499 26401
rect 17920 26336 18000 26364
rect 20594 26364 20622 26404
rect 22278 26392 22284 26404
rect 22336 26392 22342 26444
rect 25869 26435 25927 26441
rect 25869 26401 25881 26435
rect 25915 26432 25927 26435
rect 26513 26435 26571 26441
rect 26513 26432 26525 26435
rect 25915 26404 26525 26432
rect 25915 26401 25927 26404
rect 25869 26395 25927 26401
rect 26513 26401 26525 26404
rect 26559 26432 26571 26435
rect 26694 26432 26700 26444
rect 26559 26404 26700 26432
rect 26559 26401 26571 26404
rect 26513 26395 26571 26401
rect 26694 26392 26700 26404
rect 26752 26392 26758 26444
rect 27157 26435 27215 26441
rect 27157 26401 27169 26435
rect 27203 26401 27215 26435
rect 27798 26432 27804 26444
rect 27759 26404 27804 26432
rect 27157 26395 27215 26401
rect 27172 26364 27200 26395
rect 27798 26392 27804 26404
rect 27856 26392 27862 26444
rect 29273 26435 29331 26441
rect 29273 26401 29285 26435
rect 29319 26432 29331 26435
rect 29525 26435 29583 26441
rect 29525 26432 29537 26435
rect 29319 26404 29537 26432
rect 29319 26401 29331 26404
rect 29273 26395 29331 26401
rect 29525 26401 29537 26404
rect 29571 26401 29583 26435
rect 29525 26395 29583 26401
rect 30374 26392 30380 26444
rect 30432 26432 30438 26444
rect 30653 26435 30711 26441
rect 30653 26432 30665 26435
rect 30432 26404 30665 26432
rect 30432 26392 30438 26404
rect 30653 26401 30665 26404
rect 30699 26432 30711 26435
rect 31113 26435 31171 26441
rect 31113 26432 31125 26435
rect 30699 26404 31125 26432
rect 30699 26401 30711 26404
rect 30653 26395 30711 26401
rect 31113 26401 31125 26404
rect 31159 26401 31171 26435
rect 31113 26395 31171 26401
rect 33965 26435 34023 26441
rect 33965 26401 33977 26435
rect 34011 26432 34023 26435
rect 34054 26432 34060 26444
rect 34011 26404 34060 26432
rect 34011 26401 34023 26404
rect 33965 26395 34023 26401
rect 34054 26392 34060 26404
rect 34112 26392 34118 26444
rect 34330 26392 34336 26444
rect 34388 26432 34394 26444
rect 34609 26435 34667 26441
rect 34609 26432 34621 26435
rect 34388 26404 34621 26432
rect 34388 26392 34394 26404
rect 34609 26401 34621 26404
rect 34655 26401 34667 26435
rect 35710 26432 35716 26444
rect 35671 26404 35716 26432
rect 34609 26395 34667 26401
rect 35710 26392 35716 26404
rect 35768 26392 35774 26444
rect 36354 26392 36360 26444
rect 36412 26432 36418 26444
rect 36541 26435 36599 26441
rect 36541 26432 36553 26435
rect 36412 26404 36553 26432
rect 36412 26392 36418 26404
rect 36541 26401 36553 26404
rect 36587 26401 36599 26435
rect 36541 26395 36599 26401
rect 37274 26392 37280 26444
rect 37332 26432 37338 26444
rect 37369 26435 37427 26441
rect 37369 26432 37381 26435
rect 37332 26404 37381 26432
rect 37332 26392 37338 26404
rect 37369 26401 37381 26404
rect 37415 26401 37427 26435
rect 37369 26395 37427 26401
rect 37458 26392 37464 26444
rect 37516 26432 37522 26444
rect 37553 26435 37611 26441
rect 37553 26432 37565 26435
rect 37516 26404 37565 26432
rect 37516 26392 37522 26404
rect 37553 26401 37565 26404
rect 37599 26401 37611 26435
rect 37553 26395 37611 26401
rect 38194 26392 38200 26444
rect 38252 26432 38258 26444
rect 38562 26432 38568 26444
rect 38252 26404 38568 26432
rect 38252 26392 38258 26404
rect 38562 26392 38568 26404
rect 38620 26432 38626 26444
rect 39577 26435 39635 26441
rect 39577 26432 39589 26435
rect 38620 26404 39589 26432
rect 38620 26392 38626 26404
rect 39577 26401 39589 26404
rect 39623 26401 39635 26435
rect 39577 26395 39635 26401
rect 40494 26392 40500 26444
rect 40552 26432 40558 26444
rect 41138 26432 41144 26444
rect 40552 26404 41144 26432
rect 40552 26392 40558 26404
rect 41138 26392 41144 26404
rect 41196 26392 41202 26444
rect 55030 26392 55036 26444
rect 55088 26432 55094 26444
rect 56873 26435 56931 26441
rect 56873 26432 56885 26435
rect 55088 26404 56885 26432
rect 55088 26392 55094 26404
rect 56873 26401 56885 26404
rect 56919 26401 56931 26435
rect 56873 26395 56931 26401
rect 56962 26392 56968 26444
rect 57020 26432 57026 26444
rect 57977 26435 58035 26441
rect 57977 26432 57989 26435
rect 57020 26404 57989 26432
rect 57020 26392 57026 26404
rect 57977 26401 57989 26404
rect 58023 26401 58035 26435
rect 57977 26395 58035 26401
rect 38654 26364 38660 26376
rect 20594 26336 26464 26364
rect 27172 26336 37780 26364
rect 38615 26336 38660 26364
rect 17920 26324 17926 26336
rect 19886 26296 19892 26308
rect 16531 26268 19892 26296
rect 16531 26265 16543 26268
rect 16485 26259 16543 26265
rect 19886 26256 19892 26268
rect 19944 26256 19950 26308
rect 24486 26256 24492 26308
rect 24544 26296 24550 26308
rect 26329 26299 26387 26305
rect 26329 26296 26341 26299
rect 24544 26268 26341 26296
rect 24544 26256 24550 26268
rect 26329 26265 26341 26268
rect 26375 26265 26387 26299
rect 26436 26296 26464 26336
rect 37642 26296 37648 26308
rect 26436 26268 36492 26296
rect 37603 26268 37648 26296
rect 26329 26259 26387 26265
rect 6362 26228 6368 26240
rect 6323 26200 6368 26228
rect 6362 26188 6368 26200
rect 6420 26188 6426 26240
rect 11241 26231 11299 26237
rect 11241 26197 11253 26231
rect 11287 26228 11299 26231
rect 11514 26228 11520 26240
rect 11287 26200 11520 26228
rect 11287 26197 11299 26200
rect 11241 26191 11299 26197
rect 11514 26188 11520 26200
rect 11572 26188 11578 26240
rect 13538 26228 13544 26240
rect 13499 26200 13544 26228
rect 13538 26188 13544 26200
rect 13596 26188 13602 26240
rect 15010 26188 15016 26240
rect 15068 26228 15074 26240
rect 15289 26231 15347 26237
rect 15289 26228 15301 26231
rect 15068 26200 15301 26228
rect 15068 26188 15074 26200
rect 15289 26197 15301 26200
rect 15335 26197 15347 26231
rect 15289 26191 15347 26197
rect 16942 26188 16948 26240
rect 17000 26228 17006 26240
rect 18046 26228 18052 26240
rect 17000 26200 18052 26228
rect 17000 26188 17006 26200
rect 18046 26188 18052 26200
rect 18104 26188 18110 26240
rect 19061 26231 19119 26237
rect 19061 26197 19073 26231
rect 19107 26228 19119 26231
rect 19518 26228 19524 26240
rect 19107 26200 19524 26228
rect 19107 26197 19119 26200
rect 19061 26191 19119 26197
rect 19518 26188 19524 26200
rect 19576 26188 19582 26240
rect 22373 26231 22431 26237
rect 22373 26197 22385 26231
rect 22419 26228 22431 26231
rect 22830 26228 22836 26240
rect 22419 26200 22836 26228
rect 22419 26197 22431 26200
rect 22373 26191 22431 26197
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 23198 26228 23204 26240
rect 23159 26200 23204 26228
rect 23198 26188 23204 26200
rect 23256 26188 23262 26240
rect 25317 26231 25375 26237
rect 25317 26197 25329 26231
rect 25363 26228 25375 26231
rect 26878 26228 26884 26240
rect 25363 26200 26884 26228
rect 25363 26197 25375 26200
rect 25317 26191 25375 26197
rect 26878 26188 26884 26200
rect 26936 26228 26942 26240
rect 28353 26231 28411 26237
rect 28353 26228 28365 26231
rect 26936 26200 28365 26228
rect 26936 26188 26942 26200
rect 28353 26197 28365 26200
rect 28399 26197 28411 26231
rect 28353 26191 28411 26197
rect 29273 26231 29331 26237
rect 29273 26197 29285 26231
rect 29319 26228 29331 26231
rect 30469 26231 30527 26237
rect 30469 26228 30481 26231
rect 29319 26200 30481 26228
rect 29319 26197 29331 26200
rect 29273 26191 29331 26197
rect 30469 26197 30481 26200
rect 30515 26197 30527 26231
rect 32582 26228 32588 26240
rect 32543 26200 32588 26228
rect 30469 26191 30527 26197
rect 32582 26188 32588 26200
rect 32640 26188 32646 26240
rect 34698 26228 34704 26240
rect 34659 26200 34704 26228
rect 34698 26188 34704 26200
rect 34756 26188 34762 26240
rect 36464 26228 36492 26268
rect 37642 26256 37648 26268
rect 37700 26256 37706 26308
rect 37752 26296 37780 26336
rect 38654 26324 38660 26336
rect 38712 26324 38718 26376
rect 40586 26324 40592 26376
rect 40644 26364 40650 26376
rect 57238 26364 57244 26376
rect 40644 26336 57244 26364
rect 40644 26324 40650 26336
rect 57238 26324 57244 26336
rect 57296 26324 57302 26376
rect 39393 26299 39451 26305
rect 39393 26296 39405 26299
rect 37752 26268 39405 26296
rect 39393 26265 39405 26268
rect 39439 26265 39451 26299
rect 49418 26296 49424 26308
rect 49379 26268 49424 26296
rect 39393 26259 39451 26265
rect 49418 26256 49424 26268
rect 49476 26256 49482 26308
rect 38289 26231 38347 26237
rect 38289 26228 38301 26231
rect 36464 26200 38301 26228
rect 38289 26197 38301 26200
rect 38335 26197 38347 26231
rect 38289 26191 38347 26197
rect 38838 26188 38844 26240
rect 38896 26228 38902 26240
rect 40957 26231 41015 26237
rect 40957 26228 40969 26231
rect 38896 26200 40969 26228
rect 38896 26188 38902 26200
rect 40957 26197 40969 26200
rect 41003 26197 41015 26231
rect 42334 26228 42340 26240
rect 42295 26200 42340 26228
rect 40957 26191 41015 26197
rect 42334 26188 42340 26200
rect 42392 26188 42398 26240
rect 44450 26228 44456 26240
rect 44411 26200 44456 26228
rect 44450 26188 44456 26200
rect 44508 26188 44514 26240
rect 45830 26228 45836 26240
rect 45791 26200 45836 26228
rect 45830 26188 45836 26200
rect 45888 26188 45894 26240
rect 49970 26228 49976 26240
rect 49931 26200 49976 26228
rect 49970 26188 49976 26200
rect 50028 26188 50034 26240
rect 1104 26138 58880 26160
rect 1104 26086 10614 26138
rect 10666 26086 10678 26138
rect 10730 26086 10742 26138
rect 10794 26086 10806 26138
rect 10858 26086 29878 26138
rect 29930 26086 29942 26138
rect 29994 26086 30006 26138
rect 30058 26086 30070 26138
rect 30122 26086 49142 26138
rect 49194 26086 49206 26138
rect 49258 26086 49270 26138
rect 49322 26086 49334 26138
rect 49386 26086 58880 26138
rect 1104 26064 58880 26086
rect 2314 25984 2320 26036
rect 2372 26024 2378 26036
rect 2593 26027 2651 26033
rect 2593 26024 2605 26027
rect 2372 25996 2605 26024
rect 2372 25984 2378 25996
rect 2593 25993 2605 25996
rect 2639 25993 2651 26027
rect 2593 25987 2651 25993
rect 3234 25984 3240 26036
rect 3292 26024 3298 26036
rect 3421 26027 3479 26033
rect 3421 26024 3433 26027
rect 3292 25996 3433 26024
rect 3292 25984 3298 25996
rect 3421 25993 3433 25996
rect 3467 26024 3479 26027
rect 3510 26024 3516 26036
rect 3467 25996 3516 26024
rect 3467 25993 3479 25996
rect 3421 25987 3479 25993
rect 3510 25984 3516 25996
rect 3568 25984 3574 26036
rect 4430 25984 4436 26036
rect 4488 26024 4494 26036
rect 4488 25996 19472 26024
rect 4488 25984 4494 25996
rect 5166 25956 5172 25968
rect 5127 25928 5172 25956
rect 5166 25916 5172 25928
rect 5224 25916 5230 25968
rect 8757 25959 8815 25965
rect 8757 25925 8769 25959
rect 8803 25956 8815 25959
rect 8846 25956 8852 25968
rect 8803 25928 8852 25956
rect 8803 25925 8815 25928
rect 8757 25919 8815 25925
rect 1394 25888 1400 25900
rect 1355 25860 1400 25888
rect 1394 25848 1400 25860
rect 1452 25848 1458 25900
rect 6362 25848 6368 25900
rect 6420 25888 6426 25900
rect 8772 25888 8800 25919
rect 8846 25916 8852 25928
rect 8904 25916 8910 25968
rect 9309 25959 9367 25965
rect 9309 25925 9321 25959
rect 9355 25956 9367 25959
rect 10226 25956 10232 25968
rect 9355 25928 10232 25956
rect 9355 25925 9367 25928
rect 9309 25919 9367 25925
rect 10226 25916 10232 25928
rect 10284 25916 10290 25968
rect 11057 25959 11115 25965
rect 11057 25925 11069 25959
rect 11103 25956 11115 25959
rect 11238 25956 11244 25968
rect 11103 25928 11244 25956
rect 11103 25925 11115 25928
rect 11057 25919 11115 25925
rect 11238 25916 11244 25928
rect 11296 25916 11302 25968
rect 11793 25959 11851 25965
rect 11793 25925 11805 25959
rect 11839 25956 11851 25959
rect 12894 25956 12900 25968
rect 11839 25928 12900 25956
rect 11839 25925 11851 25928
rect 11793 25919 11851 25925
rect 12894 25916 12900 25928
rect 12952 25916 12958 25968
rect 16390 25916 16396 25968
rect 16448 25956 16454 25968
rect 17497 25959 17555 25965
rect 17497 25956 17509 25959
rect 16448 25928 17509 25956
rect 16448 25916 16454 25928
rect 17497 25925 17509 25928
rect 17543 25925 17555 25959
rect 17497 25919 17555 25925
rect 17678 25916 17684 25968
rect 17736 25916 17742 25968
rect 18325 25959 18383 25965
rect 18325 25925 18337 25959
rect 18371 25956 18383 25959
rect 18598 25956 18604 25968
rect 18371 25928 18604 25956
rect 18371 25925 18383 25928
rect 18325 25919 18383 25925
rect 18598 25916 18604 25928
rect 18656 25916 18662 25968
rect 18877 25959 18935 25965
rect 18877 25925 18889 25959
rect 18923 25956 18935 25959
rect 18966 25956 18972 25968
rect 18923 25928 18972 25956
rect 18923 25925 18935 25928
rect 18877 25919 18935 25925
rect 18966 25916 18972 25928
rect 19024 25916 19030 25968
rect 6420 25860 8800 25888
rect 10505 25891 10563 25897
rect 6420 25848 6454 25860
rect 10505 25857 10517 25891
rect 10551 25888 10563 25891
rect 16942 25888 16948 25900
rect 10551 25860 16948 25888
rect 10551 25857 10563 25860
rect 10505 25851 10563 25857
rect 1581 25823 1639 25829
rect 1581 25789 1593 25823
rect 1627 25820 1639 25823
rect 2498 25820 2504 25832
rect 1627 25792 2504 25820
rect 1627 25789 1639 25792
rect 1581 25783 1639 25789
rect 2498 25780 2504 25792
rect 2556 25780 2562 25832
rect 4890 25780 4896 25832
rect 4948 25820 4954 25832
rect 5629 25823 5687 25829
rect 5629 25820 5641 25823
rect 4948 25792 5641 25820
rect 4948 25780 4954 25792
rect 5629 25789 5641 25792
rect 5675 25820 5687 25823
rect 6426 25820 6454 25848
rect 9766 25820 9772 25832
rect 9824 25829 9830 25832
rect 5675 25792 6454 25820
rect 9733 25792 9772 25820
rect 5675 25789 5687 25792
rect 5629 25783 5687 25789
rect 9766 25780 9772 25792
rect 9824 25783 9833 25829
rect 9953 25823 10011 25829
rect 9953 25789 9965 25823
rect 9999 25820 10011 25823
rect 10520 25820 10548 25851
rect 16942 25848 16948 25860
rect 17000 25848 17006 25900
rect 17037 25891 17095 25897
rect 17037 25857 17049 25891
rect 17083 25888 17095 25891
rect 17696 25888 17724 25916
rect 17083 25860 17724 25888
rect 17083 25857 17095 25860
rect 17037 25851 17095 25857
rect 9999 25792 10548 25820
rect 9999 25789 10011 25792
rect 9953 25783 10011 25789
rect 9824 25780 9830 25783
rect 17586 25780 17592 25832
rect 17644 25820 17650 25832
rect 19444 25829 19472 25996
rect 23198 25984 23204 26036
rect 23256 26024 23262 26036
rect 33870 26024 33876 26036
rect 23256 25996 33876 26024
rect 23256 25984 23262 25996
rect 33870 25984 33876 25996
rect 33928 25984 33934 26036
rect 33965 26027 34023 26033
rect 33965 25993 33977 26027
rect 34011 26024 34023 26027
rect 34054 26024 34060 26036
rect 34011 25996 34060 26024
rect 34011 25993 34023 25996
rect 33965 25987 34023 25993
rect 34054 25984 34060 25996
rect 34112 25984 34118 26036
rect 34422 26024 34428 26036
rect 34383 25996 34428 26024
rect 34422 25984 34428 25996
rect 34480 25984 34486 26036
rect 36354 25984 36360 26036
rect 36412 26024 36418 26036
rect 36633 26027 36691 26033
rect 36633 26024 36645 26027
rect 36412 25996 36645 26024
rect 36412 25984 36418 25996
rect 36633 25993 36645 25996
rect 36679 25993 36691 26027
rect 36633 25987 36691 25993
rect 37185 26027 37243 26033
rect 37185 25993 37197 26027
rect 37231 26024 37243 26027
rect 37826 26024 37832 26036
rect 37231 25996 37832 26024
rect 37231 25993 37243 25996
rect 37185 25987 37243 25993
rect 37826 25984 37832 25996
rect 37884 25984 37890 26036
rect 38470 26024 38476 26036
rect 38431 25996 38476 26024
rect 38470 25984 38476 25996
rect 38528 25984 38534 26036
rect 38562 25984 38568 26036
rect 38620 26024 38626 26036
rect 39209 26027 39267 26033
rect 39209 26024 39221 26027
rect 38620 25996 39221 26024
rect 38620 25984 38626 25996
rect 39209 25993 39221 25996
rect 39255 25993 39267 26027
rect 39209 25987 39267 25993
rect 40126 25984 40132 26036
rect 40184 26024 40190 26036
rect 40310 26024 40316 26036
rect 40184 25996 40316 26024
rect 40184 25984 40190 25996
rect 40310 25984 40316 25996
rect 40368 25984 40374 26036
rect 40954 26024 40960 26036
rect 40915 25996 40960 26024
rect 40954 25984 40960 25996
rect 41012 25984 41018 26036
rect 41138 25984 41144 26036
rect 41196 26024 41202 26036
rect 41509 26027 41567 26033
rect 41509 26024 41521 26027
rect 41196 25996 41521 26024
rect 41196 25984 41202 25996
rect 41509 25993 41521 25996
rect 41555 25993 41567 26027
rect 41509 25987 41567 25993
rect 41598 25984 41604 26036
rect 41656 26024 41662 26036
rect 55490 26024 55496 26036
rect 41656 25996 55496 26024
rect 41656 25984 41662 25996
rect 55490 25984 55496 25996
rect 55548 25984 55554 26036
rect 57238 26024 57244 26036
rect 57199 25996 57244 26024
rect 57238 25984 57244 25996
rect 57296 25984 57302 26036
rect 19518 25916 19524 25968
rect 19576 25956 19582 25968
rect 19576 25928 32260 25956
rect 19576 25916 19582 25928
rect 19610 25848 19616 25900
rect 19668 25888 19674 25900
rect 20073 25891 20131 25897
rect 20073 25888 20085 25891
rect 19668 25860 20085 25888
rect 19668 25848 19674 25860
rect 20073 25857 20085 25860
rect 20119 25857 20131 25891
rect 32232 25888 32260 25928
rect 32306 25916 32312 25968
rect 32364 25956 32370 25968
rect 34977 25959 35035 25965
rect 34977 25956 34989 25959
rect 32364 25928 34989 25956
rect 32364 25916 32370 25928
rect 34977 25925 34989 25928
rect 35023 25925 35035 25959
rect 34977 25919 35035 25925
rect 38657 25959 38715 25965
rect 38657 25925 38669 25959
rect 38703 25956 38715 25959
rect 50430 25956 50436 25968
rect 38703 25928 50436 25956
rect 38703 25925 38715 25928
rect 38657 25919 38715 25925
rect 50430 25916 50436 25928
rect 50488 25916 50494 25968
rect 55030 25956 55036 25968
rect 54991 25928 55036 25956
rect 55030 25916 55036 25928
rect 55088 25916 55094 25968
rect 56689 25959 56747 25965
rect 56689 25925 56701 25959
rect 56735 25956 56747 25959
rect 57974 25956 57980 25968
rect 56735 25928 57980 25956
rect 56735 25925 56747 25928
rect 56689 25919 56747 25925
rect 57974 25916 57980 25928
rect 58032 25916 58038 25968
rect 32232 25860 37320 25888
rect 20073 25851 20131 25857
rect 17681 25823 17739 25829
rect 17681 25820 17693 25823
rect 17644 25792 17693 25820
rect 17644 25780 17650 25792
rect 17681 25789 17693 25792
rect 17727 25789 17739 25823
rect 17681 25783 17739 25789
rect 19429 25823 19487 25829
rect 19429 25789 19441 25823
rect 19475 25789 19487 25823
rect 19429 25783 19487 25789
rect 19521 25823 19579 25829
rect 19521 25789 19533 25823
rect 19567 25820 19579 25823
rect 20530 25820 20536 25832
rect 19567 25792 20536 25820
rect 19567 25789 19579 25792
rect 19521 25783 19579 25789
rect 20530 25780 20536 25792
rect 20588 25780 20594 25832
rect 21082 25780 21088 25832
rect 21140 25820 21146 25832
rect 21177 25823 21235 25829
rect 21177 25820 21189 25823
rect 21140 25792 21189 25820
rect 21140 25780 21146 25792
rect 21177 25789 21189 25792
rect 21223 25789 21235 25823
rect 21177 25783 21235 25789
rect 23661 25823 23719 25829
rect 23661 25789 23673 25823
rect 23707 25820 23719 25823
rect 23750 25820 23756 25832
rect 23707 25792 23756 25820
rect 23707 25789 23719 25792
rect 23661 25783 23719 25789
rect 23750 25780 23756 25792
rect 23808 25780 23814 25832
rect 26326 25820 26332 25832
rect 26287 25792 26332 25820
rect 26326 25780 26332 25792
rect 26384 25780 26390 25832
rect 26786 25820 26792 25832
rect 26747 25792 26792 25820
rect 26786 25780 26792 25792
rect 26844 25780 26850 25832
rect 29365 25823 29423 25829
rect 29365 25789 29377 25823
rect 29411 25820 29423 25823
rect 29454 25820 29460 25832
rect 29411 25792 29460 25820
rect 29411 25789 29423 25792
rect 29365 25783 29423 25789
rect 29454 25780 29460 25792
rect 29512 25820 29518 25832
rect 32769 25823 32827 25829
rect 32769 25820 32781 25823
rect 29512 25792 32781 25820
rect 29512 25780 29518 25792
rect 32769 25789 32781 25792
rect 32815 25820 32827 25823
rect 33318 25820 33324 25832
rect 32815 25792 33180 25820
rect 33279 25792 33324 25820
rect 32815 25789 32827 25792
rect 32769 25783 32827 25789
rect 5718 25712 5724 25764
rect 5776 25752 5782 25764
rect 30926 25752 30932 25764
rect 5776 25724 30932 25752
rect 5776 25712 5782 25724
rect 30926 25712 30932 25724
rect 30984 25712 30990 25764
rect 33152 25752 33180 25792
rect 33318 25780 33324 25792
rect 33376 25780 33382 25832
rect 34974 25780 34980 25832
rect 35032 25820 35038 25832
rect 35161 25823 35219 25829
rect 35161 25820 35173 25823
rect 35032 25792 35173 25820
rect 35032 25780 35038 25792
rect 35161 25789 35173 25792
rect 35207 25820 35219 25823
rect 35621 25823 35679 25829
rect 35621 25820 35633 25823
rect 35207 25792 35633 25820
rect 35207 25789 35219 25792
rect 35161 25783 35219 25789
rect 35621 25789 35633 25792
rect 35667 25789 35679 25823
rect 35621 25783 35679 25789
rect 36814 25780 36820 25832
rect 36872 25820 36878 25832
rect 37185 25823 37243 25829
rect 37185 25820 37197 25823
rect 36872 25792 37197 25820
rect 36872 25780 36878 25792
rect 37185 25789 37197 25792
rect 37231 25789 37243 25823
rect 37185 25783 37243 25789
rect 33502 25752 33508 25764
rect 33152 25724 33508 25752
rect 33502 25712 33508 25724
rect 33560 25712 33566 25764
rect 37292 25752 37320 25860
rect 37642 25848 37648 25900
rect 37700 25888 37706 25900
rect 55493 25891 55551 25897
rect 55493 25888 55505 25891
rect 37700 25860 55505 25888
rect 37700 25848 37706 25860
rect 55493 25857 55505 25860
rect 55539 25888 55551 25891
rect 56042 25888 56048 25900
rect 55539 25860 56048 25888
rect 55539 25857 55551 25860
rect 55493 25851 55551 25857
rect 56042 25848 56048 25860
rect 56100 25848 56106 25900
rect 56137 25891 56195 25897
rect 56137 25857 56149 25891
rect 56183 25888 56195 25891
rect 57701 25891 57759 25897
rect 57701 25888 57713 25891
rect 56183 25860 57713 25888
rect 56183 25857 56195 25860
rect 56137 25851 56195 25857
rect 57701 25857 57713 25860
rect 57747 25888 57759 25891
rect 58066 25888 58072 25900
rect 57747 25860 58072 25888
rect 57747 25857 57759 25860
rect 57701 25851 57759 25857
rect 58066 25848 58072 25860
rect 58124 25848 58130 25900
rect 37369 25823 37427 25829
rect 37369 25789 37381 25823
rect 37415 25820 37427 25823
rect 37550 25820 37556 25832
rect 37415 25792 37556 25820
rect 37415 25789 37427 25792
rect 37369 25783 37427 25789
rect 37550 25780 37556 25792
rect 37608 25820 37614 25832
rect 37734 25820 37740 25832
rect 37608 25792 37740 25820
rect 37608 25780 37614 25792
rect 37734 25780 37740 25792
rect 37792 25780 37798 25832
rect 38654 25780 38660 25832
rect 38712 25820 38718 25832
rect 39850 25820 39856 25832
rect 38712 25792 39856 25820
rect 38712 25780 38718 25792
rect 39850 25780 39856 25792
rect 39908 25780 39914 25832
rect 39942 25780 39948 25832
rect 40000 25820 40006 25832
rect 41598 25820 41604 25832
rect 40000 25792 41604 25820
rect 40000 25780 40006 25792
rect 41598 25780 41604 25792
rect 41656 25780 41662 25832
rect 38010 25752 38016 25764
rect 37292 25724 38016 25752
rect 38010 25712 38016 25724
rect 38068 25752 38074 25764
rect 38562 25761 38568 25764
rect 38289 25755 38347 25761
rect 38289 25752 38301 25755
rect 38068 25724 38301 25752
rect 38068 25712 38074 25724
rect 38289 25721 38301 25724
rect 38335 25721 38347 25755
rect 38289 25715 38347 25721
rect 38505 25755 38568 25761
rect 38505 25721 38517 25755
rect 38551 25721 38568 25755
rect 38505 25715 38568 25721
rect 38562 25712 38568 25715
rect 38620 25712 38626 25764
rect 56686 25712 56692 25764
rect 56744 25752 56750 25764
rect 57793 25755 57851 25761
rect 57793 25752 57805 25755
rect 56744 25724 57805 25752
rect 56744 25712 56750 25724
rect 57793 25721 57805 25724
rect 57839 25721 57851 25755
rect 57793 25715 57851 25721
rect 9858 25684 9864 25696
rect 9819 25656 9864 25684
rect 9858 25644 9864 25656
rect 9916 25644 9922 25696
rect 23658 25644 23664 25696
rect 23716 25684 23722 25696
rect 26605 25687 26663 25693
rect 26605 25684 26617 25687
rect 23716 25656 26617 25684
rect 23716 25644 23722 25656
rect 26605 25653 26617 25656
rect 26651 25653 26663 25687
rect 26605 25647 26663 25653
rect 57422 25644 57428 25696
rect 57480 25684 57486 25696
rect 57701 25687 57759 25693
rect 57701 25684 57713 25687
rect 57480 25656 57713 25684
rect 57480 25644 57486 25656
rect 57701 25653 57713 25656
rect 57747 25653 57759 25687
rect 57701 25647 57759 25653
rect 1104 25594 58880 25616
rect 1104 25542 20246 25594
rect 20298 25542 20310 25594
rect 20362 25542 20374 25594
rect 20426 25542 20438 25594
rect 20490 25542 39510 25594
rect 39562 25542 39574 25594
rect 39626 25542 39638 25594
rect 39690 25542 39702 25594
rect 39754 25542 58880 25594
rect 1104 25520 58880 25542
rect 2777 25483 2835 25489
rect 2777 25449 2789 25483
rect 2823 25480 2835 25483
rect 3326 25480 3332 25492
rect 2823 25452 3332 25480
rect 2823 25449 2835 25452
rect 2777 25443 2835 25449
rect 3326 25440 3332 25452
rect 3384 25440 3390 25492
rect 9398 25440 9404 25492
rect 9456 25480 9462 25492
rect 9953 25483 10011 25489
rect 9953 25480 9965 25483
rect 9456 25452 9965 25480
rect 9456 25440 9462 25452
rect 9953 25449 9965 25452
rect 9999 25449 10011 25483
rect 9953 25443 10011 25449
rect 16758 25440 16764 25492
rect 16816 25480 16822 25492
rect 16945 25483 17003 25489
rect 16945 25480 16957 25483
rect 16816 25452 16957 25480
rect 16816 25440 16822 25452
rect 16945 25449 16957 25452
rect 16991 25449 17003 25483
rect 16945 25443 17003 25449
rect 17586 25440 17592 25492
rect 17644 25480 17650 25492
rect 17773 25483 17831 25489
rect 17773 25480 17785 25483
rect 17644 25452 17785 25480
rect 17644 25440 17650 25452
rect 17773 25449 17785 25452
rect 17819 25449 17831 25483
rect 32582 25480 32588 25492
rect 17773 25443 17831 25449
rect 17880 25452 32588 25480
rect 12250 25372 12256 25424
rect 12308 25412 12314 25424
rect 17880 25412 17908 25452
rect 32582 25440 32588 25452
rect 32640 25440 32646 25492
rect 33870 25440 33876 25492
rect 33928 25480 33934 25492
rect 34241 25483 34299 25489
rect 34241 25480 34253 25483
rect 33928 25452 34253 25480
rect 33928 25440 33934 25452
rect 34241 25449 34253 25452
rect 34287 25449 34299 25483
rect 34241 25443 34299 25449
rect 35621 25483 35679 25489
rect 35621 25449 35633 25483
rect 35667 25480 35679 25483
rect 35710 25480 35716 25492
rect 35667 25452 35716 25480
rect 35667 25449 35679 25452
rect 35621 25443 35679 25449
rect 35710 25440 35716 25452
rect 35768 25440 35774 25492
rect 37458 25440 37464 25492
rect 37516 25480 37522 25492
rect 37645 25483 37703 25489
rect 37645 25480 37657 25483
rect 37516 25452 37657 25480
rect 37516 25440 37522 25452
rect 37645 25449 37657 25452
rect 37691 25449 37703 25483
rect 37645 25443 37703 25449
rect 38746 25440 38752 25492
rect 38804 25480 38810 25492
rect 39669 25483 39727 25489
rect 39669 25480 39681 25483
rect 38804 25452 39681 25480
rect 38804 25440 38810 25452
rect 39669 25449 39681 25452
rect 39715 25449 39727 25483
rect 57422 25480 57428 25492
rect 57383 25452 57428 25480
rect 39669 25443 39727 25449
rect 57422 25440 57428 25452
rect 57480 25440 57486 25492
rect 12308 25384 17908 25412
rect 12308 25372 12314 25384
rect 17954 25372 17960 25424
rect 18012 25412 18018 25424
rect 56870 25412 56876 25424
rect 18012 25384 56876 25412
rect 18012 25372 18018 25384
rect 56870 25372 56876 25384
rect 56928 25412 56934 25424
rect 57977 25415 58035 25421
rect 57977 25412 57989 25415
rect 56928 25384 57989 25412
rect 56928 25372 56934 25384
rect 57977 25381 57989 25384
rect 58023 25381 58035 25415
rect 57977 25375 58035 25381
rect 58161 25415 58219 25421
rect 58161 25381 58173 25415
rect 58207 25412 58219 25415
rect 58434 25412 58440 25424
rect 58207 25384 58440 25412
rect 58207 25381 58219 25384
rect 58161 25375 58219 25381
rect 58434 25372 58440 25384
rect 58492 25372 58498 25424
rect 1581 25347 1639 25353
rect 1581 25313 1593 25347
rect 1627 25344 1639 25347
rect 1627 25316 2268 25344
rect 1627 25313 1639 25316
rect 1581 25307 1639 25313
rect 1394 25208 1400 25220
rect 1355 25180 1400 25208
rect 1394 25168 1400 25180
rect 1452 25168 1458 25220
rect 2240 25217 2268 25316
rect 16758 25304 16764 25356
rect 16816 25344 16822 25356
rect 18785 25347 18843 25353
rect 18785 25344 18797 25347
rect 16816 25316 18797 25344
rect 16816 25304 16822 25316
rect 18785 25313 18797 25316
rect 18831 25313 18843 25347
rect 18785 25307 18843 25313
rect 37734 25304 37740 25356
rect 37792 25344 37798 25356
rect 38197 25347 38255 25353
rect 38197 25344 38209 25347
rect 37792 25316 38209 25344
rect 37792 25304 37798 25316
rect 38197 25313 38209 25316
rect 38243 25313 38255 25347
rect 38197 25307 38255 25313
rect 38381 25347 38439 25353
rect 38381 25313 38393 25347
rect 38427 25313 38439 25347
rect 38381 25307 38439 25313
rect 33502 25276 33508 25288
rect 33415 25248 33508 25276
rect 33502 25236 33508 25248
rect 33560 25276 33566 25288
rect 33560 25248 37596 25276
rect 33560 25236 33566 25248
rect 2225 25211 2283 25217
rect 2225 25177 2237 25211
rect 2271 25208 2283 25211
rect 23658 25208 23664 25220
rect 2271 25180 23664 25208
rect 2271 25177 2283 25180
rect 2225 25171 2283 25177
rect 23658 25168 23664 25180
rect 23716 25168 23722 25220
rect 36170 25208 36176 25220
rect 36083 25180 36176 25208
rect 36170 25168 36176 25180
rect 36228 25208 36234 25220
rect 37458 25208 37464 25220
rect 36228 25180 37464 25208
rect 36228 25168 36234 25180
rect 37458 25168 37464 25180
rect 37516 25168 37522 25220
rect 36446 25100 36452 25152
rect 36504 25140 36510 25152
rect 36722 25140 36728 25152
rect 36504 25112 36728 25140
rect 36504 25100 36510 25112
rect 36722 25100 36728 25112
rect 36780 25140 36786 25152
rect 36909 25143 36967 25149
rect 36909 25140 36921 25143
rect 36780 25112 36921 25140
rect 36780 25100 36786 25112
rect 36909 25109 36921 25112
rect 36955 25109 36967 25143
rect 37568 25140 37596 25248
rect 37918 25236 37924 25288
rect 37976 25276 37982 25288
rect 38396 25276 38424 25307
rect 38562 25304 38568 25356
rect 38620 25344 38626 25356
rect 39013 25347 39071 25353
rect 39013 25344 39025 25347
rect 38620 25316 39025 25344
rect 38620 25304 38626 25316
rect 39013 25313 39025 25316
rect 39059 25313 39071 25347
rect 39013 25307 39071 25313
rect 39209 25347 39267 25353
rect 39209 25313 39221 25347
rect 39255 25344 39267 25347
rect 39298 25344 39304 25356
rect 39255 25316 39304 25344
rect 39255 25313 39267 25316
rect 39209 25307 39267 25313
rect 39298 25304 39304 25316
rect 39356 25304 39362 25356
rect 39390 25304 39396 25356
rect 39448 25344 39454 25356
rect 40589 25347 40647 25353
rect 40589 25344 40601 25347
rect 39448 25316 40601 25344
rect 39448 25304 39454 25316
rect 40589 25313 40601 25316
rect 40635 25313 40647 25347
rect 40589 25307 40647 25313
rect 56781 25347 56839 25353
rect 56781 25313 56793 25347
rect 56827 25344 56839 25347
rect 57238 25344 57244 25356
rect 56827 25316 57244 25344
rect 56827 25313 56839 25316
rect 56781 25307 56839 25313
rect 57238 25304 57244 25316
rect 57296 25304 57302 25356
rect 39114 25276 39120 25288
rect 37976 25248 38424 25276
rect 39075 25248 39120 25276
rect 37976 25236 37982 25248
rect 39114 25236 39120 25248
rect 39172 25236 39178 25288
rect 38473 25211 38531 25217
rect 38473 25177 38485 25211
rect 38519 25208 38531 25211
rect 47854 25208 47860 25220
rect 38519 25180 47860 25208
rect 38519 25177 38531 25180
rect 38473 25171 38531 25177
rect 47854 25168 47860 25180
rect 47912 25168 47918 25220
rect 39390 25140 39396 25152
rect 37568 25112 39396 25140
rect 36909 25103 36967 25109
rect 39390 25100 39396 25112
rect 39448 25100 39454 25152
rect 55674 25140 55680 25152
rect 55635 25112 55680 25140
rect 55674 25100 55680 25112
rect 55732 25100 55738 25152
rect 1104 25050 58880 25072
rect 1104 24998 10614 25050
rect 10666 24998 10678 25050
rect 10730 24998 10742 25050
rect 10794 24998 10806 25050
rect 10858 24998 29878 25050
rect 29930 24998 29942 25050
rect 29994 24998 30006 25050
rect 30058 24998 30070 25050
rect 30122 24998 49142 25050
rect 49194 24998 49206 25050
rect 49258 24998 49270 25050
rect 49322 24998 49334 25050
rect 49386 24998 58880 25050
rect 1104 24976 58880 24998
rect 1486 24936 1492 24948
rect 1447 24908 1492 24936
rect 1486 24896 1492 24908
rect 1544 24896 1550 24948
rect 1578 24896 1584 24948
rect 1636 24936 1642 24948
rect 1949 24939 2007 24945
rect 1949 24936 1961 24939
rect 1636 24908 1961 24936
rect 1636 24896 1642 24908
rect 1949 24905 1961 24908
rect 1995 24905 2007 24939
rect 1949 24899 2007 24905
rect 34330 24896 34336 24948
rect 34388 24936 34394 24948
rect 34425 24939 34483 24945
rect 34425 24936 34437 24939
rect 34388 24908 34437 24936
rect 34388 24896 34394 24908
rect 34425 24905 34437 24908
rect 34471 24905 34483 24939
rect 34425 24899 34483 24905
rect 34532 24908 42518 24936
rect 29638 24828 29644 24880
rect 29696 24868 29702 24880
rect 34532 24868 34560 24908
rect 38010 24868 38016 24880
rect 29696 24840 34560 24868
rect 37971 24840 38016 24868
rect 29696 24828 29702 24840
rect 38010 24828 38016 24840
rect 38068 24828 38074 24880
rect 38470 24828 38476 24880
rect 38528 24868 38534 24880
rect 39117 24871 39175 24877
rect 39117 24868 39129 24871
rect 38528 24840 39129 24868
rect 38528 24828 38534 24840
rect 39117 24837 39129 24840
rect 39163 24868 39175 24871
rect 39669 24871 39727 24877
rect 39669 24868 39681 24871
rect 39163 24840 39681 24868
rect 39163 24837 39175 24840
rect 39117 24831 39175 24837
rect 39669 24837 39681 24840
rect 39715 24868 39727 24871
rect 39942 24868 39948 24880
rect 39715 24840 39948 24868
rect 39715 24837 39727 24840
rect 39669 24831 39727 24837
rect 39942 24828 39948 24840
rect 40000 24828 40006 24880
rect 42490 24868 42518 24908
rect 54386 24896 54392 24948
rect 54444 24936 54450 24948
rect 56413 24939 56471 24945
rect 56413 24936 56425 24939
rect 54444 24908 56425 24936
rect 54444 24896 54450 24908
rect 56413 24905 56425 24908
rect 56459 24936 56471 24939
rect 56686 24936 56692 24948
rect 56459 24908 56692 24936
rect 56459 24905 56471 24908
rect 56413 24899 56471 24905
rect 56686 24896 56692 24908
rect 56744 24896 56750 24948
rect 56778 24896 56784 24948
rect 56836 24936 56842 24948
rect 56962 24936 56968 24948
rect 56836 24908 56968 24936
rect 56836 24896 56842 24908
rect 56962 24896 56968 24908
rect 57020 24896 57026 24948
rect 55674 24868 55680 24880
rect 42490 24840 55680 24868
rect 55674 24828 55680 24840
rect 55732 24828 55738 24880
rect 38028 24800 38056 24828
rect 38565 24803 38623 24809
rect 38565 24800 38577 24803
rect 38028 24772 38577 24800
rect 38565 24769 38577 24772
rect 38611 24769 38623 24803
rect 38565 24763 38623 24769
rect 39390 24760 39396 24812
rect 39448 24800 39454 24812
rect 40129 24803 40187 24809
rect 40129 24800 40141 24803
rect 39448 24772 40141 24800
rect 39448 24760 39454 24772
rect 40129 24769 40141 24772
rect 40175 24769 40187 24803
rect 40129 24763 40187 24769
rect 23566 24732 23572 24744
rect 23527 24704 23572 24732
rect 23566 24692 23572 24704
rect 23624 24692 23630 24744
rect 28997 24735 29055 24741
rect 28997 24701 29009 24735
rect 29043 24732 29055 24735
rect 32306 24732 32312 24744
rect 29043 24704 32312 24732
rect 29043 24701 29055 24704
rect 28997 24695 29055 24701
rect 32306 24692 32312 24704
rect 32364 24692 32370 24744
rect 57517 24735 57575 24741
rect 57517 24701 57529 24735
rect 57563 24732 57575 24735
rect 57882 24732 57888 24744
rect 57563 24704 57888 24732
rect 57563 24701 57575 24704
rect 57517 24695 57575 24701
rect 57882 24692 57888 24704
rect 57940 24732 57946 24744
rect 58161 24735 58219 24741
rect 58161 24732 58173 24735
rect 57940 24704 58173 24732
rect 57940 24692 57946 24704
rect 58161 24701 58173 24704
rect 58207 24701 58219 24735
rect 58161 24695 58219 24701
rect 39850 24624 39856 24676
rect 39908 24664 39914 24676
rect 39908 24636 58020 24664
rect 39908 24624 39914 24636
rect 23474 24596 23480 24608
rect 23435 24568 23480 24596
rect 23474 24556 23480 24568
rect 23532 24556 23538 24608
rect 28902 24596 28908 24608
rect 28863 24568 28908 24596
rect 28902 24556 28908 24568
rect 28960 24556 28966 24608
rect 36722 24596 36728 24608
rect 36683 24568 36728 24596
rect 36722 24556 36728 24568
rect 36780 24556 36786 24608
rect 37274 24596 37280 24608
rect 37235 24568 37280 24596
rect 37274 24556 37280 24568
rect 37332 24556 37338 24608
rect 57992 24605 58020 24636
rect 57977 24599 58035 24605
rect 57977 24565 57989 24599
rect 58023 24565 58035 24599
rect 57977 24559 58035 24565
rect 1104 24506 58880 24528
rect 1104 24454 20246 24506
rect 20298 24454 20310 24506
rect 20362 24454 20374 24506
rect 20426 24454 20438 24506
rect 20490 24454 39510 24506
rect 39562 24454 39574 24506
rect 39626 24454 39638 24506
rect 39690 24454 39702 24506
rect 39754 24454 58880 24506
rect 1104 24432 58880 24454
rect 37550 24352 37556 24404
rect 37608 24392 37614 24404
rect 39025 24395 39083 24401
rect 39025 24392 39037 24395
rect 37608 24364 39037 24392
rect 37608 24352 37614 24364
rect 39025 24361 39037 24364
rect 39071 24361 39083 24395
rect 56870 24392 56876 24404
rect 56831 24364 56876 24392
rect 39025 24355 39083 24361
rect 56870 24352 56876 24364
rect 56928 24352 56934 24404
rect 39132 24296 42518 24324
rect 22649 24259 22707 24265
rect 22649 24225 22661 24259
rect 22695 24225 22707 24259
rect 22649 24219 22707 24225
rect 22833 24259 22891 24265
rect 22833 24225 22845 24259
rect 22879 24256 22891 24259
rect 23106 24256 23112 24268
rect 22879 24228 23112 24256
rect 22879 24225 22891 24228
rect 22833 24219 22891 24225
rect 22664 24188 22692 24219
rect 23106 24216 23112 24228
rect 23164 24216 23170 24268
rect 27430 24216 27436 24268
rect 27488 24256 27494 24268
rect 28169 24259 28227 24265
rect 28169 24256 28181 24259
rect 27488 24228 28181 24256
rect 27488 24216 27494 24228
rect 28169 24225 28181 24228
rect 28215 24225 28227 24259
rect 28169 24219 28227 24225
rect 28353 24259 28411 24265
rect 28353 24225 28365 24259
rect 28399 24256 28411 24259
rect 28442 24256 28448 24268
rect 28399 24228 28448 24256
rect 28399 24225 28411 24228
rect 28353 24219 28411 24225
rect 28442 24216 28448 24228
rect 28500 24256 28506 24268
rect 28902 24256 28908 24268
rect 28500 24228 28908 24256
rect 28500 24216 28506 24228
rect 28902 24216 28908 24228
rect 28960 24216 28966 24268
rect 37734 24256 37740 24268
rect 37695 24228 37740 24256
rect 37734 24216 37740 24228
rect 37792 24216 37798 24268
rect 39132 24265 39160 24296
rect 38289 24259 38347 24265
rect 38289 24225 38301 24259
rect 38335 24256 38347 24259
rect 39117 24259 39175 24265
rect 38335 24228 39068 24256
rect 38335 24225 38347 24228
rect 38289 24219 38347 24225
rect 23474 24188 23480 24200
rect 22664 24160 23480 24188
rect 23474 24148 23480 24160
rect 23532 24148 23538 24200
rect 38470 24188 38476 24200
rect 38431 24160 38476 24188
rect 38470 24148 38476 24160
rect 38528 24148 38534 24200
rect 39040 24188 39068 24228
rect 39117 24225 39129 24259
rect 39163 24256 39175 24259
rect 39206 24256 39212 24268
rect 39163 24228 39212 24256
rect 39163 24225 39175 24228
rect 39117 24219 39175 24225
rect 39206 24216 39212 24228
rect 39264 24216 39270 24268
rect 39761 24259 39819 24265
rect 39761 24225 39773 24259
rect 39807 24256 39819 24259
rect 39807 24228 40724 24256
rect 39807 24225 39819 24228
rect 39761 24219 39819 24225
rect 39298 24188 39304 24200
rect 39040 24160 39304 24188
rect 39298 24148 39304 24160
rect 39356 24188 39362 24200
rect 39669 24191 39727 24197
rect 39669 24188 39681 24191
rect 39356 24160 39681 24188
rect 39356 24148 39362 24160
rect 39669 24157 39681 24160
rect 39715 24157 39727 24191
rect 39669 24151 39727 24157
rect 3510 24080 3516 24132
rect 3568 24120 3574 24132
rect 22557 24123 22615 24129
rect 22557 24120 22569 24123
rect 3568 24092 22569 24120
rect 3568 24080 3574 24092
rect 22557 24089 22569 24092
rect 22603 24089 22615 24123
rect 28350 24120 28356 24132
rect 28311 24092 28356 24120
rect 22557 24083 22615 24089
rect 28350 24080 28356 24092
rect 28408 24080 28414 24132
rect 40696 24064 40724 24228
rect 42490 24188 42518 24296
rect 57517 24259 57575 24265
rect 57517 24225 57529 24259
rect 57563 24256 57575 24259
rect 57882 24256 57888 24268
rect 57563 24228 57888 24256
rect 57563 24225 57575 24228
rect 57517 24219 57575 24225
rect 57882 24216 57888 24228
rect 57940 24256 57946 24268
rect 58161 24259 58219 24265
rect 58161 24256 58173 24259
rect 57940 24228 58173 24256
rect 57940 24216 57946 24228
rect 58161 24225 58173 24228
rect 58207 24225 58219 24259
rect 58161 24219 58219 24225
rect 57790 24188 57796 24200
rect 42490 24160 57796 24188
rect 57790 24148 57796 24160
rect 57848 24148 57854 24200
rect 40678 24052 40684 24064
rect 40639 24024 40684 24052
rect 40678 24012 40684 24024
rect 40736 24012 40742 24064
rect 57974 24052 57980 24064
rect 57935 24024 57980 24052
rect 57974 24012 57980 24024
rect 58032 24012 58038 24064
rect 1104 23962 58880 23984
rect 1104 23910 10614 23962
rect 10666 23910 10678 23962
rect 10730 23910 10742 23962
rect 10794 23910 10806 23962
rect 10858 23910 29878 23962
rect 29930 23910 29942 23962
rect 29994 23910 30006 23962
rect 30058 23910 30070 23962
rect 30122 23910 49142 23962
rect 49194 23910 49206 23962
rect 49258 23910 49270 23962
rect 49322 23910 49334 23962
rect 49386 23910 58880 23962
rect 1104 23888 58880 23910
rect 1486 23848 1492 23860
rect 1447 23820 1492 23848
rect 1486 23808 1492 23820
rect 1544 23808 1550 23860
rect 22557 23851 22615 23857
rect 22557 23817 22569 23851
rect 22603 23848 22615 23851
rect 22738 23848 22744 23860
rect 22603 23820 22744 23848
rect 22603 23817 22615 23820
rect 22557 23811 22615 23817
rect 22738 23808 22744 23820
rect 22796 23808 22802 23860
rect 39206 23848 39212 23860
rect 39167 23820 39212 23848
rect 39206 23808 39212 23820
rect 39264 23808 39270 23860
rect 40678 23808 40684 23860
rect 40736 23848 40742 23860
rect 57974 23848 57980 23860
rect 40736 23820 57980 23848
rect 40736 23808 40742 23820
rect 57974 23808 57980 23820
rect 58032 23808 58038 23860
rect 37001 23783 37059 23789
rect 37001 23749 37013 23783
rect 37047 23780 37059 23783
rect 37734 23780 37740 23792
rect 37047 23752 37740 23780
rect 37047 23749 37059 23752
rect 37001 23743 37059 23749
rect 37734 23740 37740 23752
rect 37792 23740 37798 23792
rect 23474 23672 23480 23724
rect 23532 23712 23538 23724
rect 28442 23712 28448 23724
rect 23532 23684 26004 23712
rect 23532 23672 23538 23684
rect 22554 23644 22560 23656
rect 22515 23616 22560 23644
rect 22554 23604 22560 23616
rect 22612 23604 22618 23656
rect 22738 23644 22744 23656
rect 22699 23616 22744 23644
rect 22738 23604 22744 23616
rect 22796 23644 22802 23656
rect 25976 23653 26004 23684
rect 28092 23684 28448 23712
rect 28092 23653 28120 23684
rect 28442 23672 28448 23684
rect 28500 23672 28506 23724
rect 25777 23647 25835 23653
rect 25777 23644 25789 23647
rect 22796 23616 25789 23644
rect 22796 23604 22802 23616
rect 25777 23613 25789 23616
rect 25823 23613 25835 23647
rect 25777 23607 25835 23613
rect 25961 23647 26019 23653
rect 25961 23613 25973 23647
rect 26007 23613 26019 23647
rect 25961 23607 26019 23613
rect 28077 23647 28135 23653
rect 28077 23613 28089 23647
rect 28123 23613 28135 23647
rect 28534 23644 28540 23656
rect 28495 23616 28540 23644
rect 28077 23607 28135 23613
rect 1581 23579 1639 23585
rect 1581 23545 1593 23579
rect 1627 23576 1639 23579
rect 1627 23548 2176 23576
rect 1627 23545 1639 23548
rect 1581 23539 1639 23545
rect 2148 23520 2176 23548
rect 2130 23508 2136 23520
rect 2091 23480 2136 23508
rect 2130 23468 2136 23480
rect 2188 23468 2194 23520
rect 25792 23508 25820 23607
rect 28534 23604 28540 23616
rect 28592 23604 28598 23656
rect 57517 23647 57575 23653
rect 57517 23613 57529 23647
rect 57563 23644 57575 23647
rect 58158 23644 58164 23656
rect 57563 23616 58164 23644
rect 57563 23613 57575 23616
rect 57517 23607 57575 23613
rect 58158 23604 58164 23616
rect 58216 23604 58222 23656
rect 26145 23579 26203 23585
rect 26145 23545 26157 23579
rect 26191 23576 26203 23579
rect 26234 23576 26240 23588
rect 26191 23548 26240 23576
rect 26191 23545 26203 23548
rect 26145 23539 26203 23545
rect 26234 23536 26240 23548
rect 26292 23536 26298 23588
rect 35894 23536 35900 23588
rect 35952 23576 35958 23588
rect 36817 23579 36875 23585
rect 36817 23576 36829 23579
rect 35952 23548 36829 23576
rect 35952 23536 35958 23548
rect 36817 23545 36829 23548
rect 36863 23545 36875 23579
rect 36817 23539 36875 23545
rect 27430 23508 27436 23520
rect 25792 23480 27436 23508
rect 27430 23468 27436 23480
rect 27488 23468 27494 23520
rect 28258 23508 28264 23520
rect 28219 23480 28264 23508
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 36722 23468 36728 23520
rect 36780 23508 36786 23520
rect 39942 23508 39948 23520
rect 36780 23480 39948 23508
rect 36780 23468 36786 23480
rect 39942 23468 39948 23480
rect 40000 23468 40006 23520
rect 57790 23468 57796 23520
rect 57848 23508 57854 23520
rect 57977 23511 58035 23517
rect 57977 23508 57989 23511
rect 57848 23480 57989 23508
rect 57848 23468 57854 23480
rect 57977 23477 57989 23480
rect 58023 23477 58035 23511
rect 57977 23471 58035 23477
rect 1104 23418 58880 23440
rect 1104 23366 20246 23418
rect 20298 23366 20310 23418
rect 20362 23366 20374 23418
rect 20426 23366 20438 23418
rect 20490 23366 39510 23418
rect 39562 23366 39574 23418
rect 39626 23366 39638 23418
rect 39690 23366 39702 23418
rect 39754 23366 58880 23418
rect 1104 23344 58880 23366
rect 23106 23264 23112 23316
rect 23164 23304 23170 23316
rect 28534 23304 28540 23316
rect 23164 23276 28540 23304
rect 23164 23264 23170 23276
rect 28534 23264 28540 23276
rect 28592 23264 28598 23316
rect 27430 23236 27436 23248
rect 27391 23208 27436 23236
rect 27430 23196 27436 23208
rect 27488 23196 27494 23248
rect 27614 23236 27620 23248
rect 27575 23208 27620 23236
rect 27614 23196 27620 23208
rect 27672 23196 27678 23248
rect 1394 23168 1400 23180
rect 1355 23140 1400 23168
rect 1394 23128 1400 23140
rect 1452 23128 1458 23180
rect 1581 23171 1639 23177
rect 1581 23137 1593 23171
rect 1627 23168 1639 23171
rect 1627 23140 2268 23168
rect 1627 23137 1639 23140
rect 1581 23131 1639 23137
rect 2240 23041 2268 23140
rect 4154 23128 4160 23180
rect 4212 23168 4218 23180
rect 5077 23171 5135 23177
rect 5077 23168 5089 23171
rect 4212 23140 5089 23168
rect 4212 23128 4218 23140
rect 5077 23137 5089 23140
rect 5123 23137 5135 23171
rect 5077 23131 5135 23137
rect 19981 23171 20039 23177
rect 19981 23137 19993 23171
rect 20027 23168 20039 23171
rect 20625 23171 20683 23177
rect 20625 23168 20637 23171
rect 20027 23140 20637 23168
rect 20027 23137 20039 23140
rect 19981 23131 20039 23137
rect 20625 23137 20637 23140
rect 20671 23137 20683 23171
rect 20625 23131 20683 23137
rect 20717 23171 20775 23177
rect 20717 23137 20729 23171
rect 20763 23168 20775 23171
rect 21174 23168 21180 23180
rect 20763 23140 21180 23168
rect 20763 23137 20775 23140
rect 20717 23131 20775 23137
rect 21174 23128 21180 23140
rect 21232 23168 21238 23180
rect 21545 23171 21603 23177
rect 21545 23168 21557 23171
rect 21232 23140 21557 23168
rect 21232 23128 21238 23140
rect 21545 23137 21557 23140
rect 21591 23137 21603 23171
rect 21545 23131 21603 23137
rect 21821 23171 21879 23177
rect 21821 23137 21833 23171
rect 21867 23168 21879 23171
rect 23106 23168 23112 23180
rect 21867 23140 23112 23168
rect 21867 23137 21879 23140
rect 21821 23131 21879 23137
rect 23106 23128 23112 23140
rect 23164 23128 23170 23180
rect 4890 23100 4896 23112
rect 4851 23072 4896 23100
rect 4890 23060 4896 23072
rect 4948 23060 4954 23112
rect 6426 23072 29638 23100
rect 2225 23035 2283 23041
rect 2225 23001 2237 23035
rect 2271 23032 2283 23035
rect 6426 23032 6454 23072
rect 21542 23032 21548 23044
rect 2271 23004 6454 23032
rect 21503 23004 21548 23032
rect 2271 23001 2283 23004
rect 2225 22995 2283 23001
rect 21542 22992 21548 23004
rect 21600 22992 21606 23044
rect 29610 23032 29638 23072
rect 52454 23032 52460 23044
rect 29610 23004 52460 23032
rect 52454 22992 52460 23004
rect 52512 22992 52518 23044
rect 1670 22924 1676 22976
rect 1728 22964 1734 22976
rect 19981 22967 20039 22973
rect 19981 22964 19993 22967
rect 1728 22936 19993 22964
rect 1728 22924 1734 22936
rect 19981 22933 19993 22936
rect 20027 22964 20039 22967
rect 20073 22967 20131 22973
rect 20073 22964 20085 22967
rect 20027 22936 20085 22964
rect 20027 22933 20039 22936
rect 19981 22927 20039 22933
rect 20073 22933 20085 22936
rect 20119 22933 20131 22967
rect 20073 22927 20131 22933
rect 1104 22874 58880 22896
rect 1104 22822 10614 22874
rect 10666 22822 10678 22874
rect 10730 22822 10742 22874
rect 10794 22822 10806 22874
rect 10858 22822 29878 22874
rect 29930 22822 29942 22874
rect 29994 22822 30006 22874
rect 30058 22822 30070 22874
rect 30122 22822 49142 22874
rect 49194 22822 49206 22874
rect 49258 22822 49270 22874
rect 49322 22822 49334 22874
rect 49386 22822 58880 22874
rect 1104 22800 58880 22822
rect 4154 22760 4160 22772
rect 4115 22732 4160 22760
rect 4154 22720 4160 22732
rect 4212 22720 4218 22772
rect 34606 22720 34612 22772
rect 34664 22760 34670 22772
rect 34885 22763 34943 22769
rect 34885 22760 34897 22763
rect 34664 22732 34897 22760
rect 34664 22720 34670 22732
rect 34885 22729 34897 22732
rect 34931 22729 34943 22763
rect 34885 22723 34943 22729
rect 36449 22763 36507 22769
rect 36449 22729 36461 22763
rect 36495 22760 36507 22763
rect 40218 22760 40224 22772
rect 36495 22732 40224 22760
rect 36495 22729 36507 22732
rect 36449 22723 36507 22729
rect 21174 22556 21180 22568
rect 21135 22528 21180 22556
rect 21174 22516 21180 22528
rect 21232 22516 21238 22568
rect 21453 22559 21511 22565
rect 21453 22525 21465 22559
rect 21499 22556 21511 22559
rect 22738 22556 22744 22568
rect 21499 22528 22744 22556
rect 21499 22525 21511 22528
rect 21453 22519 21511 22525
rect 22738 22516 22744 22528
rect 22796 22516 22802 22568
rect 25958 22516 25964 22568
rect 26016 22556 26022 22568
rect 26421 22559 26479 22565
rect 26421 22556 26433 22559
rect 26016 22528 26433 22556
rect 26016 22516 26022 22528
rect 26421 22525 26433 22528
rect 26467 22525 26479 22559
rect 34900 22556 34928 22723
rect 40218 22720 40224 22732
rect 40276 22720 40282 22772
rect 35437 22559 35495 22565
rect 35437 22556 35449 22559
rect 34900 22528 35449 22556
rect 26421 22519 26479 22525
rect 35437 22525 35449 22528
rect 35483 22525 35495 22559
rect 35437 22519 35495 22525
rect 35529 22559 35587 22565
rect 35529 22525 35541 22559
rect 35575 22556 35587 22559
rect 35986 22556 35992 22568
rect 35575 22528 35992 22556
rect 35575 22525 35587 22528
rect 35529 22519 35587 22525
rect 35986 22516 35992 22528
rect 36044 22556 36050 22568
rect 36449 22559 36507 22565
rect 36449 22556 36461 22559
rect 36044 22528 36461 22556
rect 36044 22516 36050 22528
rect 36449 22525 36461 22528
rect 36495 22525 36507 22559
rect 36449 22519 36507 22525
rect 36538 22516 36544 22568
rect 36596 22556 36602 22568
rect 36633 22559 36691 22565
rect 36633 22556 36645 22559
rect 36596 22528 36645 22556
rect 36596 22516 36602 22528
rect 36633 22525 36645 22528
rect 36679 22525 36691 22559
rect 36633 22519 36691 22525
rect 57517 22559 57575 22565
rect 57517 22525 57529 22559
rect 57563 22556 57575 22559
rect 58158 22556 58164 22568
rect 57563 22528 58164 22556
rect 57563 22525 57575 22528
rect 57517 22519 57575 22525
rect 58158 22516 58164 22528
rect 58216 22516 58222 22568
rect 1394 22488 1400 22500
rect 1355 22460 1400 22488
rect 1394 22448 1400 22460
rect 1452 22448 1458 22500
rect 1581 22491 1639 22497
rect 1581 22457 1593 22491
rect 1627 22488 1639 22491
rect 2225 22491 2283 22497
rect 2225 22488 2237 22491
rect 1627 22460 2237 22488
rect 1627 22457 1639 22460
rect 1581 22451 1639 22457
rect 2225 22457 2237 22460
rect 2271 22488 2283 22491
rect 21085 22491 21143 22497
rect 21085 22488 21097 22491
rect 2271 22460 21097 22488
rect 2271 22457 2283 22460
rect 2225 22451 2283 22457
rect 21085 22457 21097 22460
rect 21131 22457 21143 22491
rect 21085 22451 21143 22457
rect 26513 22423 26571 22429
rect 26513 22389 26525 22423
rect 26559 22420 26571 22423
rect 27430 22420 27436 22432
rect 26559 22392 27436 22420
rect 26559 22389 26571 22392
rect 26513 22383 26571 22389
rect 27430 22380 27436 22392
rect 27488 22380 27494 22432
rect 57977 22423 58035 22429
rect 57977 22389 57989 22423
rect 58023 22420 58035 22423
rect 58250 22420 58256 22432
rect 58023 22392 58256 22420
rect 58023 22389 58035 22392
rect 57977 22383 58035 22389
rect 58250 22380 58256 22392
rect 58308 22380 58314 22432
rect 1104 22330 58880 22352
rect 1104 22278 20246 22330
rect 20298 22278 20310 22330
rect 20362 22278 20374 22330
rect 20426 22278 20438 22330
rect 20490 22278 39510 22330
rect 39562 22278 39574 22330
rect 39626 22278 39638 22330
rect 39690 22278 39702 22330
rect 39754 22278 58880 22330
rect 1104 22256 58880 22278
rect 27341 22219 27399 22225
rect 27341 22185 27353 22219
rect 27387 22216 27399 22219
rect 27798 22216 27804 22228
rect 27387 22188 27804 22216
rect 27387 22185 27399 22188
rect 27341 22179 27399 22185
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 27246 22080 27252 22092
rect 27207 22052 27252 22080
rect 27246 22040 27252 22052
rect 27304 22040 27310 22092
rect 27430 22080 27436 22092
rect 27391 22052 27436 22080
rect 27430 22040 27436 22052
rect 27488 22040 27494 22092
rect 36262 22080 36268 22092
rect 36223 22052 36268 22080
rect 36262 22040 36268 22052
rect 36320 22080 36326 22092
rect 36909 22083 36967 22089
rect 36909 22080 36921 22083
rect 36320 22052 36921 22080
rect 36320 22040 36326 22052
rect 36909 22049 36921 22052
rect 36955 22049 36967 22083
rect 57977 22083 58035 22089
rect 57977 22080 57989 22083
rect 36909 22043 36967 22049
rect 57348 22052 57989 22080
rect 57348 21956 57376 22052
rect 57977 22049 57989 22052
rect 58023 22049 58035 22083
rect 57977 22043 58035 22049
rect 36449 21947 36507 21953
rect 36449 21913 36461 21947
rect 36495 21944 36507 21947
rect 36538 21944 36544 21956
rect 36495 21916 36544 21944
rect 36495 21913 36507 21916
rect 36449 21907 36507 21913
rect 36538 21904 36544 21916
rect 36596 21904 36602 21956
rect 37093 21947 37151 21953
rect 37093 21913 37105 21947
rect 37139 21944 37151 21947
rect 38102 21944 38108 21956
rect 37139 21916 38108 21944
rect 37139 21913 37151 21916
rect 37093 21907 37151 21913
rect 38102 21904 38108 21916
rect 38160 21944 38166 21956
rect 38562 21944 38568 21956
rect 38160 21916 38568 21944
rect 38160 21904 38166 21916
rect 38562 21904 38568 21916
rect 38620 21904 38626 21956
rect 57330 21944 57336 21956
rect 57291 21916 57336 21944
rect 57330 21904 57336 21916
rect 57388 21904 57394 21956
rect 57882 21904 57888 21956
rect 57940 21944 57946 21956
rect 58161 21947 58219 21953
rect 58161 21944 58173 21947
rect 57940 21916 58173 21944
rect 57940 21904 57946 21916
rect 58161 21913 58173 21916
rect 58207 21913 58219 21947
rect 58161 21907 58219 21913
rect 1104 21786 58880 21808
rect 1104 21734 10614 21786
rect 10666 21734 10678 21786
rect 10730 21734 10742 21786
rect 10794 21734 10806 21786
rect 10858 21734 29878 21786
rect 29930 21734 29942 21786
rect 29994 21734 30006 21786
rect 30058 21734 30070 21786
rect 30122 21734 49142 21786
rect 49194 21734 49206 21786
rect 49258 21734 49270 21786
rect 49322 21734 49334 21786
rect 49386 21734 58880 21786
rect 1104 21712 58880 21734
rect 19794 21672 19800 21684
rect 19755 21644 19800 21672
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 19978 21632 19984 21684
rect 20036 21672 20042 21684
rect 20441 21675 20499 21681
rect 20441 21672 20453 21675
rect 20036 21644 20453 21672
rect 20036 21632 20042 21644
rect 20441 21641 20453 21644
rect 20487 21641 20499 21675
rect 29454 21672 29460 21684
rect 29415 21644 29460 21672
rect 20441 21635 20499 21641
rect 29454 21632 29460 21644
rect 29512 21632 29518 21684
rect 31018 21632 31024 21684
rect 31076 21672 31082 21684
rect 31389 21675 31447 21681
rect 31389 21672 31401 21675
rect 31076 21644 31401 21672
rect 31076 21632 31082 21644
rect 31389 21641 31401 21644
rect 31435 21641 31447 21675
rect 31389 21635 31447 21641
rect 23750 21564 23756 21616
rect 23808 21604 23814 21616
rect 36725 21607 36783 21613
rect 36725 21604 36737 21607
rect 23808 21576 36737 21604
rect 23808 21564 23814 21576
rect 36725 21573 36737 21576
rect 36771 21573 36783 21607
rect 36725 21567 36783 21573
rect 20070 21536 20076 21548
rect 19812 21508 20076 21536
rect 19812 21477 19840 21508
rect 20070 21496 20076 21508
rect 20128 21536 20134 21548
rect 38378 21536 38384 21548
rect 20128 21508 20484 21536
rect 20128 21496 20134 21508
rect 20456 21477 20484 21508
rect 27264 21508 30788 21536
rect 27264 21480 27292 21508
rect 19797 21471 19855 21477
rect 19797 21437 19809 21471
rect 19843 21437 19855 21471
rect 19797 21431 19855 21437
rect 19981 21471 20039 21477
rect 19981 21437 19993 21471
rect 20027 21437 20039 21471
rect 19981 21431 20039 21437
rect 20441 21471 20499 21477
rect 20441 21437 20453 21471
rect 20487 21437 20499 21471
rect 20441 21431 20499 21437
rect 20625 21471 20683 21477
rect 20625 21437 20637 21471
rect 20671 21468 20683 21471
rect 27246 21468 27252 21480
rect 20671 21440 27252 21468
rect 20671 21437 20683 21440
rect 20625 21431 20683 21437
rect 19996 21400 20024 21431
rect 27246 21428 27252 21440
rect 27304 21428 27310 21480
rect 27614 21428 27620 21480
rect 27672 21468 27678 21480
rect 28721 21471 28779 21477
rect 27672 21440 28304 21468
rect 27672 21428 27678 21440
rect 28166 21400 28172 21412
rect 19996 21372 28172 21400
rect 28166 21360 28172 21372
rect 28224 21360 28230 21412
rect 28276 21400 28304 21440
rect 28721 21437 28733 21471
rect 28767 21468 28779 21471
rect 29454 21468 29460 21480
rect 28767 21440 29460 21468
rect 28767 21437 28779 21440
rect 28721 21431 28779 21437
rect 29454 21428 29460 21440
rect 29512 21428 29518 21480
rect 30760 21409 30788 21508
rect 36832 21508 38384 21536
rect 31205 21471 31263 21477
rect 31205 21437 31217 21471
rect 31251 21437 31263 21471
rect 31386 21468 31392 21480
rect 31347 21440 31392 21468
rect 31205 21431 31263 21437
rect 30561 21403 30619 21409
rect 30561 21400 30573 21403
rect 28276 21372 30573 21400
rect 30561 21369 30573 21372
rect 30607 21369 30619 21403
rect 30561 21363 30619 21369
rect 30745 21403 30803 21409
rect 30745 21369 30757 21403
rect 30791 21400 30803 21403
rect 31220 21400 31248 21431
rect 31386 21428 31392 21440
rect 31444 21428 31450 21480
rect 35894 21468 35900 21480
rect 35855 21440 35900 21468
rect 35894 21428 35900 21440
rect 35952 21428 35958 21480
rect 36832 21477 36860 21508
rect 38378 21496 38384 21508
rect 38436 21536 38442 21548
rect 38436 21508 38792 21536
rect 38436 21496 38442 21508
rect 36817 21471 36875 21477
rect 36817 21437 36829 21471
rect 36863 21437 36875 21471
rect 36817 21431 36875 21437
rect 36909 21471 36967 21477
rect 36909 21437 36921 21471
rect 36955 21437 36967 21471
rect 36909 21431 36967 21437
rect 31294 21400 31300 21412
rect 30791 21372 31300 21400
rect 30791 21369 30803 21372
rect 30745 21363 30803 21369
rect 28905 21335 28963 21341
rect 28905 21301 28917 21335
rect 28951 21332 28963 21335
rect 29270 21332 29276 21344
rect 28951 21304 29276 21332
rect 28951 21301 28963 21304
rect 28905 21295 28963 21301
rect 29270 21292 29276 21304
rect 29328 21292 29334 21344
rect 30576 21332 30604 21363
rect 31294 21360 31300 21372
rect 31352 21360 31358 21412
rect 35912 21332 35940 21428
rect 36538 21360 36544 21412
rect 36596 21400 36602 21412
rect 36924 21400 36952 21431
rect 37826 21428 37832 21480
rect 37884 21468 37890 21480
rect 38764 21477 38792 21508
rect 38289 21471 38347 21477
rect 38289 21468 38301 21471
rect 37884 21440 38301 21468
rect 37884 21428 37890 21440
rect 38289 21437 38301 21440
rect 38335 21437 38347 21471
rect 38289 21431 38347 21437
rect 38749 21471 38807 21477
rect 38749 21437 38761 21471
rect 38795 21437 38807 21471
rect 38749 21431 38807 21437
rect 36596 21372 36952 21400
rect 39025 21403 39083 21409
rect 36596 21360 36602 21372
rect 39025 21369 39037 21403
rect 39071 21369 39083 21403
rect 39025 21363 39083 21369
rect 36078 21332 36084 21344
rect 30576 21304 35940 21332
rect 36039 21304 36084 21332
rect 36078 21292 36084 21304
rect 36136 21292 36142 21344
rect 39040 21332 39068 21363
rect 56778 21332 56784 21344
rect 39040 21304 56784 21332
rect 56778 21292 56784 21304
rect 56836 21292 56842 21344
rect 1104 21242 58880 21264
rect 1104 21190 20246 21242
rect 20298 21190 20310 21242
rect 20362 21190 20374 21242
rect 20426 21190 20438 21242
rect 20490 21190 39510 21242
rect 39562 21190 39574 21242
rect 39626 21190 39638 21242
rect 39690 21190 39702 21242
rect 39754 21190 58880 21242
rect 1104 21168 58880 21190
rect 1486 21128 1492 21140
rect 1447 21100 1492 21128
rect 1486 21088 1492 21100
rect 1544 21088 1550 21140
rect 20070 21128 20076 21140
rect 20031 21100 20076 21128
rect 20070 21088 20076 21100
rect 20128 21088 20134 21140
rect 28166 21088 28172 21140
rect 28224 21128 28230 21140
rect 54570 21128 54576 21140
rect 28224 21100 29638 21128
rect 28224 21088 28230 21100
rect 28534 21020 28540 21072
rect 28592 21060 28598 21072
rect 28905 21063 28963 21069
rect 28905 21060 28917 21063
rect 28592 21032 28917 21060
rect 28592 21020 28598 21032
rect 28905 21029 28917 21032
rect 28951 21029 28963 21063
rect 29270 21060 29276 21072
rect 29231 21032 29276 21060
rect 28905 21023 28963 21029
rect 29270 21020 29276 21032
rect 29328 21020 29334 21072
rect 29610 21060 29638 21100
rect 32416 21100 54576 21128
rect 32416 21069 32444 21100
rect 54570 21088 54576 21100
rect 54628 21088 54634 21140
rect 32401 21063 32459 21069
rect 29610 21032 31064 21060
rect 1578 20992 1584 21004
rect 1539 20964 1584 20992
rect 1578 20952 1584 20964
rect 1636 20952 1642 21004
rect 20070 20952 20076 21004
rect 20128 20992 20134 21004
rect 20165 20995 20223 21001
rect 20165 20992 20177 20995
rect 20128 20964 20177 20992
rect 20128 20952 20134 20964
rect 20165 20961 20177 20964
rect 20211 20992 20223 20995
rect 20625 20995 20683 21001
rect 20625 20992 20637 20995
rect 20211 20964 20637 20992
rect 20211 20961 20223 20964
rect 20165 20955 20223 20961
rect 20625 20961 20637 20964
rect 20671 20961 20683 20995
rect 20625 20955 20683 20961
rect 27430 20952 27436 21004
rect 27488 20992 27494 21004
rect 27893 20995 27951 21001
rect 27893 20992 27905 20995
rect 27488 20964 27905 20992
rect 27488 20952 27494 20964
rect 27893 20961 27905 20964
rect 27939 20961 27951 20995
rect 28166 20992 28172 21004
rect 28127 20964 28172 20992
rect 27893 20955 27951 20961
rect 28166 20952 28172 20964
rect 28224 20952 28230 21004
rect 29288 20992 29316 21020
rect 30929 20995 30987 21001
rect 30929 20992 30941 20995
rect 29288 20964 30941 20992
rect 27706 20924 27712 20936
rect 27667 20896 27712 20924
rect 27706 20884 27712 20896
rect 27764 20884 27770 20936
rect 30576 20856 30604 20964
rect 30929 20961 30941 20964
rect 30975 20961 30987 20995
rect 30929 20955 30987 20961
rect 30653 20927 30711 20933
rect 30653 20893 30665 20927
rect 30699 20924 30711 20927
rect 31036 20924 31064 21032
rect 32401 21029 32413 21063
rect 32447 21029 32459 21063
rect 32401 21023 32459 21029
rect 36078 21020 36084 21072
rect 36136 21060 36142 21072
rect 50801 21063 50859 21069
rect 36136 21032 37412 21060
rect 36136 21020 36142 21032
rect 31665 20995 31723 21001
rect 31665 20961 31677 20995
rect 31711 20961 31723 20995
rect 32214 20992 32220 21004
rect 32175 20964 32220 20992
rect 31665 20955 31723 20961
rect 31110 20924 31116 20936
rect 30699 20896 31116 20924
rect 30699 20893 30711 20896
rect 30653 20887 30711 20893
rect 31110 20884 31116 20896
rect 31168 20924 31174 20936
rect 31680 20924 31708 20955
rect 32214 20952 32220 20964
rect 32272 20952 32278 21004
rect 35986 20992 35992 21004
rect 35947 20964 35992 20992
rect 35986 20952 35992 20964
rect 36044 20952 36050 21004
rect 36556 21001 36584 21032
rect 37384 21001 37412 21032
rect 50801 21029 50813 21063
rect 50847 21060 50859 21063
rect 50847 21032 51534 21060
rect 50847 21029 50859 21032
rect 50801 21023 50859 21029
rect 36541 20995 36599 21001
rect 36541 20961 36553 20995
rect 36587 20961 36599 20995
rect 36541 20955 36599 20961
rect 37185 20995 37243 21001
rect 37185 20961 37197 20995
rect 37231 20961 37243 20995
rect 37185 20955 37243 20961
rect 37369 20995 37427 21001
rect 37369 20961 37381 20995
rect 37415 20992 37427 20995
rect 37826 20992 37832 21004
rect 37415 20964 37832 20992
rect 37415 20961 37427 20964
rect 37369 20955 37427 20961
rect 36078 20924 36084 20936
rect 31168 20896 31708 20924
rect 36039 20896 36084 20924
rect 31168 20884 31174 20896
rect 36078 20884 36084 20896
rect 36136 20884 36142 20936
rect 36630 20884 36636 20936
rect 36688 20924 36694 20936
rect 37001 20927 37059 20933
rect 37001 20924 37013 20927
rect 36688 20896 37013 20924
rect 36688 20884 36694 20896
rect 37001 20893 37013 20896
rect 37047 20893 37059 20927
rect 37001 20887 37059 20893
rect 37090 20884 37096 20936
rect 37148 20924 37154 20936
rect 37200 20924 37228 20955
rect 37826 20952 37832 20964
rect 37884 20952 37890 21004
rect 38010 20992 38016 21004
rect 37971 20964 38016 20992
rect 38010 20952 38016 20964
rect 38068 20952 38074 21004
rect 38838 20992 38844 21004
rect 38799 20964 38844 20992
rect 38838 20952 38844 20964
rect 38896 20952 38902 21004
rect 47210 20952 47216 21004
rect 47268 20992 47274 21004
rect 48133 20995 48191 21001
rect 48133 20992 48145 20995
rect 47268 20964 48145 20992
rect 47268 20952 47274 20964
rect 48133 20961 48145 20964
rect 48179 20961 48191 20995
rect 48133 20955 48191 20961
rect 48225 20995 48283 21001
rect 48225 20961 48237 20995
rect 48271 20992 48283 20995
rect 51506 20992 51534 21032
rect 54386 20992 54392 21004
rect 48271 20964 51120 20992
rect 51506 20964 54392 20992
rect 48271 20961 48283 20964
rect 48225 20955 48283 20961
rect 38749 20927 38807 20933
rect 38749 20924 38761 20927
rect 37148 20896 38761 20924
rect 37148 20884 37154 20896
rect 38749 20893 38761 20896
rect 38795 20893 38807 20927
rect 38749 20887 38807 20893
rect 47394 20884 47400 20936
rect 47452 20924 47458 20936
rect 48317 20927 48375 20933
rect 48317 20924 48329 20927
rect 47452 20896 48329 20924
rect 47452 20884 47458 20896
rect 48317 20893 48329 20896
rect 48363 20924 48375 20927
rect 50801 20927 50859 20933
rect 50801 20924 50813 20927
rect 48363 20896 50813 20924
rect 48363 20893 48375 20896
rect 48317 20887 48375 20893
rect 50801 20893 50813 20896
rect 50847 20893 50859 20927
rect 51092 20924 51120 20964
rect 54386 20952 54392 20964
rect 54444 20952 54450 21004
rect 57517 20995 57575 21001
rect 57517 20961 57529 20995
rect 57563 20992 57575 20995
rect 58158 20992 58164 21004
rect 57563 20964 58164 20992
rect 57563 20961 57575 20964
rect 57517 20955 57575 20961
rect 58158 20952 58164 20964
rect 58216 20952 58222 21004
rect 51092 20896 58020 20924
rect 50801 20887 50859 20893
rect 36262 20856 36268 20868
rect 30576 20828 36268 20856
rect 36262 20816 36268 20828
rect 36320 20816 36326 20868
rect 38105 20859 38163 20865
rect 38105 20825 38117 20859
rect 38151 20856 38163 20859
rect 57330 20856 57336 20868
rect 38151 20828 57336 20856
rect 38151 20825 38163 20828
rect 38105 20819 38163 20825
rect 57330 20816 57336 20828
rect 57388 20816 57394 20868
rect 57992 20865 58020 20896
rect 57977 20859 58035 20865
rect 57977 20825 57989 20859
rect 58023 20825 58035 20859
rect 57977 20819 58035 20825
rect 47210 20788 47216 20800
rect 47171 20760 47216 20788
rect 47210 20748 47216 20760
rect 47268 20748 47274 20800
rect 47762 20788 47768 20800
rect 47723 20760 47768 20788
rect 47762 20748 47768 20760
rect 47820 20748 47826 20800
rect 1104 20698 58880 20720
rect 1104 20646 10614 20698
rect 10666 20646 10678 20698
rect 10730 20646 10742 20698
rect 10794 20646 10806 20698
rect 10858 20646 29878 20698
rect 29930 20646 29942 20698
rect 29994 20646 30006 20698
rect 30058 20646 30070 20698
rect 30122 20646 49142 20698
rect 49194 20646 49206 20698
rect 49258 20646 49270 20698
rect 49322 20646 49334 20698
rect 49386 20646 58880 20698
rect 1104 20624 58880 20646
rect 1581 20587 1639 20593
rect 1581 20553 1593 20587
rect 1627 20584 1639 20587
rect 4522 20584 4528 20596
rect 1627 20556 4528 20584
rect 1627 20553 1639 20556
rect 1581 20547 1639 20553
rect 4522 20544 4528 20556
rect 4580 20544 4586 20596
rect 38378 20584 38384 20596
rect 38339 20556 38384 20584
rect 38378 20544 38384 20556
rect 38436 20544 38442 20596
rect 47394 20584 47400 20596
rect 47355 20556 47400 20584
rect 47394 20544 47400 20556
rect 47452 20544 47458 20596
rect 1394 20380 1400 20392
rect 1355 20352 1400 20380
rect 1394 20340 1400 20352
rect 1452 20380 1458 20392
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1452 20352 2053 20380
rect 1452 20340 1458 20352
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 21910 20340 21916 20392
rect 21968 20380 21974 20392
rect 22554 20380 22560 20392
rect 21968 20352 22560 20380
rect 21968 20340 21974 20352
rect 22554 20340 22560 20352
rect 22612 20380 22618 20392
rect 22833 20383 22891 20389
rect 22833 20380 22845 20383
rect 22612 20352 22845 20380
rect 22612 20340 22618 20352
rect 22833 20349 22845 20352
rect 22879 20349 22891 20383
rect 23106 20380 23112 20392
rect 23067 20352 23112 20380
rect 22833 20343 22891 20349
rect 23106 20340 23112 20352
rect 23164 20340 23170 20392
rect 31294 20340 31300 20392
rect 31352 20380 31358 20392
rect 31389 20383 31447 20389
rect 31389 20380 31401 20383
rect 31352 20352 31401 20380
rect 31352 20340 31358 20352
rect 31389 20349 31401 20352
rect 31435 20349 31447 20383
rect 31389 20343 31447 20349
rect 31665 20383 31723 20389
rect 31665 20349 31677 20383
rect 31711 20380 31723 20383
rect 32214 20380 32220 20392
rect 31711 20352 32220 20380
rect 31711 20349 31723 20352
rect 31665 20343 31723 20349
rect 32214 20340 32220 20352
rect 32272 20380 32278 20392
rect 32674 20380 32680 20392
rect 32272 20352 32680 20380
rect 32272 20340 32278 20352
rect 32674 20340 32680 20352
rect 32732 20340 32738 20392
rect 36538 20380 36544 20392
rect 36499 20352 36544 20380
rect 36538 20340 36544 20352
rect 36596 20340 36602 20392
rect 36817 20383 36875 20389
rect 36817 20349 36829 20383
rect 36863 20380 36875 20383
rect 37090 20380 37096 20392
rect 36863 20352 37096 20380
rect 36863 20349 36875 20352
rect 36817 20343 36875 20349
rect 37090 20340 37096 20352
rect 37148 20340 37154 20392
rect 38473 20383 38531 20389
rect 38473 20349 38485 20383
rect 38519 20380 38531 20383
rect 38519 20352 38976 20380
rect 38519 20349 38531 20352
rect 38473 20343 38531 20349
rect 31757 20315 31815 20321
rect 31757 20281 31769 20315
rect 31803 20312 31815 20315
rect 31938 20312 31944 20324
rect 31803 20284 31944 20312
rect 31803 20281 31815 20284
rect 31757 20275 31815 20281
rect 31938 20272 31944 20284
rect 31996 20272 32002 20324
rect 38948 20256 38976 20352
rect 2682 20244 2688 20256
rect 2643 20216 2688 20244
rect 2682 20204 2688 20216
rect 2740 20204 2746 20256
rect 23290 20244 23296 20256
rect 23251 20216 23296 20244
rect 23290 20204 23296 20216
rect 23348 20204 23354 20256
rect 36354 20244 36360 20256
rect 36315 20216 36360 20244
rect 36354 20204 36360 20216
rect 36412 20204 36418 20256
rect 38930 20244 38936 20256
rect 38891 20216 38936 20244
rect 38930 20204 38936 20216
rect 38988 20204 38994 20256
rect 1104 20154 58880 20176
rect 1104 20102 20246 20154
rect 20298 20102 20310 20154
rect 20362 20102 20374 20154
rect 20426 20102 20438 20154
rect 20490 20102 39510 20154
rect 39562 20102 39574 20154
rect 39626 20102 39638 20154
rect 39690 20102 39702 20154
rect 39754 20102 58880 20154
rect 1104 20080 58880 20102
rect 1578 20000 1584 20052
rect 1636 20040 1642 20052
rect 2409 20043 2467 20049
rect 2409 20040 2421 20043
rect 1636 20012 2421 20040
rect 1636 20000 1642 20012
rect 2409 20009 2421 20012
rect 2455 20009 2467 20043
rect 2409 20003 2467 20009
rect 2498 20000 2504 20052
rect 2556 20040 2562 20052
rect 3053 20043 3111 20049
rect 3053 20040 3065 20043
rect 2556 20012 3065 20040
rect 2556 20000 2562 20012
rect 3053 20009 3065 20012
rect 3099 20009 3111 20043
rect 3053 20003 3111 20009
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 15933 20043 15991 20049
rect 15933 20040 15945 20043
rect 15896 20012 15945 20040
rect 15896 20000 15902 20012
rect 15933 20009 15945 20012
rect 15979 20009 15991 20043
rect 15933 20003 15991 20009
rect 17865 20043 17923 20049
rect 17865 20009 17877 20043
rect 17911 20009 17923 20043
rect 21910 20040 21916 20052
rect 21871 20012 21916 20040
rect 17865 20003 17923 20009
rect 2332 19944 16804 19972
rect 2332 19916 2360 19944
rect 2314 19904 2320 19916
rect 2227 19876 2320 19904
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 2501 19907 2559 19913
rect 2501 19873 2513 19907
rect 2547 19904 2559 19907
rect 2682 19904 2688 19916
rect 2547 19876 2688 19904
rect 2547 19873 2559 19876
rect 2501 19867 2559 19873
rect 2682 19864 2688 19876
rect 2740 19904 2746 19916
rect 2961 19907 3019 19913
rect 2961 19904 2973 19907
rect 2740 19876 2973 19904
rect 2740 19864 2746 19876
rect 2961 19873 2973 19876
rect 3007 19873 3019 19907
rect 2961 19867 3019 19873
rect 3145 19907 3203 19913
rect 3145 19873 3157 19907
rect 3191 19904 3203 19907
rect 8754 19904 8760 19916
rect 3191 19876 8760 19904
rect 3191 19873 3203 19876
rect 3145 19867 3203 19873
rect 2976 19836 3004 19867
rect 8754 19864 8760 19876
rect 8812 19904 8818 19916
rect 16776 19913 16804 19944
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 8812 19876 15853 19904
rect 8812 19864 8818 19876
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 15841 19867 15899 19873
rect 16025 19907 16083 19913
rect 16025 19873 16037 19907
rect 16071 19873 16083 19907
rect 16025 19867 16083 19873
rect 16761 19907 16819 19913
rect 16761 19873 16773 19907
rect 16807 19873 16819 19907
rect 16761 19867 16819 19873
rect 17773 19907 17831 19913
rect 17773 19873 17785 19907
rect 17819 19873 17831 19907
rect 17773 19867 17831 19873
rect 16040 19836 16068 19867
rect 16206 19836 16212 19848
rect 2976 19808 4016 19836
rect 16040 19808 16212 19836
rect 3988 19712 4016 19808
rect 16206 19796 16212 19808
rect 16264 19836 16270 19848
rect 17788 19836 17816 19867
rect 16264 19808 17816 19836
rect 17880 19836 17908 20003
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 23290 20000 23296 20052
rect 23348 20040 23354 20052
rect 57790 20040 57796 20052
rect 23348 20012 57796 20040
rect 23348 20000 23354 20012
rect 57790 20000 57796 20012
rect 57848 20000 57854 20052
rect 32674 19972 32680 19984
rect 32635 19944 32680 19972
rect 32674 19932 32680 19944
rect 32732 19932 32738 19984
rect 36449 19975 36507 19981
rect 36449 19941 36461 19975
rect 36495 19972 36507 19975
rect 36495 19944 37320 19972
rect 36495 19941 36507 19944
rect 36449 19935 36507 19941
rect 21818 19904 21824 19916
rect 21779 19876 21824 19904
rect 21818 19864 21824 19876
rect 21876 19904 21882 19916
rect 22465 19907 22523 19913
rect 22465 19904 22477 19907
rect 21876 19876 22477 19904
rect 21876 19864 21882 19876
rect 22465 19873 22477 19876
rect 22511 19873 22523 19907
rect 31110 19904 31116 19916
rect 31071 19876 31116 19904
rect 22465 19867 22523 19873
rect 31110 19864 31116 19876
rect 31168 19864 31174 19916
rect 31386 19904 31392 19916
rect 31347 19876 31392 19904
rect 31386 19864 31392 19876
rect 31444 19904 31450 19916
rect 32033 19907 32091 19913
rect 32033 19904 32045 19907
rect 31444 19876 32045 19904
rect 31444 19864 31450 19876
rect 32033 19873 32045 19876
rect 32079 19873 32091 19907
rect 32033 19867 32091 19873
rect 32125 19907 32183 19913
rect 32125 19873 32137 19907
rect 32171 19904 32183 19907
rect 32214 19904 32220 19916
rect 32171 19876 32220 19904
rect 32171 19873 32183 19876
rect 32125 19867 32183 19873
rect 32214 19864 32220 19876
rect 32272 19864 32278 19916
rect 32398 19864 32404 19916
rect 32456 19904 32462 19916
rect 32585 19907 32643 19913
rect 32585 19904 32597 19907
rect 32456 19876 32597 19904
rect 32456 19864 32462 19876
rect 32585 19873 32597 19876
rect 32631 19873 32643 19907
rect 32585 19867 32643 19873
rect 35802 19864 35808 19916
rect 35860 19904 35866 19916
rect 36357 19907 36415 19913
rect 36357 19904 36369 19907
rect 35860 19876 36369 19904
rect 35860 19864 35866 19876
rect 36357 19873 36369 19876
rect 36403 19873 36415 19907
rect 36357 19867 36415 19873
rect 36538 19864 36544 19916
rect 36596 19904 36602 19916
rect 37292 19913 37320 19944
rect 37001 19907 37059 19913
rect 37001 19904 37013 19907
rect 36596 19876 37013 19904
rect 36596 19864 36602 19876
rect 37001 19873 37013 19876
rect 37047 19873 37059 19907
rect 37001 19867 37059 19873
rect 37277 19907 37335 19913
rect 37277 19873 37289 19907
rect 37323 19904 37335 19907
rect 38010 19904 38016 19916
rect 37323 19876 38016 19904
rect 37323 19873 37335 19876
rect 37277 19867 37335 19873
rect 38010 19864 38016 19876
rect 38068 19864 38074 19916
rect 57977 19907 58035 19913
rect 57977 19904 57989 19907
rect 57348 19876 57989 19904
rect 54938 19836 54944 19848
rect 17880 19808 54944 19836
rect 16264 19796 16270 19808
rect 17788 19768 17816 19808
rect 54938 19796 54944 19808
rect 54996 19796 55002 19848
rect 31389 19771 31447 19777
rect 17788 19740 18552 19768
rect 3970 19700 3976 19712
rect 3931 19672 3976 19700
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 18524 19709 18552 19740
rect 31389 19737 31401 19771
rect 31435 19768 31447 19771
rect 31478 19768 31484 19780
rect 31435 19740 31484 19768
rect 31435 19737 31447 19740
rect 31389 19731 31447 19737
rect 31478 19728 31484 19740
rect 31536 19728 31542 19780
rect 57348 19777 57376 19876
rect 57977 19873 57989 19876
rect 58023 19873 58035 19907
rect 57977 19867 58035 19873
rect 37277 19771 37335 19777
rect 37277 19737 37289 19771
rect 37323 19768 37335 19771
rect 57333 19771 57391 19777
rect 57333 19768 57345 19771
rect 37323 19740 57345 19768
rect 37323 19737 37335 19740
rect 37277 19731 37335 19737
rect 57333 19737 57345 19740
rect 57379 19737 57391 19771
rect 58158 19768 58164 19780
rect 58119 19740 58164 19768
rect 57333 19731 57391 19737
rect 58158 19728 58164 19740
rect 58216 19728 58222 19780
rect 18509 19703 18567 19709
rect 18509 19669 18521 19703
rect 18555 19700 18567 19703
rect 19334 19700 19340 19712
rect 18555 19672 19340 19700
rect 18555 19669 18567 19672
rect 18509 19663 18567 19669
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 35802 19700 35808 19712
rect 35763 19672 35808 19700
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 1104 19610 58880 19632
rect 1104 19558 10614 19610
rect 10666 19558 10678 19610
rect 10730 19558 10742 19610
rect 10794 19558 10806 19610
rect 10858 19558 29878 19610
rect 29930 19558 29942 19610
rect 29994 19558 30006 19610
rect 30058 19558 30070 19610
rect 30122 19558 49142 19610
rect 49194 19558 49206 19610
rect 49258 19558 49270 19610
rect 49322 19558 49334 19610
rect 49386 19558 58880 19610
rect 1104 19536 58880 19558
rect 2314 19496 2320 19508
rect 2275 19468 2320 19496
rect 2314 19456 2320 19468
rect 2372 19456 2378 19508
rect 3970 19456 3976 19508
rect 4028 19496 4034 19508
rect 25682 19496 25688 19508
rect 4028 19468 25688 19496
rect 4028 19456 4034 19468
rect 25682 19456 25688 19468
rect 25740 19456 25746 19508
rect 7006 19388 7012 19440
rect 7064 19428 7070 19440
rect 35802 19428 35808 19440
rect 7064 19400 35808 19428
rect 7064 19388 7070 19400
rect 35802 19388 35808 19400
rect 35860 19388 35866 19440
rect 16206 19360 16212 19372
rect 16167 19332 16212 19360
rect 16206 19320 16212 19332
rect 16264 19320 16270 19372
rect 1394 19292 1400 19304
rect 1355 19264 1400 19292
rect 1394 19252 1400 19264
rect 1452 19252 1458 19304
rect 2222 19292 2228 19304
rect 2183 19264 2228 19292
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 8662 19292 8668 19304
rect 8623 19264 8668 19292
rect 8662 19252 8668 19264
rect 8720 19252 8726 19304
rect 8754 19252 8760 19304
rect 8812 19292 8818 19304
rect 8812 19264 8857 19292
rect 8812 19252 8818 19264
rect 57977 19227 58035 19233
rect 57977 19224 57989 19227
rect 57348 19196 57989 19224
rect 57348 19168 57376 19196
rect 57977 19193 57989 19196
rect 58023 19193 58035 19227
rect 58158 19224 58164 19236
rect 58119 19196 58164 19224
rect 57977 19187 58035 19193
rect 58158 19184 58164 19196
rect 58216 19184 58222 19236
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 32214 19116 32220 19168
rect 32272 19156 32278 19168
rect 32769 19159 32827 19165
rect 32769 19156 32781 19159
rect 32272 19128 32781 19156
rect 32272 19116 32278 19128
rect 32769 19125 32781 19128
rect 32815 19156 32827 19159
rect 45738 19156 45744 19168
rect 32815 19128 45744 19156
rect 32815 19125 32827 19128
rect 32769 19119 32827 19125
rect 45738 19116 45744 19128
rect 45796 19116 45802 19168
rect 57330 19156 57336 19168
rect 57291 19128 57336 19156
rect 57330 19116 57336 19128
rect 57388 19116 57394 19168
rect 1104 19066 58880 19088
rect 1104 19014 20246 19066
rect 20298 19014 20310 19066
rect 20362 19014 20374 19066
rect 20426 19014 20438 19066
rect 20490 19014 39510 19066
rect 39562 19014 39574 19066
rect 39626 19014 39638 19066
rect 39690 19014 39702 19066
rect 39754 19014 58880 19066
rect 1104 18992 58880 19014
rect 1394 18952 1400 18964
rect 1355 18924 1400 18952
rect 1394 18912 1400 18924
rect 1452 18912 1458 18964
rect 1578 18912 1584 18964
rect 1636 18952 1642 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 1636 18924 2329 18952
rect 1636 18912 1642 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 26513 18955 26571 18961
rect 26513 18921 26525 18955
rect 26559 18952 26571 18955
rect 26602 18952 26608 18964
rect 26559 18924 26608 18952
rect 26559 18921 26571 18924
rect 26513 18915 26571 18921
rect 26602 18912 26608 18924
rect 26660 18912 26666 18964
rect 25774 18776 25780 18828
rect 25832 18816 25838 18828
rect 26421 18819 26479 18825
rect 26421 18816 26433 18819
rect 25832 18788 26433 18816
rect 25832 18776 25838 18788
rect 26421 18785 26433 18788
rect 26467 18785 26479 18819
rect 26421 18779 26479 18785
rect 26605 18819 26663 18825
rect 26605 18785 26617 18819
rect 26651 18816 26663 18819
rect 26786 18816 26792 18828
rect 26651 18788 26792 18816
rect 26651 18785 26663 18788
rect 26605 18779 26663 18785
rect 26786 18776 26792 18788
rect 26844 18816 26850 18828
rect 27062 18816 27068 18828
rect 26844 18788 27068 18816
rect 26844 18776 26850 18788
rect 27062 18776 27068 18788
rect 27120 18816 27126 18828
rect 27433 18819 27491 18825
rect 27433 18816 27445 18819
rect 27120 18788 27445 18816
rect 27120 18776 27126 18788
rect 27433 18785 27445 18788
rect 27479 18785 27491 18819
rect 27890 18816 27896 18828
rect 27851 18788 27896 18816
rect 27433 18779 27491 18785
rect 27890 18776 27896 18788
rect 27948 18776 27954 18828
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18717 2467 18751
rect 2409 18711 2467 18717
rect 2424 18680 2452 18711
rect 2498 18708 2504 18760
rect 2556 18748 2562 18760
rect 2593 18751 2651 18757
rect 2593 18748 2605 18751
rect 2556 18720 2605 18748
rect 2556 18708 2562 18720
rect 2593 18717 2605 18720
rect 2639 18748 2651 18751
rect 4154 18748 4160 18760
rect 2639 18720 4160 18748
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 4154 18708 4160 18720
rect 4212 18708 4218 18760
rect 28169 18751 28227 18757
rect 28169 18717 28181 18751
rect 28215 18748 28227 18751
rect 44450 18748 44456 18760
rect 28215 18720 44456 18748
rect 28215 18717 28227 18720
rect 28169 18711 28227 18717
rect 44450 18708 44456 18720
rect 44508 18708 44514 18760
rect 3237 18683 3295 18689
rect 3237 18680 3249 18683
rect 2424 18652 3249 18680
rect 3237 18649 3249 18652
rect 3283 18680 3295 18683
rect 34882 18680 34888 18692
rect 3283 18652 34888 18680
rect 3283 18649 3295 18652
rect 3237 18643 3295 18649
rect 34882 18640 34888 18652
rect 34940 18640 34946 18692
rect 42334 18640 42340 18692
rect 42392 18680 42398 18692
rect 57146 18680 57152 18692
rect 42392 18652 57152 18680
rect 42392 18640 42398 18652
rect 57146 18640 57152 18652
rect 57204 18640 57210 18692
rect 1949 18615 2007 18621
rect 1949 18581 1961 18615
rect 1995 18612 2007 18615
rect 2038 18612 2044 18624
rect 1995 18584 2044 18612
rect 1995 18581 2007 18584
rect 1949 18575 2007 18581
rect 2038 18572 2044 18584
rect 2096 18572 2102 18624
rect 1104 18522 58880 18544
rect 1104 18470 10614 18522
rect 10666 18470 10678 18522
rect 10730 18470 10742 18522
rect 10794 18470 10806 18522
rect 10858 18470 29878 18522
rect 29930 18470 29942 18522
rect 29994 18470 30006 18522
rect 30058 18470 30070 18522
rect 30122 18470 49142 18522
rect 49194 18470 49206 18522
rect 49258 18470 49270 18522
rect 49322 18470 49334 18522
rect 49386 18470 58880 18522
rect 1104 18448 58880 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 2222 18408 2228 18420
rect 1627 18380 2228 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 2222 18368 2228 18380
rect 2280 18368 2286 18420
rect 2498 18368 2504 18420
rect 2556 18408 2562 18420
rect 2593 18411 2651 18417
rect 2593 18408 2605 18411
rect 2556 18380 2605 18408
rect 2556 18368 2562 18380
rect 2593 18377 2605 18380
rect 2639 18377 2651 18411
rect 2593 18371 2651 18377
rect 1394 18204 1400 18216
rect 1355 18176 1400 18204
rect 1394 18164 1400 18176
rect 1452 18204 1458 18216
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1452 18176 2053 18204
rect 1452 18164 1458 18176
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 1104 17978 58880 18000
rect 1104 17926 20246 17978
rect 20298 17926 20310 17978
rect 20362 17926 20374 17978
rect 20426 17926 20438 17978
rect 20490 17926 39510 17978
rect 39562 17926 39574 17978
rect 39626 17926 39638 17978
rect 39690 17926 39702 17978
rect 39754 17926 58880 17978
rect 1104 17904 58880 17926
rect 27062 17864 27068 17876
rect 27023 17836 27068 17864
rect 27062 17824 27068 17836
rect 27120 17824 27126 17876
rect 27614 17824 27620 17876
rect 27672 17864 27678 17876
rect 27893 17867 27951 17873
rect 27893 17864 27905 17867
rect 27672 17836 27905 17864
rect 27672 17824 27678 17836
rect 27893 17833 27905 17836
rect 27939 17833 27951 17867
rect 27893 17827 27951 17833
rect 55217 17867 55275 17873
rect 55217 17833 55229 17867
rect 55263 17864 55275 17867
rect 57977 17867 58035 17873
rect 57977 17864 57989 17867
rect 55263 17836 57989 17864
rect 55263 17833 55275 17836
rect 55217 17827 55275 17833
rect 57977 17833 57989 17836
rect 58023 17833 58035 17867
rect 57977 17827 58035 17833
rect 25406 17756 25412 17808
rect 25464 17796 25470 17808
rect 26329 17799 26387 17805
rect 26329 17796 26341 17799
rect 25464 17768 26341 17796
rect 25464 17756 25470 17768
rect 26329 17765 26341 17768
rect 26375 17796 26387 17799
rect 27801 17799 27859 17805
rect 27801 17796 27813 17799
rect 26375 17768 27813 17796
rect 26375 17765 26387 17768
rect 26329 17759 26387 17765
rect 27801 17765 27813 17768
rect 27847 17765 27859 17799
rect 27801 17759 27859 17765
rect 1394 17728 1400 17740
rect 1355 17700 1400 17728
rect 1394 17688 1400 17700
rect 1452 17688 1458 17740
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 2222 17728 2228 17740
rect 1627 17700 2228 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 27249 17731 27307 17737
rect 27249 17697 27261 17731
rect 27295 17697 27307 17731
rect 27249 17691 27307 17697
rect 26513 17663 26571 17669
rect 26513 17629 26525 17663
rect 26559 17660 26571 17663
rect 26602 17660 26608 17672
rect 26559 17632 26608 17660
rect 26559 17629 26571 17632
rect 26513 17623 26571 17629
rect 26602 17620 26608 17632
rect 26660 17660 26666 17672
rect 27264 17660 27292 17691
rect 28718 17688 28724 17740
rect 28776 17728 28782 17740
rect 54205 17731 54263 17737
rect 54205 17728 54217 17731
rect 28776 17700 54217 17728
rect 28776 17688 28782 17700
rect 54205 17697 54217 17700
rect 54251 17728 54263 17731
rect 55125 17731 55183 17737
rect 55125 17728 55137 17731
rect 54251 17700 55137 17728
rect 54251 17697 54263 17700
rect 54205 17691 54263 17697
rect 55125 17697 55137 17700
rect 55171 17697 55183 17731
rect 55125 17691 55183 17697
rect 57517 17731 57575 17737
rect 57517 17697 57529 17731
rect 57563 17728 57575 17731
rect 58158 17728 58164 17740
rect 57563 17700 58164 17728
rect 57563 17697 57575 17700
rect 57517 17691 57575 17697
rect 58158 17688 58164 17700
rect 58216 17688 58222 17740
rect 36262 17660 36268 17672
rect 26660 17632 36268 17660
rect 26660 17620 26666 17632
rect 36262 17620 36268 17632
rect 36320 17620 36326 17672
rect 54386 17620 54392 17672
rect 54444 17660 54450 17672
rect 55309 17663 55367 17669
rect 55309 17660 55321 17663
rect 54444 17632 55321 17660
rect 54444 17620 54450 17632
rect 55309 17629 55321 17632
rect 55355 17629 55367 17663
rect 55309 17623 55367 17629
rect 2222 17524 2228 17536
rect 2183 17496 2228 17524
rect 2222 17484 2228 17496
rect 2280 17484 2286 17536
rect 54757 17527 54815 17533
rect 54757 17493 54769 17527
rect 54803 17524 54815 17527
rect 54938 17524 54944 17536
rect 54803 17496 54944 17524
rect 54803 17493 54815 17496
rect 54757 17487 54815 17493
rect 54938 17484 54944 17496
rect 54996 17484 55002 17536
rect 1104 17434 58880 17456
rect 1104 17382 10614 17434
rect 10666 17382 10678 17434
rect 10730 17382 10742 17434
rect 10794 17382 10806 17434
rect 10858 17382 29878 17434
rect 29930 17382 29942 17434
rect 29994 17382 30006 17434
rect 30058 17382 30070 17434
rect 30122 17382 49142 17434
rect 49194 17382 49206 17434
rect 49258 17382 49270 17434
rect 49322 17382 49334 17434
rect 49386 17382 58880 17434
rect 1104 17360 58880 17382
rect 25406 17320 25412 17332
rect 25367 17292 25412 17320
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 54386 17320 54392 17332
rect 54347 17292 54392 17320
rect 54386 17280 54392 17292
rect 54444 17280 54450 17332
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 19392 17156 26065 17184
rect 19392 17144 19398 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 8018 17116 8024 17128
rect 7979 17088 8024 17116
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 24857 17119 24915 17125
rect 24857 17085 24869 17119
rect 24903 17116 24915 17119
rect 25314 17116 25320 17128
rect 24903 17088 25320 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 25314 17076 25320 17088
rect 25372 17076 25378 17128
rect 26602 17116 26608 17128
rect 26563 17088 26608 17116
rect 26602 17076 26608 17088
rect 26660 17076 26666 17128
rect 36262 17116 36268 17128
rect 36223 17088 36268 17116
rect 36262 17076 36268 17088
rect 36320 17076 36326 17128
rect 57882 17116 57888 17128
rect 57843 17088 57888 17116
rect 57882 17076 57888 17088
rect 57940 17076 57946 17128
rect 36446 17008 36452 17060
rect 36504 17048 36510 17060
rect 36541 17051 36599 17057
rect 36541 17048 36553 17051
rect 36504 17020 36553 17048
rect 36504 17008 36510 17020
rect 36541 17017 36553 17020
rect 36587 17048 36599 17051
rect 37642 17048 37648 17060
rect 36587 17020 37648 17048
rect 36587 17017 36599 17020
rect 36541 17011 36599 17017
rect 37642 17008 37648 17020
rect 37700 17008 37706 17060
rect 57425 17051 57483 17057
rect 57425 17017 57437 17051
rect 57471 17048 57483 17051
rect 58066 17048 58072 17060
rect 57471 17020 58072 17048
rect 57471 17017 57483 17020
rect 57425 17011 57483 17017
rect 58066 17008 58072 17020
rect 58124 17008 58130 17060
rect 8113 16983 8171 16989
rect 8113 16949 8125 16983
rect 8159 16980 8171 16983
rect 8478 16980 8484 16992
rect 8159 16952 8484 16980
rect 8159 16949 8171 16952
rect 8113 16943 8171 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 1104 16890 58880 16912
rect 1104 16838 20246 16890
rect 20298 16838 20310 16890
rect 20362 16838 20374 16890
rect 20426 16838 20438 16890
rect 20490 16838 39510 16890
rect 39562 16838 39574 16890
rect 39626 16838 39638 16890
rect 39690 16838 39702 16890
rect 39754 16838 58880 16890
rect 1104 16816 58880 16838
rect 10318 16776 10324 16788
rect 10279 16748 10324 16776
rect 10318 16736 10324 16748
rect 10376 16736 10382 16788
rect 21269 16779 21327 16785
rect 21269 16745 21281 16779
rect 21315 16776 21327 16779
rect 21358 16776 21364 16788
rect 21315 16748 21364 16776
rect 21315 16745 21327 16748
rect 21269 16739 21327 16745
rect 21358 16736 21364 16748
rect 21416 16776 21422 16788
rect 22738 16776 22744 16788
rect 21416 16748 22744 16776
rect 21416 16736 21422 16748
rect 1394 16600 1400 16652
rect 1452 16640 1458 16652
rect 1489 16643 1547 16649
rect 1489 16640 1501 16643
rect 1452 16612 1501 16640
rect 1452 16600 1458 16612
rect 1489 16609 1501 16612
rect 1535 16609 1547 16643
rect 1489 16603 1547 16609
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 10321 16643 10379 16649
rect 10321 16640 10333 16643
rect 8536 16612 10333 16640
rect 8536 16600 8542 16612
rect 10321 16609 10333 16612
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 10597 16643 10655 16649
rect 10597 16609 10609 16643
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 21085 16643 21143 16649
rect 21085 16609 21097 16643
rect 21131 16640 21143 16643
rect 21174 16640 21180 16652
rect 21131 16612 21180 16640
rect 21131 16609 21143 16612
rect 21085 16603 21143 16609
rect 10612 16572 10640 16603
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21744 16649 21772 16748
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 22005 16711 22063 16717
rect 22005 16708 22017 16711
rect 21928 16680 22017 16708
rect 21729 16643 21787 16649
rect 21729 16609 21741 16643
rect 21775 16609 21787 16643
rect 21729 16603 21787 16609
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 10612 16544 11161 16572
rect 11149 16541 11161 16544
rect 11195 16572 11207 16575
rect 14366 16572 14372 16584
rect 11195 16544 14372 16572
rect 11195 16541 11207 16544
rect 11149 16535 11207 16541
rect 14366 16532 14372 16544
rect 14424 16572 14430 16584
rect 21928 16572 21956 16680
rect 22005 16677 22017 16680
rect 22051 16708 22063 16711
rect 29454 16708 29460 16720
rect 22051 16680 28672 16708
rect 22051 16677 22063 16680
rect 22005 16671 22063 16677
rect 22738 16640 22744 16652
rect 22699 16612 22744 16640
rect 22738 16600 22744 16612
rect 22796 16600 22802 16652
rect 25406 16600 25412 16652
rect 25464 16640 25470 16652
rect 25685 16643 25743 16649
rect 25685 16640 25697 16643
rect 25464 16612 25697 16640
rect 25464 16600 25470 16612
rect 25685 16609 25697 16612
rect 25731 16609 25743 16643
rect 26786 16640 26792 16652
rect 26747 16612 26792 16640
rect 25685 16603 25743 16609
rect 26786 16600 26792 16612
rect 26844 16600 26850 16652
rect 28644 16649 28672 16680
rect 29196 16680 29460 16708
rect 29196 16649 29224 16680
rect 29454 16668 29460 16680
rect 29512 16668 29518 16720
rect 57882 16708 57888 16720
rect 42490 16680 57888 16708
rect 28629 16643 28687 16649
rect 28629 16609 28641 16643
rect 28675 16640 28687 16643
rect 29181 16643 29239 16649
rect 29181 16640 29193 16643
rect 28675 16612 29193 16640
rect 28675 16609 28687 16612
rect 28629 16603 28687 16609
rect 29181 16609 29193 16612
rect 29227 16609 29239 16643
rect 29362 16640 29368 16652
rect 29323 16612 29368 16640
rect 29181 16603 29239 16609
rect 29362 16600 29368 16612
rect 29420 16600 29426 16652
rect 37090 16640 37096 16652
rect 37003 16612 37096 16640
rect 37090 16600 37096 16612
rect 37148 16640 37154 16652
rect 38013 16643 38071 16649
rect 38013 16640 38025 16643
rect 37148 16612 38025 16640
rect 37148 16600 37154 16612
rect 38013 16609 38025 16612
rect 38059 16609 38071 16643
rect 38013 16603 38071 16609
rect 37369 16575 37427 16581
rect 14424 16544 21956 16572
rect 22388 16544 29638 16572
rect 14424 16532 14430 16544
rect 13538 16464 13544 16516
rect 13596 16504 13602 16516
rect 22388 16504 22416 16544
rect 25314 16504 25320 16516
rect 13596 16476 22416 16504
rect 22480 16476 25320 16504
rect 13596 16464 13602 16476
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 20625 16439 20683 16445
rect 20625 16405 20637 16439
rect 20671 16436 20683 16439
rect 21174 16436 21180 16448
rect 20671 16408 21180 16436
rect 20671 16405 20683 16408
rect 20625 16399 20683 16405
rect 21174 16396 21180 16408
rect 21232 16436 21238 16448
rect 22480 16436 22508 16476
rect 25314 16464 25320 16476
rect 25372 16504 25378 16516
rect 25372 16476 27016 16504
rect 25372 16464 25378 16476
rect 21232 16408 22508 16436
rect 23017 16439 23075 16445
rect 21232 16396 21238 16408
rect 23017 16405 23029 16439
rect 23063 16436 23075 16439
rect 23290 16436 23296 16448
rect 23063 16408 23296 16436
rect 23063 16405 23075 16408
rect 23017 16399 23075 16405
rect 23290 16396 23296 16408
rect 23348 16396 23354 16448
rect 24394 16396 24400 16448
rect 24452 16436 24458 16448
rect 25501 16439 25559 16445
rect 25501 16436 25513 16439
rect 24452 16408 25513 16436
rect 24452 16396 24458 16408
rect 25501 16405 25513 16408
rect 25547 16405 25559 16439
rect 25501 16399 25559 16405
rect 26510 16396 26516 16448
rect 26568 16436 26574 16448
rect 26605 16439 26663 16445
rect 26605 16436 26617 16439
rect 26568 16408 26617 16436
rect 26568 16396 26574 16408
rect 26605 16405 26617 16408
rect 26651 16436 26663 16439
rect 26878 16436 26884 16448
rect 26651 16408 26884 16436
rect 26651 16405 26663 16408
rect 26605 16399 26663 16405
rect 26878 16396 26884 16408
rect 26936 16396 26942 16448
rect 26988 16436 27016 16476
rect 29270 16464 29276 16516
rect 29328 16504 29334 16516
rect 29365 16507 29423 16513
rect 29365 16504 29377 16507
rect 29328 16476 29377 16504
rect 29328 16464 29334 16476
rect 29365 16473 29377 16476
rect 29411 16473 29423 16507
rect 29610 16504 29638 16544
rect 37369 16541 37381 16575
rect 37415 16572 37427 16575
rect 37458 16572 37464 16584
rect 37415 16544 37464 16572
rect 37415 16541 37427 16544
rect 37369 16535 37427 16541
rect 37458 16532 37464 16544
rect 37516 16532 37522 16584
rect 37550 16532 37556 16584
rect 37608 16572 37614 16584
rect 42490 16572 42518 16680
rect 57882 16668 57888 16680
rect 57940 16668 57946 16720
rect 44637 16643 44695 16649
rect 44637 16609 44649 16643
rect 44683 16640 44695 16643
rect 57974 16640 57980 16652
rect 44683 16612 45232 16640
rect 57935 16612 57980 16640
rect 44683 16609 44695 16612
rect 44637 16603 44695 16609
rect 37608 16544 42518 16572
rect 37608 16532 37614 16544
rect 40862 16504 40868 16516
rect 29610 16476 40868 16504
rect 29365 16467 29423 16473
rect 40862 16464 40868 16476
rect 40920 16464 40926 16516
rect 29546 16436 29552 16448
rect 26988 16408 29552 16436
rect 29546 16396 29552 16408
rect 29604 16396 29610 16448
rect 38194 16436 38200 16448
rect 38155 16408 38200 16436
rect 38194 16396 38200 16408
rect 38252 16396 38258 16448
rect 44542 16436 44548 16448
rect 44503 16408 44548 16436
rect 44542 16396 44548 16408
rect 44600 16396 44606 16448
rect 45204 16445 45232 16612
rect 57974 16600 57980 16612
rect 58032 16600 58038 16652
rect 58158 16504 58164 16516
rect 58119 16476 58164 16504
rect 58158 16464 58164 16476
rect 58216 16464 58222 16516
rect 45189 16439 45247 16445
rect 45189 16405 45201 16439
rect 45235 16436 45247 16439
rect 57698 16436 57704 16448
rect 45235 16408 57704 16436
rect 45235 16405 45247 16408
rect 45189 16399 45247 16405
rect 57698 16396 57704 16408
rect 57756 16396 57762 16448
rect 1104 16346 58880 16368
rect 1104 16294 10614 16346
rect 10666 16294 10678 16346
rect 10730 16294 10742 16346
rect 10794 16294 10806 16346
rect 10858 16294 29878 16346
rect 29930 16294 29942 16346
rect 29994 16294 30006 16346
rect 30058 16294 30070 16346
rect 30122 16294 49142 16346
rect 49194 16294 49206 16346
rect 49258 16294 49270 16346
rect 49322 16294 49334 16346
rect 49386 16294 58880 16346
rect 1104 16272 58880 16294
rect 1394 16232 1400 16244
rect 1355 16204 1400 16232
rect 1394 16192 1400 16204
rect 1452 16192 1458 16244
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 29730 16232 29736 16244
rect 1636 16204 29736 16232
rect 1636 16192 1642 16204
rect 29730 16192 29736 16204
rect 29788 16192 29794 16244
rect 29917 16235 29975 16241
rect 29917 16201 29929 16235
rect 29963 16232 29975 16235
rect 30190 16232 30196 16244
rect 29963 16204 30196 16232
rect 29963 16201 29975 16204
rect 29917 16195 29975 16201
rect 30190 16192 30196 16204
rect 30248 16232 30254 16244
rect 37090 16232 37096 16244
rect 30248 16204 37096 16232
rect 30248 16192 30254 16204
rect 37090 16192 37096 16204
rect 37148 16192 37154 16244
rect 17862 16124 17868 16176
rect 17920 16164 17926 16176
rect 18325 16167 18383 16173
rect 18325 16164 18337 16167
rect 17920 16136 18337 16164
rect 17920 16124 17926 16136
rect 18325 16133 18337 16136
rect 18371 16133 18383 16167
rect 18325 16127 18383 16133
rect 25682 16124 25688 16176
rect 25740 16164 25746 16176
rect 25961 16167 26019 16173
rect 25961 16164 25973 16167
rect 25740 16136 25973 16164
rect 25740 16124 25746 16136
rect 25961 16133 25973 16136
rect 26007 16133 26019 16167
rect 25961 16127 26019 16133
rect 29178 16124 29184 16176
rect 29236 16164 29242 16176
rect 29365 16167 29423 16173
rect 29365 16164 29377 16167
rect 29236 16136 29377 16164
rect 29236 16124 29242 16136
rect 29365 16133 29377 16136
rect 29411 16133 29423 16167
rect 57330 16164 57336 16176
rect 29365 16127 29423 16133
rect 29840 16136 57336 16164
rect 21082 16096 21088 16108
rect 21043 16068 21088 16096
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16096 23351 16099
rect 29840 16096 29868 16136
rect 57330 16124 57336 16136
rect 57388 16124 57394 16176
rect 37550 16096 37556 16108
rect 23339 16068 29868 16096
rect 36004 16068 37556 16096
rect 23339 16065 23351 16068
rect 23293 16059 23351 16065
rect 36004 16040 36032 16068
rect 37550 16056 37556 16068
rect 37608 16056 37614 16108
rect 38194 16056 38200 16108
rect 38252 16096 38258 16108
rect 40862 16096 40868 16108
rect 38252 16068 40724 16096
rect 40823 16068 40868 16096
rect 38252 16056 38258 16068
rect 8478 16028 8484 16040
rect 8439 16000 8484 16028
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 18509 16031 18567 16037
rect 18509 15997 18521 16031
rect 18555 16028 18567 16031
rect 18782 16028 18788 16040
rect 18555 16000 18788 16028
rect 18555 15997 18567 16000
rect 18509 15991 18567 15997
rect 8294 15920 8300 15972
rect 8352 15960 8358 15972
rect 8389 15963 8447 15969
rect 8389 15960 8401 15963
rect 8352 15932 8401 15960
rect 8352 15920 8358 15932
rect 8389 15929 8401 15932
rect 8435 15929 8447 15963
rect 8772 15960 8800 15991
rect 18782 15988 18788 16000
rect 18840 15988 18846 16040
rect 21358 16028 21364 16040
rect 21319 16000 21364 16028
rect 21358 15988 21364 16000
rect 21416 15988 21422 16040
rect 23198 16028 23204 16040
rect 23159 16000 23204 16028
rect 23198 15988 23204 16000
rect 23256 15988 23262 16040
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 25498 16028 25504 16040
rect 23799 16000 25504 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 9309 15963 9367 15969
rect 9309 15960 9321 15963
rect 8772 15932 9321 15960
rect 8389 15923 8447 15929
rect 9309 15929 9321 15932
rect 9355 15960 9367 15963
rect 15470 15960 15476 15972
rect 9355 15932 15476 15960
rect 9355 15929 9367 15932
rect 9309 15923 9367 15929
rect 15470 15920 15476 15932
rect 15528 15960 15534 15972
rect 15528 15932 20622 15960
rect 15528 15920 15534 15932
rect 20594 15892 20622 15932
rect 22002 15920 22008 15972
rect 22060 15960 22066 15972
rect 22557 15963 22615 15969
rect 22557 15960 22569 15963
rect 22060 15932 22569 15960
rect 22060 15920 22066 15932
rect 22557 15929 22569 15932
rect 22603 15960 22615 15963
rect 23768 15960 23796 15991
rect 25498 15988 25504 16000
rect 25556 15988 25562 16040
rect 29086 16028 29092 16040
rect 29047 16000 29092 16028
rect 29086 15988 29092 16000
rect 29144 15988 29150 16040
rect 29270 16028 29276 16040
rect 29231 16000 29276 16028
rect 29270 15988 29276 16000
rect 29328 15988 29334 16040
rect 29546 15988 29552 16040
rect 29604 16028 29610 16040
rect 30101 16031 30159 16037
rect 30101 16028 30113 16031
rect 29604 16000 30113 16028
rect 29604 15988 29610 16000
rect 30101 15997 30113 16000
rect 30147 16028 30159 16031
rect 30561 16031 30619 16037
rect 30561 16028 30573 16031
rect 30147 16000 30573 16028
rect 30147 15997 30159 16000
rect 30101 15991 30159 15997
rect 30561 15997 30573 16000
rect 30607 15997 30619 16031
rect 35986 16028 35992 16040
rect 35899 16000 35992 16028
rect 30561 15991 30619 15997
rect 35986 15988 35992 16000
rect 36044 15988 36050 16040
rect 36262 15988 36268 16040
rect 36320 16028 36326 16040
rect 38764 16037 38792 16068
rect 40696 16037 40724 16068
rect 40862 16056 40868 16068
rect 40920 16056 40926 16108
rect 43530 16096 43536 16108
rect 43491 16068 43536 16096
rect 43530 16056 43536 16068
rect 43588 16056 43594 16108
rect 37001 16031 37059 16037
rect 37001 16028 37013 16031
rect 36320 16000 37013 16028
rect 36320 15988 36326 16000
rect 37001 15997 37013 16000
rect 37047 15997 37059 16031
rect 37001 15991 37059 15997
rect 38749 16031 38807 16037
rect 38749 15997 38761 16031
rect 38795 15997 38807 16031
rect 38749 15991 38807 15997
rect 38841 16031 38899 16037
rect 38841 15997 38853 16031
rect 38887 15997 38899 16031
rect 38841 15991 38899 15997
rect 40681 16031 40739 16037
rect 40681 15997 40693 16031
rect 40727 15997 40739 16031
rect 40681 15991 40739 15997
rect 40957 16031 41015 16037
rect 40957 15997 40969 16031
rect 41003 16028 41015 16031
rect 41138 16028 41144 16040
rect 41003 16000 41144 16028
rect 41003 15997 41015 16000
rect 40957 15991 41015 15997
rect 26237 15963 26295 15969
rect 22603 15932 23796 15960
rect 25424 15932 26188 15960
rect 22603 15929 22615 15932
rect 22557 15923 22615 15929
rect 25424 15904 25452 15932
rect 25406 15892 25412 15904
rect 20594 15864 25412 15892
rect 25406 15852 25412 15864
rect 25464 15852 25470 15904
rect 26160 15892 26188 15932
rect 26237 15929 26249 15963
rect 26283 15960 26295 15963
rect 26786 15960 26792 15972
rect 26283 15932 26792 15960
rect 26283 15929 26295 15932
rect 26237 15923 26295 15929
rect 26786 15920 26792 15932
rect 26844 15960 26850 15972
rect 30190 15960 30196 15972
rect 26844 15932 30196 15960
rect 26844 15920 26850 15932
rect 30190 15920 30196 15932
rect 30248 15920 30254 15972
rect 37090 15960 37096 15972
rect 30300 15932 37096 15960
rect 28537 15895 28595 15901
rect 28537 15892 28549 15895
rect 26160 15864 28549 15892
rect 28537 15861 28549 15864
rect 28583 15892 28595 15895
rect 28902 15892 28908 15904
rect 28583 15864 28908 15892
rect 28583 15861 28595 15864
rect 28537 15855 28595 15861
rect 28902 15852 28908 15864
rect 28960 15892 28966 15904
rect 29086 15892 29092 15904
rect 28960 15864 29092 15892
rect 28960 15852 28966 15864
rect 29086 15852 29092 15864
rect 29144 15852 29150 15904
rect 29730 15852 29736 15904
rect 29788 15892 29794 15904
rect 30300 15892 30328 15932
rect 37090 15920 37096 15932
rect 37148 15920 37154 15972
rect 38378 15920 38384 15972
rect 38436 15960 38442 15972
rect 38856 15960 38884 15991
rect 38436 15932 38884 15960
rect 39025 15963 39083 15969
rect 38436 15920 38442 15932
rect 39025 15929 39037 15963
rect 39071 15960 39083 15963
rect 40696 15960 40724 15991
rect 41138 15988 41144 16000
rect 41196 15988 41202 16040
rect 43622 16028 43628 16040
rect 43583 16000 43628 16028
rect 43622 15988 43628 16000
rect 43680 15988 43686 16040
rect 43809 16031 43867 16037
rect 43809 15997 43821 16031
rect 43855 16028 43867 16031
rect 44361 16031 44419 16037
rect 44361 16028 44373 16031
rect 43855 16000 44373 16028
rect 43855 15997 43867 16000
rect 43809 15991 43867 15997
rect 44361 15997 44373 16000
rect 44407 15997 44419 16031
rect 44542 16028 44548 16040
rect 44503 16000 44548 16028
rect 44361 15991 44419 15997
rect 43824 15960 43852 15991
rect 44542 15988 44548 16000
rect 44600 15988 44606 16040
rect 39071 15932 40632 15960
rect 40696 15932 43852 15960
rect 44729 15963 44787 15969
rect 39071 15929 39083 15932
rect 39025 15923 39083 15929
rect 35894 15892 35900 15904
rect 29788 15864 30328 15892
rect 35855 15864 35900 15892
rect 29788 15852 29794 15864
rect 35894 15852 35900 15864
rect 35952 15852 35958 15904
rect 37277 15895 37335 15901
rect 37277 15861 37289 15895
rect 37323 15892 37335 15895
rect 39850 15892 39856 15904
rect 37323 15864 39856 15892
rect 37323 15861 37335 15864
rect 37277 15855 37335 15861
rect 39850 15852 39856 15864
rect 39908 15852 39914 15904
rect 40604 15892 40632 15932
rect 44729 15929 44741 15963
rect 44775 15960 44787 15963
rect 57974 15960 57980 15972
rect 44775 15932 57980 15960
rect 44775 15929 44787 15932
rect 44729 15923 44787 15929
rect 57974 15920 57980 15932
rect 58032 15920 58038 15972
rect 45830 15892 45836 15904
rect 40604 15864 45836 15892
rect 45830 15852 45836 15864
rect 45888 15852 45894 15904
rect 1104 15802 58880 15824
rect 1104 15750 20246 15802
rect 20298 15750 20310 15802
rect 20362 15750 20374 15802
rect 20426 15750 20438 15802
rect 20490 15750 39510 15802
rect 39562 15750 39574 15802
rect 39626 15750 39638 15802
rect 39690 15750 39702 15802
rect 39754 15750 58880 15802
rect 1104 15728 58880 15750
rect 1578 15688 1584 15700
rect 1539 15660 1584 15688
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 18874 15688 18880 15700
rect 17696 15660 18880 15688
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 17696 15561 17724 15660
rect 18874 15648 18880 15660
rect 18932 15688 18938 15700
rect 18932 15660 20622 15688
rect 18932 15648 18938 15660
rect 20594 15620 20622 15660
rect 21174 15648 21180 15700
rect 21232 15688 21238 15700
rect 22002 15688 22008 15700
rect 21232 15660 22008 15688
rect 21232 15648 21238 15660
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 28537 15691 28595 15697
rect 28537 15657 28549 15691
rect 28583 15688 28595 15691
rect 29270 15688 29276 15700
rect 28583 15660 29276 15688
rect 28583 15657 28595 15660
rect 28537 15651 28595 15657
rect 29270 15648 29276 15660
rect 29328 15648 29334 15700
rect 35986 15648 35992 15700
rect 36044 15688 36050 15700
rect 36081 15691 36139 15697
rect 36081 15688 36093 15691
rect 36044 15660 36093 15688
rect 36044 15648 36050 15660
rect 36081 15657 36093 15660
rect 36127 15657 36139 15691
rect 37090 15688 37096 15700
rect 37051 15660 37096 15688
rect 36081 15651 36139 15657
rect 37090 15648 37096 15660
rect 37148 15648 37154 15700
rect 37737 15691 37795 15697
rect 37737 15657 37749 15691
rect 37783 15688 37795 15691
rect 37826 15688 37832 15700
rect 37783 15660 37832 15688
rect 37783 15657 37795 15660
rect 37737 15651 37795 15657
rect 37826 15648 37832 15660
rect 37884 15648 37890 15700
rect 33689 15623 33747 15629
rect 33689 15620 33701 15623
rect 20594 15592 33701 15620
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15521 17739 15555
rect 17862 15552 17868 15564
rect 17823 15524 17868 15552
rect 17681 15515 17739 15521
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 18782 15552 18788 15564
rect 18743 15524 18788 15552
rect 18782 15512 18788 15524
rect 18840 15552 18846 15564
rect 18840 15524 21312 15552
rect 18840 15512 18846 15524
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 17589 15487 17647 15493
rect 17589 15484 17601 15487
rect 10376 15456 17601 15484
rect 10376 15444 10382 15456
rect 17589 15453 17601 15456
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 19978 15444 19984 15496
rect 20036 15484 20042 15496
rect 21174 15484 21180 15496
rect 20036 15456 21180 15484
rect 20036 15444 20042 15456
rect 21174 15444 21180 15456
rect 21232 15444 21238 15496
rect 21284 15484 21312 15524
rect 21358 15512 21364 15564
rect 21416 15552 21422 15564
rect 22097 15555 22155 15561
rect 22097 15552 22109 15555
rect 21416 15524 22109 15552
rect 21416 15512 21422 15524
rect 22097 15521 22109 15524
rect 22143 15521 22155 15555
rect 24394 15552 24400 15564
rect 22097 15515 22155 15521
rect 23676 15524 24400 15552
rect 23676 15496 23704 15524
rect 24394 15512 24400 15524
rect 24452 15552 24458 15564
rect 25225 15555 25283 15561
rect 25225 15552 25237 15555
rect 24452 15524 25237 15552
rect 24452 15512 24458 15524
rect 25225 15521 25237 15524
rect 25271 15521 25283 15555
rect 25225 15515 25283 15521
rect 28350 15512 28356 15564
rect 28408 15552 28414 15564
rect 33060 15561 33088 15592
rect 33689 15589 33701 15592
rect 33735 15620 33747 15623
rect 35894 15620 35900 15632
rect 33735 15592 35900 15620
rect 33735 15589 33747 15592
rect 33689 15583 33747 15589
rect 35894 15580 35900 15592
rect 35952 15580 35958 15632
rect 28445 15555 28503 15561
rect 28445 15552 28457 15555
rect 28408 15524 28457 15552
rect 28408 15512 28414 15524
rect 28445 15521 28457 15524
rect 28491 15552 28503 15555
rect 29089 15555 29147 15561
rect 29089 15552 29101 15555
rect 28491 15524 29101 15552
rect 28491 15521 28503 15524
rect 28445 15515 28503 15521
rect 29089 15521 29101 15524
rect 29135 15521 29147 15555
rect 32401 15555 32459 15561
rect 32401 15552 32413 15555
rect 29089 15515 29147 15521
rect 29610 15524 32413 15552
rect 23658 15484 23664 15496
rect 21284 15456 23664 15484
rect 23658 15444 23664 15456
rect 23716 15444 23722 15496
rect 25406 15484 25412 15496
rect 25367 15456 25412 15484
rect 25406 15444 25412 15456
rect 25464 15444 25470 15496
rect 25498 15444 25504 15496
rect 25556 15484 25562 15496
rect 29610 15484 29638 15524
rect 32401 15521 32413 15524
rect 32447 15552 32459 15555
rect 32953 15555 33011 15561
rect 32953 15552 32965 15555
rect 32447 15524 32965 15552
rect 32447 15521 32459 15524
rect 32401 15515 32459 15521
rect 32953 15521 32965 15524
rect 32999 15521 33011 15555
rect 32953 15515 33011 15521
rect 33045 15555 33103 15561
rect 33045 15521 33057 15555
rect 33091 15521 33103 15555
rect 37108 15552 37136 15648
rect 37645 15555 37703 15561
rect 37645 15552 37657 15555
rect 37108 15524 37657 15552
rect 33045 15515 33103 15521
rect 37645 15521 37657 15524
rect 37691 15521 37703 15555
rect 37844 15552 37872 15648
rect 38102 15580 38108 15632
rect 38160 15620 38166 15632
rect 38160 15592 38884 15620
rect 38160 15580 38166 15592
rect 38856 15561 38884 15592
rect 38565 15555 38623 15561
rect 38565 15552 38577 15555
rect 37844 15524 38577 15552
rect 37645 15515 37703 15521
rect 38565 15521 38577 15524
rect 38611 15521 38623 15555
rect 38565 15515 38623 15521
rect 38841 15555 38899 15561
rect 38841 15521 38853 15555
rect 38887 15521 38899 15555
rect 38841 15515 38899 15521
rect 25556 15456 29638 15484
rect 32968 15484 32996 15515
rect 39850 15512 39856 15564
rect 39908 15552 39914 15564
rect 40957 15555 41015 15561
rect 40957 15552 40969 15555
rect 39908 15524 40969 15552
rect 39908 15512 39914 15524
rect 40957 15521 40969 15524
rect 41003 15521 41015 15555
rect 40957 15515 41015 15521
rect 41509 15555 41567 15561
rect 41509 15521 41521 15555
rect 41555 15552 41567 15555
rect 44542 15552 44548 15564
rect 41555 15524 44548 15552
rect 41555 15521 41567 15524
rect 41509 15515 41567 15521
rect 44542 15512 44548 15524
rect 44600 15512 44606 15564
rect 33226 15484 33232 15496
rect 32968 15456 33088 15484
rect 33187 15456 33232 15484
rect 25556 15444 25562 15456
rect 33060 15416 33088 15456
rect 33226 15444 33232 15456
rect 33284 15444 33290 15496
rect 37274 15484 37280 15496
rect 33336 15456 37280 15484
rect 33336 15416 33364 15456
rect 37274 15444 37280 15456
rect 37332 15444 37338 15496
rect 38654 15484 38660 15496
rect 38615 15456 38660 15484
rect 38654 15444 38660 15456
rect 38712 15444 38718 15496
rect 41414 15484 41420 15496
rect 41375 15456 41420 15484
rect 41414 15444 41420 15456
rect 41472 15444 41478 15496
rect 33060 15388 33364 15416
rect 18966 15348 18972 15360
rect 18927 15320 18972 15348
rect 18966 15308 18972 15320
rect 19024 15308 19030 15360
rect 1104 15258 58880 15280
rect 1104 15206 10614 15258
rect 10666 15206 10678 15258
rect 10730 15206 10742 15258
rect 10794 15206 10806 15258
rect 10858 15206 29878 15258
rect 29930 15206 29942 15258
rect 29994 15206 30006 15258
rect 30058 15206 30070 15258
rect 30122 15206 49142 15258
rect 49194 15206 49206 15258
rect 49258 15206 49270 15258
rect 49322 15206 49334 15258
rect 49386 15206 58880 15258
rect 1104 15184 58880 15206
rect 1394 15144 1400 15156
rect 1355 15116 1400 15144
rect 1394 15104 1400 15116
rect 1452 15104 1458 15156
rect 18874 15144 18880 15156
rect 18835 15116 18880 15144
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 18138 15008 18144 15020
rect 18099 14980 18144 15008
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 17862 14940 17868 14952
rect 17823 14912 17868 14940
rect 17862 14900 17868 14912
rect 17920 14900 17926 14952
rect 18046 14940 18052 14952
rect 18007 14912 18052 14940
rect 18046 14900 18052 14912
rect 18104 14900 18110 14952
rect 36814 14940 36820 14952
rect 36775 14912 36820 14940
rect 36814 14900 36820 14912
rect 36872 14900 36878 14952
rect 37001 14943 37059 14949
rect 37001 14909 37013 14943
rect 37047 14940 37059 14943
rect 38102 14940 38108 14952
rect 37047 14912 38108 14940
rect 37047 14909 37059 14912
rect 37001 14903 37059 14909
rect 38102 14900 38108 14912
rect 38160 14900 38166 14952
rect 57425 14943 57483 14949
rect 57425 14909 57437 14943
rect 57471 14940 57483 14943
rect 58158 14940 58164 14952
rect 57471 14912 58164 14940
rect 57471 14909 57483 14912
rect 57425 14903 57483 14909
rect 58158 14900 58164 14912
rect 58216 14900 58222 14952
rect 35434 14832 35440 14884
rect 35492 14872 35498 14884
rect 36633 14875 36691 14881
rect 36633 14872 36645 14875
rect 35492 14844 36645 14872
rect 35492 14832 35498 14844
rect 36633 14841 36645 14844
rect 36679 14841 36691 14875
rect 36633 14835 36691 14841
rect 57974 14804 57980 14816
rect 57935 14776 57980 14804
rect 57974 14764 57980 14776
rect 58032 14764 58038 14816
rect 1104 14714 58880 14736
rect 1104 14662 20246 14714
rect 20298 14662 20310 14714
rect 20362 14662 20374 14714
rect 20426 14662 20438 14714
rect 20490 14662 39510 14714
rect 39562 14662 39574 14714
rect 39626 14662 39638 14714
rect 39690 14662 39702 14714
rect 39754 14662 58880 14714
rect 1104 14640 58880 14662
rect 57974 14600 57980 14612
rect 18432 14572 57980 14600
rect 1394 14464 1400 14476
rect 1355 14436 1400 14464
rect 1394 14424 1400 14436
rect 1452 14464 1458 14476
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1452 14436 2053 14464
rect 1452 14424 1458 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 14921 14467 14979 14473
rect 14921 14433 14933 14467
rect 14967 14464 14979 14467
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 14967 14436 15485 14464
rect 14967 14433 14979 14436
rect 14921 14427 14979 14433
rect 15473 14433 15485 14436
rect 15519 14464 15531 14467
rect 18432 14464 18460 14572
rect 57974 14560 57980 14572
rect 58032 14560 58038 14612
rect 23658 14532 23664 14544
rect 23619 14504 23664 14532
rect 23658 14492 23664 14504
rect 23716 14492 23722 14544
rect 52454 14532 52460 14544
rect 52415 14504 52460 14532
rect 52454 14492 52460 14504
rect 52512 14492 52518 14544
rect 54386 14532 54392 14544
rect 52932 14504 54392 14532
rect 15519 14436 18460 14464
rect 22465 14467 22523 14473
rect 15519 14433 15531 14436
rect 15473 14427 15531 14433
rect 22465 14433 22477 14467
rect 22511 14464 22523 14467
rect 22554 14464 22560 14476
rect 22511 14436 22560 14464
rect 22511 14433 22523 14436
rect 22465 14427 22523 14433
rect 22554 14424 22560 14436
rect 22612 14424 22618 14476
rect 36998 14424 37004 14476
rect 37056 14464 37062 14476
rect 52932 14473 52960 14504
rect 54386 14492 54392 14504
rect 54444 14492 54450 14544
rect 37093 14467 37151 14473
rect 37093 14464 37105 14467
rect 37056 14436 37105 14464
rect 37056 14424 37062 14436
rect 37093 14433 37105 14436
rect 37139 14433 37151 14467
rect 37093 14427 37151 14433
rect 51997 14467 52055 14473
rect 51997 14433 52009 14467
rect 52043 14464 52055 14467
rect 52917 14467 52975 14473
rect 52917 14464 52929 14467
rect 52043 14436 52929 14464
rect 52043 14433 52055 14436
rect 51997 14427 52055 14433
rect 52917 14433 52929 14436
rect 52963 14433 52975 14467
rect 53098 14464 53104 14476
rect 53059 14436 53104 14464
rect 52917 14427 52975 14433
rect 53098 14424 53104 14436
rect 53156 14424 53162 14476
rect 57517 14467 57575 14473
rect 57517 14433 57529 14467
rect 57563 14464 57575 14467
rect 58158 14464 58164 14476
rect 57563 14436 58164 14464
rect 57563 14433 57575 14436
rect 57517 14427 57575 14433
rect 58158 14424 58164 14436
rect 58216 14424 58222 14476
rect 53193 14399 53251 14405
rect 53193 14365 53205 14399
rect 53239 14365 53251 14399
rect 53193 14359 53251 14365
rect 1581 14331 1639 14337
rect 1581 14297 1593 14331
rect 1627 14328 1639 14331
rect 17678 14328 17684 14340
rect 1627 14300 17684 14328
rect 1627 14297 1639 14300
rect 1581 14291 1639 14297
rect 17678 14288 17684 14300
rect 17736 14288 17742 14340
rect 18046 14288 18052 14340
rect 18104 14328 18110 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 18104 14300 22569 14328
rect 18104 14288 18110 14300
rect 22557 14297 22569 14300
rect 22603 14328 22615 14331
rect 23198 14328 23204 14340
rect 22603 14300 23204 14328
rect 22603 14297 22615 14300
rect 22557 14291 22615 14297
rect 23198 14288 23204 14300
rect 23256 14288 23262 14340
rect 36814 14288 36820 14340
rect 36872 14328 36878 14340
rect 37001 14331 37059 14337
rect 37001 14328 37013 14331
rect 36872 14300 37013 14328
rect 36872 14288 36878 14300
rect 37001 14297 37013 14300
rect 37047 14297 37059 14331
rect 53208 14328 53236 14359
rect 57977 14331 58035 14337
rect 57977 14328 57989 14331
rect 53208 14300 57989 14328
rect 37001 14291 37059 14297
rect 57977 14297 57989 14300
rect 58023 14297 58035 14331
rect 57977 14291 58035 14297
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 14829 14263 14887 14269
rect 14829 14260 14841 14263
rect 13780 14232 14841 14260
rect 13780 14220 13786 14232
rect 14829 14229 14841 14232
rect 14875 14229 14887 14263
rect 23566 14260 23572 14272
rect 23527 14232 23572 14260
rect 14829 14223 14887 14229
rect 23566 14220 23572 14232
rect 23624 14220 23630 14272
rect 54386 14220 54392 14272
rect 54444 14260 54450 14272
rect 56318 14260 56324 14272
rect 54444 14232 56324 14260
rect 54444 14220 54450 14232
rect 56318 14220 56324 14232
rect 56376 14220 56382 14272
rect 1104 14170 58880 14192
rect 1104 14118 10614 14170
rect 10666 14118 10678 14170
rect 10730 14118 10742 14170
rect 10794 14118 10806 14170
rect 10858 14118 29878 14170
rect 29930 14118 29942 14170
rect 29994 14118 30006 14170
rect 30058 14118 30070 14170
rect 30122 14118 49142 14170
rect 49194 14118 49206 14170
rect 49258 14118 49270 14170
rect 49322 14118 49334 14170
rect 49386 14118 58880 14170
rect 1104 14096 58880 14118
rect 13556 13892 14412 13920
rect 1394 13852 1400 13864
rect 1355 13824 1400 13852
rect 1394 13812 1400 13824
rect 1452 13852 1458 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1452 13824 2053 13852
rect 1452 13812 1458 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 10594 13852 10600 13864
rect 10555 13824 10600 13852
rect 2041 13815 2099 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 13556 13861 13584 13892
rect 10781 13855 10839 13861
rect 10781 13821 10793 13855
rect 10827 13852 10839 13855
rect 11793 13855 11851 13861
rect 11793 13852 11805 13855
rect 10827 13824 11805 13852
rect 10827 13821 10839 13824
rect 10781 13815 10839 13821
rect 11793 13821 11805 13824
rect 11839 13852 11851 13855
rect 13541 13855 13599 13861
rect 13541 13852 13553 13855
rect 11839 13824 13553 13852
rect 11839 13821 11851 13824
rect 11793 13815 11851 13821
rect 13541 13821 13553 13824
rect 13587 13821 13599 13855
rect 13722 13852 13728 13864
rect 13683 13824 13728 13852
rect 13541 13815 13599 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14384 13861 14412 13892
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13852 14427 13855
rect 21082 13852 21088 13864
rect 14415 13824 21088 13852
rect 14415 13821 14427 13824
rect 14369 13815 14427 13821
rect 21082 13812 21088 13824
rect 21140 13812 21146 13864
rect 22830 13852 22836 13864
rect 22791 13824 22836 13852
rect 22830 13812 22836 13824
rect 22888 13812 22894 13864
rect 23017 13855 23075 13861
rect 23017 13821 23029 13855
rect 23063 13852 23075 13855
rect 23566 13852 23572 13864
rect 23063 13824 23572 13852
rect 23063 13821 23075 13824
rect 23017 13815 23075 13821
rect 23566 13812 23572 13824
rect 23624 13812 23630 13864
rect 34698 13812 34704 13864
rect 34756 13852 34762 13864
rect 35345 13855 35403 13861
rect 35345 13852 35357 13855
rect 34756 13824 35357 13852
rect 34756 13812 34762 13824
rect 35345 13821 35357 13824
rect 35391 13821 35403 13855
rect 35345 13815 35403 13821
rect 35621 13855 35679 13861
rect 35621 13821 35633 13855
rect 35667 13821 35679 13855
rect 35621 13815 35679 13821
rect 2130 13744 2136 13796
rect 2188 13784 2194 13796
rect 10413 13787 10471 13793
rect 10413 13784 10425 13787
rect 2188 13756 10425 13784
rect 2188 13744 2194 13756
rect 10413 13753 10425 13756
rect 10459 13753 10471 13787
rect 13814 13784 13820 13796
rect 13775 13756 13820 13784
rect 10413 13747 10471 13753
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 19886 13744 19892 13796
rect 19944 13784 19950 13796
rect 22649 13787 22707 13793
rect 22649 13784 22661 13787
rect 19944 13756 22661 13784
rect 19944 13744 19950 13756
rect 22649 13753 22661 13756
rect 22695 13753 22707 13787
rect 22649 13747 22707 13753
rect 1581 13719 1639 13725
rect 1581 13685 1593 13719
rect 1627 13716 1639 13719
rect 2406 13716 2412 13728
rect 1627 13688 2412 13716
rect 1627 13685 1639 13688
rect 1581 13679 1639 13685
rect 2406 13676 2412 13688
rect 2464 13676 2470 13728
rect 23566 13716 23572 13728
rect 23479 13688 23572 13716
rect 23566 13676 23572 13688
rect 23624 13716 23630 13728
rect 34606 13716 34612 13728
rect 23624 13688 34612 13716
rect 23624 13676 23630 13688
rect 34606 13676 34612 13688
rect 34664 13716 34670 13728
rect 35636 13716 35664 13815
rect 34664 13688 35664 13716
rect 35805 13719 35863 13725
rect 34664 13676 34670 13688
rect 35805 13685 35817 13719
rect 35851 13716 35863 13719
rect 55122 13716 55128 13728
rect 35851 13688 55128 13716
rect 35851 13685 35863 13688
rect 35805 13679 35863 13685
rect 55122 13676 55128 13688
rect 55180 13676 55186 13728
rect 1104 13626 58880 13648
rect 1104 13574 20246 13626
rect 20298 13574 20310 13626
rect 20362 13574 20374 13626
rect 20426 13574 20438 13626
rect 20490 13574 39510 13626
rect 39562 13574 39574 13626
rect 39626 13574 39638 13626
rect 39690 13574 39702 13626
rect 39754 13574 58880 13626
rect 1104 13552 58880 13574
rect 2406 13512 2412 13524
rect 2367 13484 2412 13512
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 15562 13512 15568 13524
rect 10244 13484 15568 13512
rect 1489 13447 1547 13453
rect 1489 13413 1501 13447
rect 1535 13444 1547 13447
rect 1578 13444 1584 13456
rect 1535 13416 1584 13444
rect 1535 13413 1547 13416
rect 1489 13407 1547 13413
rect 1578 13404 1584 13416
rect 1636 13444 1642 13456
rect 2498 13444 2504 13456
rect 1636 13416 2504 13444
rect 1636 13404 1642 13416
rect 2498 13404 2504 13416
rect 2556 13404 2562 13456
rect 2317 13379 2375 13385
rect 2317 13345 2329 13379
rect 2363 13345 2375 13379
rect 2317 13339 2375 13345
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 1949 13175 2007 13181
rect 1949 13172 1961 13175
rect 1728 13144 1961 13172
rect 1728 13132 1734 13144
rect 1949 13141 1961 13144
rect 1995 13141 2007 13175
rect 2332 13172 2360 13339
rect 2498 13308 2504 13320
rect 2459 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13268 2562 13320
rect 10244 13308 10272 13484
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 10594 13444 10600 13456
rect 10336 13416 10600 13444
rect 10336 13385 10364 13416
rect 10594 13404 10600 13416
rect 10652 13444 10658 13456
rect 11241 13447 11299 13453
rect 11241 13444 11253 13447
rect 10652 13416 11253 13444
rect 10652 13404 10658 13416
rect 11241 13413 11253 13416
rect 11287 13413 11299 13447
rect 13722 13444 13728 13456
rect 11241 13407 11299 13413
rect 12820 13416 13728 13444
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13345 10379 13379
rect 10502 13376 10508 13388
rect 10415 13348 10508 13376
rect 10321 13339 10379 13345
rect 10502 13336 10508 13348
rect 10560 13376 10566 13388
rect 11333 13379 11391 13385
rect 10560 13348 11008 13376
rect 10560 13336 10566 13348
rect 10244 13280 10364 13308
rect 2406 13200 2412 13252
rect 2464 13240 2470 13252
rect 10229 13243 10287 13249
rect 10229 13240 10241 13243
rect 2464 13212 10241 13240
rect 2464 13200 2470 13212
rect 10229 13209 10241 13212
rect 10275 13209 10287 13243
rect 10229 13203 10287 13209
rect 3237 13175 3295 13181
rect 3237 13172 3249 13175
rect 2332 13144 3249 13172
rect 1949 13135 2007 13141
rect 3237 13141 3249 13144
rect 3283 13172 3295 13175
rect 10336 13172 10364 13280
rect 10980 13240 11008 13348
rect 11333 13345 11345 13379
rect 11379 13376 11391 13379
rect 11882 13376 11888 13388
rect 11379 13348 11888 13376
rect 11379 13345 11391 13348
rect 11333 13339 11391 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12820 13385 12848 13416
rect 13722 13404 13728 13416
rect 13780 13404 13786 13456
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 12989 13379 13047 13385
rect 12989 13345 13001 13379
rect 13035 13376 13047 13379
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13035 13348 13553 13376
rect 13035 13345 13047 13348
rect 12989 13339 13047 13345
rect 13541 13345 13553 13348
rect 13587 13376 13599 13379
rect 18966 13376 18972 13388
rect 13587 13348 18972 13376
rect 13587 13345 13599 13348
rect 13541 13339 13599 13345
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 11112 13280 12633 13308
rect 11112 13268 11118 13280
rect 12621 13277 12633 13280
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 13004 13240 13032 13339
rect 18966 13336 18972 13348
rect 19024 13336 19030 13388
rect 10980 13212 13032 13240
rect 11882 13172 11888 13184
rect 3283 13144 10364 13172
rect 11843 13144 11888 13172
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 1104 13082 58880 13104
rect 1104 13030 10614 13082
rect 10666 13030 10678 13082
rect 10730 13030 10742 13082
rect 10794 13030 10806 13082
rect 10858 13030 29878 13082
rect 29930 13030 29942 13082
rect 29994 13030 30006 13082
rect 30058 13030 30070 13082
rect 30122 13030 49142 13082
rect 49194 13030 49206 13082
rect 49258 13030 49270 13082
rect 49322 13030 49334 13082
rect 49386 13030 58880 13082
rect 1104 13008 58880 13030
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 10597 12971 10655 12977
rect 10597 12968 10609 12971
rect 10560 12940 10609 12968
rect 10560 12928 10566 12940
rect 10597 12937 10609 12940
rect 10643 12937 10655 12971
rect 10597 12931 10655 12937
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 57425 12835 57483 12841
rect 57425 12801 57437 12835
rect 57471 12832 57483 12835
rect 57882 12832 57888 12844
rect 57471 12804 57888 12832
rect 57471 12801 57483 12804
rect 57425 12795 57483 12801
rect 57882 12792 57888 12804
rect 57940 12832 57946 12844
rect 57940 12804 58112 12832
rect 57940 12792 57946 12804
rect 58084 12773 58112 12804
rect 58069 12767 58127 12773
rect 58069 12733 58081 12767
rect 58115 12733 58127 12767
rect 58069 12727 58127 12733
rect 1581 12699 1639 12705
rect 1581 12665 1593 12699
rect 1627 12665 1639 12699
rect 57885 12699 57943 12705
rect 57885 12696 57897 12699
rect 1581 12659 1639 12665
rect 42490 12668 57897 12696
rect 1596 12628 1624 12659
rect 1854 12628 1860 12640
rect 1596 12600 1860 12628
rect 1854 12588 1860 12600
rect 1912 12628 1918 12640
rect 2133 12631 2191 12637
rect 2133 12628 2145 12631
rect 1912 12600 2145 12628
rect 1912 12588 1918 12600
rect 2133 12597 2145 12600
rect 2179 12597 2191 12631
rect 2133 12591 2191 12597
rect 38930 12588 38936 12640
rect 38988 12628 38994 12640
rect 42490 12628 42518 12668
rect 57885 12665 57897 12668
rect 57931 12665 57943 12699
rect 57885 12659 57943 12665
rect 38988 12600 42518 12628
rect 38988 12588 38994 12600
rect 1104 12538 58880 12560
rect 1104 12486 20246 12538
rect 20298 12486 20310 12538
rect 20362 12486 20374 12538
rect 20426 12486 20438 12538
rect 20490 12486 39510 12538
rect 39562 12486 39574 12538
rect 39626 12486 39638 12538
rect 39690 12486 39702 12538
rect 39754 12486 58880 12538
rect 1104 12464 58880 12486
rect 57425 12291 57483 12297
rect 57425 12257 57437 12291
rect 57471 12288 57483 12291
rect 58158 12288 58164 12300
rect 57471 12260 58164 12288
rect 57471 12257 57483 12260
rect 57425 12251 57483 12257
rect 58158 12248 58164 12260
rect 58216 12248 58222 12300
rect 2222 12180 2228 12232
rect 2280 12220 2286 12232
rect 36170 12220 36176 12232
rect 2280 12192 36176 12220
rect 2280 12180 2286 12192
rect 36170 12180 36176 12192
rect 36228 12180 36234 12232
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 57977 12155 58035 12161
rect 57977 12152 57989 12155
rect 11940 12124 57989 12152
rect 11940 12112 11946 12124
rect 57977 12121 57989 12124
rect 58023 12121 58035 12155
rect 57977 12115 58035 12121
rect 1104 11994 58880 12016
rect 1104 11942 10614 11994
rect 10666 11942 10678 11994
rect 10730 11942 10742 11994
rect 10794 11942 10806 11994
rect 10858 11942 29878 11994
rect 29930 11942 29942 11994
rect 29994 11942 30006 11994
rect 30058 11942 30070 11994
rect 30122 11942 49142 11994
rect 49194 11942 49206 11994
rect 49258 11942 49270 11994
rect 49322 11942 49334 11994
rect 49386 11942 58880 11994
rect 1104 11920 58880 11942
rect 1394 11608 1400 11620
rect 1355 11580 1400 11608
rect 1394 11568 1400 11580
rect 1452 11568 1458 11620
rect 1581 11611 1639 11617
rect 1581 11577 1593 11611
rect 1627 11608 1639 11611
rect 2222 11608 2228 11620
rect 1627 11580 2228 11608
rect 1627 11577 1639 11580
rect 1581 11571 1639 11577
rect 2222 11568 2228 11580
rect 2280 11568 2286 11620
rect 57882 11568 57888 11620
rect 57940 11608 57946 11620
rect 57977 11611 58035 11617
rect 57977 11608 57989 11611
rect 57940 11580 57989 11608
rect 57940 11568 57946 11580
rect 57977 11577 57989 11580
rect 58023 11577 58035 11611
rect 58158 11608 58164 11620
rect 58119 11580 58164 11608
rect 57977 11571 58035 11577
rect 58158 11568 58164 11580
rect 58216 11568 58222 11620
rect 1104 11450 58880 11472
rect 1104 11398 20246 11450
rect 20298 11398 20310 11450
rect 20362 11398 20374 11450
rect 20426 11398 20438 11450
rect 20490 11398 39510 11450
rect 39562 11398 39574 11450
rect 39626 11398 39638 11450
rect 39690 11398 39702 11450
rect 39754 11398 58880 11450
rect 1104 11376 58880 11398
rect 57882 11336 57888 11348
rect 57843 11308 57888 11336
rect 57882 11296 57888 11308
rect 57940 11296 57946 11348
rect 57517 11271 57575 11277
rect 57517 11237 57529 11271
rect 57563 11268 57575 11271
rect 58250 11268 58256 11280
rect 57563 11240 58256 11268
rect 57563 11237 57575 11240
rect 57517 11231 57575 11237
rect 58250 11228 58256 11240
rect 58308 11228 58314 11280
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11200 1639 11203
rect 2225 11203 2283 11209
rect 2225 11200 2237 11203
rect 1627 11172 2237 11200
rect 1627 11169 1639 11172
rect 1581 11163 1639 11169
rect 2225 11169 2237 11172
rect 2271 11200 2283 11203
rect 41414 11200 41420 11212
rect 2271 11172 41420 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 41414 11160 41420 11172
rect 41472 11160 41478 11212
rect 56410 11092 56416 11144
rect 56468 11132 56474 11144
rect 57241 11135 57299 11141
rect 57241 11132 57253 11135
rect 56468 11104 57253 11132
rect 56468 11092 56474 11104
rect 57241 11101 57253 11104
rect 57287 11101 57299 11135
rect 57241 11095 57299 11101
rect 57425 11135 57483 11141
rect 57425 11101 57437 11135
rect 57471 11101 57483 11135
rect 57425 11095 57483 11101
rect 1486 10996 1492 11008
rect 1447 10968 1492 10996
rect 1486 10956 1492 10968
rect 1544 10956 1550 11008
rect 28534 10956 28540 11008
rect 28592 10996 28598 11008
rect 56689 10999 56747 11005
rect 56689 10996 56701 10999
rect 28592 10968 56701 10996
rect 28592 10956 28598 10968
rect 56689 10965 56701 10968
rect 56735 10996 56747 10999
rect 57440 10996 57468 11095
rect 56735 10968 57468 10996
rect 56735 10965 56747 10968
rect 56689 10959 56747 10965
rect 1104 10906 58880 10928
rect 1104 10854 10614 10906
rect 10666 10854 10678 10906
rect 10730 10854 10742 10906
rect 10794 10854 10806 10906
rect 10858 10854 29878 10906
rect 29930 10854 29942 10906
rect 29994 10854 30006 10906
rect 30058 10854 30070 10906
rect 30122 10854 49142 10906
rect 49194 10854 49206 10906
rect 49258 10854 49270 10906
rect 49322 10854 49334 10906
rect 49386 10854 58880 10906
rect 1104 10832 58880 10854
rect 23290 10752 23296 10804
rect 23348 10792 23354 10804
rect 23845 10795 23903 10801
rect 23845 10792 23857 10795
rect 23348 10764 23857 10792
rect 23348 10752 23354 10764
rect 23845 10761 23857 10764
rect 23891 10792 23903 10795
rect 23891 10764 24808 10792
rect 23891 10761 23903 10764
rect 23845 10755 23903 10761
rect 24780 10597 24808 10764
rect 24581 10591 24639 10597
rect 24581 10557 24593 10591
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 24765 10591 24823 10597
rect 24765 10557 24777 10591
rect 24811 10588 24823 10591
rect 30926 10588 30932 10600
rect 24811 10560 30932 10588
rect 24811 10557 24823 10560
rect 24765 10551 24823 10557
rect 24397 10523 24455 10529
rect 24397 10520 24409 10523
rect 6426 10492 24409 10520
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 6426 10452 6454 10492
rect 24397 10489 24409 10492
rect 24443 10489 24455 10523
rect 24596 10520 24624 10551
rect 30926 10548 30932 10560
rect 30984 10548 30990 10600
rect 25038 10520 25044 10532
rect 24596 10492 25044 10520
rect 24397 10483 24455 10489
rect 25038 10480 25044 10492
rect 25096 10480 25102 10532
rect 2280 10424 6454 10452
rect 2280 10412 2286 10424
rect 56410 10412 56416 10464
rect 56468 10452 56474 10464
rect 56781 10455 56839 10461
rect 56781 10452 56793 10455
rect 56468 10424 56793 10452
rect 56468 10412 56474 10424
rect 56781 10421 56793 10424
rect 56827 10421 56839 10455
rect 56781 10415 56839 10421
rect 1104 10362 58880 10384
rect 1104 10310 20246 10362
rect 20298 10310 20310 10362
rect 20362 10310 20374 10362
rect 20426 10310 20438 10362
rect 20490 10310 39510 10362
rect 39562 10310 39574 10362
rect 39626 10310 39638 10362
rect 39690 10310 39702 10362
rect 39754 10310 58880 10362
rect 1104 10288 58880 10310
rect 57425 10183 57483 10189
rect 57425 10149 57437 10183
rect 57471 10180 57483 10183
rect 57790 10180 57796 10192
rect 57471 10152 57796 10180
rect 57471 10149 57483 10152
rect 57425 10143 57483 10149
rect 57790 10140 57796 10152
rect 57848 10180 57854 10192
rect 57977 10183 58035 10189
rect 57977 10180 57989 10183
rect 57848 10152 57989 10180
rect 57848 10140 57854 10152
rect 57977 10149 57989 10152
rect 58023 10149 58035 10183
rect 58158 10180 58164 10192
rect 58119 10152 58164 10180
rect 57977 10143 58035 10149
rect 58158 10140 58164 10152
rect 58216 10140 58222 10192
rect 1486 9908 1492 9920
rect 1447 9880 1492 9908
rect 1486 9868 1492 9880
rect 1544 9868 1550 9920
rect 33318 9868 33324 9920
rect 33376 9908 33382 9920
rect 42334 9908 42340 9920
rect 33376 9880 42340 9908
rect 33376 9868 33382 9880
rect 42334 9868 42340 9880
rect 42392 9868 42398 9920
rect 1104 9818 58880 9840
rect 1104 9766 10614 9818
rect 10666 9766 10678 9818
rect 10730 9766 10742 9818
rect 10794 9766 10806 9818
rect 10858 9766 29878 9818
rect 29930 9766 29942 9818
rect 29994 9766 30006 9818
rect 30058 9766 30070 9818
rect 30122 9766 49142 9818
rect 49194 9766 49206 9818
rect 49258 9766 49270 9818
rect 49322 9766 49334 9818
rect 49386 9766 58880 9818
rect 1104 9744 58880 9766
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 49970 9704 49976 9716
rect 19116 9676 49976 9704
rect 19116 9664 19122 9676
rect 49970 9664 49976 9676
rect 50028 9664 50034 9716
rect 30926 9596 30932 9648
rect 30984 9636 30990 9648
rect 34609 9639 34667 9645
rect 34609 9636 34621 9639
rect 30984 9608 34621 9636
rect 30984 9596 30990 9608
rect 34609 9605 34621 9608
rect 34655 9605 34667 9639
rect 34609 9599 34667 9605
rect 1486 9500 1492 9512
rect 1447 9472 1492 9500
rect 1486 9460 1492 9472
rect 1544 9460 1550 9512
rect 34624 9500 34652 9599
rect 58158 9568 58164 9580
rect 58119 9540 58164 9568
rect 58158 9528 58164 9540
rect 58216 9528 58222 9580
rect 35161 9503 35219 9509
rect 35161 9500 35173 9503
rect 34624 9472 35173 9500
rect 35161 9469 35173 9472
rect 35207 9469 35219 9503
rect 35342 9500 35348 9512
rect 35303 9472 35348 9500
rect 35161 9463 35219 9469
rect 35342 9460 35348 9472
rect 35400 9460 35406 9512
rect 57977 9435 58035 9441
rect 57977 9432 57989 9435
rect 57348 9404 57989 9432
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 21818 9364 21824 9376
rect 1627 9336 21824 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 21818 9324 21824 9336
rect 21876 9324 21882 9376
rect 57348 9373 57376 9404
rect 57977 9401 57989 9404
rect 58023 9401 58035 9435
rect 57977 9395 58035 9401
rect 35437 9367 35495 9373
rect 35437 9333 35449 9367
rect 35483 9364 35495 9367
rect 57333 9367 57391 9373
rect 57333 9364 57345 9367
rect 35483 9336 57345 9364
rect 35483 9333 35495 9336
rect 35437 9327 35495 9333
rect 57333 9333 57345 9336
rect 57379 9333 57391 9367
rect 57333 9327 57391 9333
rect 1104 9274 58880 9296
rect 1104 9222 20246 9274
rect 20298 9222 20310 9274
rect 20362 9222 20374 9274
rect 20426 9222 20438 9274
rect 20490 9222 39510 9274
rect 39562 9222 39574 9274
rect 39626 9222 39638 9274
rect 39690 9222 39702 9274
rect 39754 9222 58880 9274
rect 1104 9200 58880 9222
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 9214 9092 9220 9104
rect 1627 9064 9220 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 9214 9052 9220 9064
rect 9272 9052 9278 9104
rect 1394 8888 1400 8900
rect 1355 8860 1400 8888
rect 1394 8848 1400 8860
rect 1452 8848 1458 8900
rect 1104 8730 58880 8752
rect 1104 8678 10614 8730
rect 10666 8678 10678 8730
rect 10730 8678 10742 8730
rect 10794 8678 10806 8730
rect 10858 8678 29878 8730
rect 29930 8678 29942 8730
rect 29994 8678 30006 8730
rect 30058 8678 30070 8730
rect 30122 8678 49142 8730
rect 49194 8678 49206 8730
rect 49258 8678 49270 8730
rect 49322 8678 49334 8730
rect 49386 8678 58880 8730
rect 1104 8656 58880 8678
rect 9214 8616 9220 8628
rect 9175 8588 9220 8616
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 9640 8588 10517 8616
rect 9640 8576 9646 8588
rect 10505 8585 10517 8588
rect 10551 8616 10563 8619
rect 26510 8616 26516 8628
rect 10551 8588 18046 8616
rect 26471 8588 26516 8616
rect 10551 8585 10563 8588
rect 10505 8579 10563 8585
rect 6426 8520 13860 8548
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2225 8347 2283 8353
rect 2225 8344 2237 8347
rect 1627 8316 2237 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 2225 8313 2237 8316
rect 2271 8344 2283 8347
rect 6426 8344 6454 8520
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 2271 8316 6454 8344
rect 8680 8452 8769 8480
rect 2271 8313 2283 8316
rect 2225 8307 2283 8313
rect 1486 8276 1492 8288
rect 1447 8248 1492 8276
rect 1486 8236 1492 8248
rect 1544 8236 1550 8288
rect 2498 8236 2504 8288
rect 2556 8276 2562 8288
rect 8680 8276 8708 8452
rect 8757 8449 8769 8452
rect 8803 8480 8815 8483
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 8803 8452 9873 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 9861 8449 9873 8452
rect 9907 8480 9919 8483
rect 13722 8480 13728 8492
rect 9907 8452 13728 8480
rect 9907 8449 9919 8452
rect 9861 8443 9919 8449
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 9582 8412 9588 8424
rect 9543 8384 9588 8412
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 13832 8344 13860 8520
rect 18018 8480 18046 8588
rect 26510 8576 26516 8588
rect 26568 8576 26574 8628
rect 18018 8452 20622 8480
rect 20594 8412 20622 8452
rect 41782 8412 41788 8424
rect 20594 8384 41788 8412
rect 41782 8372 41788 8384
rect 41840 8372 41846 8424
rect 25590 8344 25596 8356
rect 13832 8316 25596 8344
rect 25590 8304 25596 8316
rect 25648 8304 25654 8356
rect 38654 8304 38660 8356
rect 38712 8344 38718 8356
rect 57333 8347 57391 8353
rect 57333 8344 57345 8347
rect 38712 8316 57345 8344
rect 38712 8304 38718 8316
rect 57333 8313 57345 8316
rect 57379 8344 57391 8347
rect 57977 8347 58035 8353
rect 57977 8344 57989 8347
rect 57379 8316 57989 8344
rect 57379 8313 57391 8316
rect 57333 8307 57391 8313
rect 57977 8313 57989 8316
rect 58023 8313 58035 8347
rect 58158 8344 58164 8356
rect 58119 8316 58164 8344
rect 57977 8307 58035 8313
rect 58158 8304 58164 8316
rect 58216 8304 58222 8356
rect 2556 8248 8708 8276
rect 2556 8236 2562 8248
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 9732 8248 9777 8276
rect 9732 8236 9738 8248
rect 1104 8186 58880 8208
rect 1104 8134 20246 8186
rect 20298 8134 20310 8186
rect 20362 8134 20374 8186
rect 20426 8134 20438 8186
rect 20490 8134 39510 8186
rect 39562 8134 39574 8186
rect 39626 8134 39638 8186
rect 39690 8134 39702 8186
rect 39754 8134 58880 8186
rect 1104 8112 58880 8134
rect 25590 8032 25596 8084
rect 25648 8072 25654 8084
rect 25777 8075 25835 8081
rect 25777 8072 25789 8075
rect 25648 8044 25789 8072
rect 25648 8032 25654 8044
rect 25777 8041 25789 8044
rect 25823 8041 25835 8075
rect 25777 8035 25835 8041
rect 27890 8004 27896 8016
rect 26896 7976 27896 8004
rect 25774 7936 25780 7948
rect 25735 7908 25780 7936
rect 25774 7896 25780 7908
rect 25832 7896 25838 7948
rect 26053 7939 26111 7945
rect 26053 7905 26065 7939
rect 26099 7936 26111 7939
rect 26510 7936 26516 7948
rect 26099 7908 26516 7936
rect 26099 7905 26111 7908
rect 26053 7899 26111 7905
rect 26510 7896 26516 7908
rect 26568 7936 26574 7948
rect 26896 7945 26924 7976
rect 27890 7964 27896 7976
rect 27948 7964 27954 8016
rect 26881 7939 26939 7945
rect 26568 7908 26832 7936
rect 26568 7896 26574 7908
rect 20622 7828 20628 7880
rect 20680 7868 20686 7880
rect 26697 7871 26755 7877
rect 26697 7868 26709 7871
rect 20680 7840 26709 7868
rect 20680 7828 20686 7840
rect 26697 7837 26709 7840
rect 26743 7837 26755 7871
rect 26804 7868 26832 7908
rect 26881 7905 26893 7939
rect 26927 7905 26939 7939
rect 26881 7899 26939 7905
rect 26973 7939 27031 7945
rect 26973 7905 26985 7939
rect 27019 7905 27031 7939
rect 26973 7899 27031 7905
rect 26988 7868 27016 7899
rect 26804 7840 27016 7868
rect 26697 7831 26755 7837
rect 1104 7642 58880 7664
rect 1104 7590 10614 7642
rect 10666 7590 10678 7642
rect 10730 7590 10742 7642
rect 10794 7590 10806 7642
rect 10858 7590 29878 7642
rect 29930 7590 29942 7642
rect 29994 7590 30006 7642
rect 30058 7590 30070 7642
rect 30122 7590 49142 7642
rect 49194 7590 49206 7642
rect 49258 7590 49270 7642
rect 49322 7590 49334 7642
rect 49386 7590 58880 7642
rect 1104 7568 58880 7590
rect 26237 7531 26295 7537
rect 26237 7497 26249 7531
rect 26283 7528 26295 7531
rect 26510 7528 26516 7540
rect 26283 7500 26516 7528
rect 26283 7497 26295 7500
rect 26237 7491 26295 7497
rect 26510 7488 26516 7500
rect 26568 7488 26574 7540
rect 27890 7488 27896 7540
rect 27948 7528 27954 7540
rect 28077 7531 28135 7537
rect 28077 7528 28089 7531
rect 27948 7500 28089 7528
rect 27948 7488 27954 7500
rect 28077 7497 28089 7500
rect 28123 7497 28135 7531
rect 28077 7491 28135 7497
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7324 1458 7336
rect 2041 7327 2099 7333
rect 2041 7324 2053 7327
rect 1452 7296 2053 7324
rect 1452 7284 1458 7296
rect 2041 7293 2053 7296
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 28169 7327 28227 7333
rect 28169 7293 28181 7327
rect 28215 7293 28227 7327
rect 28169 7287 28227 7293
rect 57517 7327 57575 7333
rect 57517 7293 57529 7327
rect 57563 7324 57575 7327
rect 58158 7324 58164 7336
rect 57563 7296 58164 7324
rect 57563 7293 57575 7296
rect 57517 7287 57575 7293
rect 28184 7256 28212 7287
rect 58158 7284 58164 7296
rect 58216 7284 58222 7336
rect 28721 7259 28779 7265
rect 28721 7256 28733 7259
rect 28184 7228 28733 7256
rect 28721 7225 28733 7228
rect 28767 7256 28779 7259
rect 57882 7256 57888 7268
rect 28767 7228 57888 7256
rect 28767 7225 28779 7228
rect 28721 7219 28779 7225
rect 57882 7216 57888 7228
rect 57940 7216 57946 7268
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 57974 7188 57980 7200
rect 57935 7160 57980 7188
rect 57974 7148 57980 7160
rect 58032 7148 58038 7200
rect 1104 7098 58880 7120
rect 1104 7046 20246 7098
rect 20298 7046 20310 7098
rect 20362 7046 20374 7098
rect 20426 7046 20438 7098
rect 20490 7046 39510 7098
rect 39562 7046 39574 7098
rect 39626 7046 39638 7098
rect 39690 7046 39702 7098
rect 39754 7046 58880 7098
rect 1104 7024 58880 7046
rect 1486 6984 1492 6996
rect 1447 6956 1492 6984
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 1636 6956 2421 6984
rect 1636 6944 1642 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 1504 6916 1532 6944
rect 2498 6916 2504 6928
rect 1504 6888 2504 6916
rect 1688 6792 1716 6888
rect 2498 6876 2504 6888
rect 2556 6876 2562 6928
rect 57882 6916 57888 6928
rect 57843 6888 57888 6916
rect 57882 6876 57888 6888
rect 57940 6876 57946 6928
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 1670 6740 1676 6792
rect 1728 6740 1734 6792
rect 2332 6712 2360 6811
rect 2516 6789 2544 6876
rect 54113 6851 54171 6857
rect 54113 6817 54125 6851
rect 54159 6848 54171 6851
rect 57974 6848 57980 6860
rect 54159 6820 57980 6848
rect 54159 6817 54171 6820
rect 54113 6811 54171 6817
rect 57974 6808 57980 6820
rect 58032 6808 58038 6860
rect 58066 6808 58072 6860
rect 58124 6848 58130 6860
rect 58124 6820 58169 6848
rect 58124 6808 58130 6820
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6749 2559 6783
rect 2501 6743 2559 6749
rect 57425 6783 57483 6789
rect 57425 6749 57437 6783
rect 57471 6780 57483 6783
rect 58084 6780 58112 6808
rect 57471 6752 58112 6780
rect 57471 6749 57483 6752
rect 57425 6743 57483 6749
rect 3237 6715 3295 6721
rect 3237 6712 3249 6715
rect 2332 6684 3249 6712
rect 3237 6681 3249 6684
rect 3283 6712 3295 6715
rect 57514 6712 57520 6724
rect 3283 6684 57520 6712
rect 3283 6681 3295 6684
rect 3237 6675 3295 6681
rect 57514 6672 57520 6684
rect 57572 6672 57578 6724
rect 1946 6644 1952 6656
rect 1907 6616 1952 6644
rect 1946 6604 1952 6616
rect 2004 6604 2010 6656
rect 54018 6644 54024 6656
rect 53979 6616 54024 6644
rect 54018 6604 54024 6616
rect 54076 6604 54082 6656
rect 1104 6554 58880 6576
rect 1104 6502 10614 6554
rect 10666 6502 10678 6554
rect 10730 6502 10742 6554
rect 10794 6502 10806 6554
rect 10858 6502 29878 6554
rect 29930 6502 29942 6554
rect 29994 6502 30006 6554
rect 30058 6502 30070 6554
rect 30122 6502 49142 6554
rect 49194 6502 49206 6554
rect 49258 6502 49270 6554
rect 49322 6502 49334 6554
rect 49386 6502 58880 6554
rect 1104 6480 58880 6502
rect 1578 6236 1584 6248
rect 1539 6208 1584 6236
rect 1578 6196 1584 6208
rect 1636 6196 1642 6248
rect 1394 6168 1400 6180
rect 1355 6140 1400 6168
rect 1394 6128 1400 6140
rect 1452 6128 1458 6180
rect 57698 6100 57704 6112
rect 57659 6072 57704 6100
rect 57698 6060 57704 6072
rect 57756 6060 57762 6112
rect 1104 6010 58880 6032
rect 1104 5958 20246 6010
rect 20298 5958 20310 6010
rect 20362 5958 20374 6010
rect 20426 5958 20438 6010
rect 20490 5958 39510 6010
rect 39562 5958 39574 6010
rect 39626 5958 39638 6010
rect 39690 5958 39702 6010
rect 39754 5958 58880 6010
rect 1104 5936 58880 5958
rect 1762 5788 1768 5840
rect 1820 5828 1826 5840
rect 33962 5828 33968 5840
rect 1820 5800 33968 5828
rect 1820 5788 1826 5800
rect 33962 5788 33968 5800
rect 34020 5788 34026 5840
rect 56870 5720 56876 5772
rect 56928 5760 56934 5772
rect 57698 5760 57704 5772
rect 56928 5732 57704 5760
rect 56928 5720 56934 5732
rect 57698 5720 57704 5732
rect 57756 5760 57762 5772
rect 57977 5763 58035 5769
rect 57977 5760 57989 5763
rect 57756 5732 57989 5760
rect 57756 5720 57762 5732
rect 57977 5729 57989 5732
rect 58023 5729 58035 5763
rect 57977 5723 58035 5729
rect 58158 5624 58164 5636
rect 58119 5596 58164 5624
rect 58158 5584 58164 5596
rect 58216 5584 58222 5636
rect 40402 5516 40408 5568
rect 40460 5556 40466 5568
rect 40773 5559 40831 5565
rect 40773 5556 40785 5559
rect 40460 5528 40785 5556
rect 40460 5516 40466 5528
rect 40773 5525 40785 5528
rect 40819 5556 40831 5559
rect 53466 5556 53472 5568
rect 40819 5528 53472 5556
rect 40819 5525 40831 5528
rect 40773 5519 40831 5525
rect 53466 5516 53472 5528
rect 53524 5516 53530 5568
rect 57054 5556 57060 5568
rect 57015 5528 57060 5556
rect 57054 5516 57060 5528
rect 57112 5516 57118 5568
rect 1104 5466 58880 5488
rect 1104 5414 10614 5466
rect 10666 5414 10678 5466
rect 10730 5414 10742 5466
rect 10794 5414 10806 5466
rect 10858 5414 29878 5466
rect 29930 5414 29942 5466
rect 29994 5414 30006 5466
rect 30058 5414 30070 5466
rect 30122 5414 49142 5466
rect 49194 5414 49206 5466
rect 49258 5414 49270 5466
rect 49322 5414 49334 5466
rect 49386 5414 58880 5466
rect 1104 5392 58880 5414
rect 16850 5312 16856 5364
rect 16908 5352 16914 5364
rect 17037 5355 17095 5361
rect 17037 5352 17049 5355
rect 16908 5324 17049 5352
rect 16908 5312 16914 5324
rect 17037 5321 17049 5324
rect 17083 5352 17095 5355
rect 33962 5352 33968 5364
rect 17083 5324 24486 5352
rect 33923 5324 33968 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 1578 5244 1584 5296
rect 1636 5284 1642 5296
rect 2041 5287 2099 5293
rect 2041 5284 2053 5287
rect 1636 5256 2053 5284
rect 1636 5244 1642 5256
rect 2041 5253 2053 5256
rect 2087 5284 2099 5287
rect 18138 5284 18144 5296
rect 2087 5256 18144 5284
rect 2087 5253 2099 5256
rect 2041 5247 2099 5253
rect 18138 5244 18144 5256
rect 18196 5244 18202 5296
rect 24458 5284 24486 5324
rect 33962 5312 33968 5324
rect 34020 5312 34026 5364
rect 36078 5352 36084 5364
rect 34072 5324 36084 5352
rect 34072 5284 34100 5324
rect 36078 5312 36084 5324
rect 36136 5312 36142 5364
rect 24458 5256 34100 5284
rect 34790 5216 34796 5228
rect 34751 5188 34796 5216
rect 34790 5176 34796 5188
rect 34848 5176 34854 5228
rect 35713 5219 35771 5225
rect 35713 5185 35725 5219
rect 35759 5216 35771 5219
rect 39577 5219 39635 5225
rect 39577 5216 39589 5219
rect 35759 5188 39589 5216
rect 35759 5185 35771 5188
rect 35713 5179 35771 5185
rect 39577 5185 39589 5188
rect 39623 5216 39635 5219
rect 40221 5219 40279 5225
rect 40221 5216 40233 5219
rect 39623 5188 40233 5216
rect 39623 5185 39635 5188
rect 39577 5179 39635 5185
rect 40221 5185 40233 5188
rect 40267 5216 40279 5219
rect 41322 5216 41328 5228
rect 40267 5188 41328 5216
rect 40267 5185 40279 5188
rect 40221 5179 40279 5185
rect 21910 5108 21916 5160
rect 21968 5148 21974 5160
rect 25317 5151 25375 5157
rect 25317 5148 25329 5151
rect 21968 5120 25329 5148
rect 21968 5108 21974 5120
rect 25317 5117 25329 5120
rect 25363 5117 25375 5151
rect 25317 5111 25375 5117
rect 25409 5151 25467 5157
rect 25409 5117 25421 5151
rect 25455 5148 25467 5151
rect 25774 5148 25780 5160
rect 25455 5120 25780 5148
rect 25455 5117 25467 5120
rect 25409 5111 25467 5117
rect 25774 5108 25780 5120
rect 25832 5108 25838 5160
rect 34609 5151 34667 5157
rect 34609 5117 34621 5151
rect 34655 5148 34667 5151
rect 35728 5148 35756 5179
rect 41322 5176 41328 5188
rect 41380 5176 41386 5228
rect 41417 5219 41475 5225
rect 41417 5185 41429 5219
rect 41463 5216 41475 5219
rect 41506 5216 41512 5228
rect 41463 5188 41512 5216
rect 41463 5185 41475 5188
rect 41417 5179 41475 5185
rect 41506 5176 41512 5188
rect 41564 5176 41570 5228
rect 56410 5216 56416 5228
rect 56371 5188 56416 5216
rect 56410 5176 56416 5188
rect 56468 5176 56474 5228
rect 57517 5219 57575 5225
rect 57517 5185 57529 5219
rect 57563 5185 57575 5219
rect 57517 5179 57575 5185
rect 34655 5120 35756 5148
rect 57532 5148 57560 5179
rect 57790 5148 57796 5160
rect 57532 5120 57796 5148
rect 34655 5117 34667 5120
rect 34609 5111 34667 5117
rect 57790 5108 57796 5120
rect 57848 5148 57854 5160
rect 58161 5151 58219 5157
rect 58161 5148 58173 5151
rect 57848 5120 58173 5148
rect 57848 5108 57854 5120
rect 58161 5117 58173 5120
rect 58207 5117 58219 5151
rect 58161 5111 58219 5117
rect 56686 5040 56692 5092
rect 56744 5080 56750 5092
rect 56744 5052 58020 5080
rect 56744 5040 56750 5052
rect 1394 5012 1400 5024
rect 1355 4984 1400 5012
rect 1394 4972 1400 4984
rect 1452 4972 1458 5024
rect 33962 4972 33968 5024
rect 34020 5012 34026 5024
rect 34701 5015 34759 5021
rect 34701 5012 34713 5015
rect 34020 4984 34713 5012
rect 34020 4972 34026 4984
rect 34701 4981 34713 4984
rect 34747 4981 34759 5015
rect 34701 4975 34759 4981
rect 35179 5015 35237 5021
rect 35179 4981 35191 5015
rect 35225 5012 35237 5015
rect 35618 5012 35624 5024
rect 35225 4984 35624 5012
rect 35225 4981 35237 4984
rect 35179 4975 35237 4981
rect 35618 4972 35624 4984
rect 35676 4972 35682 5024
rect 40494 4972 40500 5024
rect 40552 5012 40558 5024
rect 40773 5015 40831 5021
rect 40773 5012 40785 5015
rect 40552 4984 40785 5012
rect 40552 4972 40558 4984
rect 40773 4981 40785 4984
rect 40819 4981 40831 5015
rect 40773 4975 40831 4981
rect 56965 5015 57023 5021
rect 56965 4981 56977 5015
rect 57011 5012 57023 5015
rect 57606 5012 57612 5024
rect 57011 4984 57612 5012
rect 57011 4981 57023 4984
rect 56965 4975 57023 4981
rect 57606 4972 57612 4984
rect 57664 4972 57670 5024
rect 57992 5021 58020 5052
rect 57977 5015 58035 5021
rect 57977 4981 57989 5015
rect 58023 4981 58035 5015
rect 57977 4975 58035 4981
rect 1104 4922 58880 4944
rect 1104 4870 20246 4922
rect 20298 4870 20310 4922
rect 20362 4870 20374 4922
rect 20426 4870 20438 4922
rect 20490 4870 39510 4922
rect 39562 4870 39574 4922
rect 39626 4870 39638 4922
rect 39690 4870 39702 4922
rect 39754 4870 58880 4922
rect 1104 4848 58880 4870
rect 2406 4808 2412 4820
rect 2367 4780 2412 4808
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 26234 4768 26240 4820
rect 26292 4808 26298 4820
rect 26421 4811 26479 4817
rect 26421 4808 26433 4811
rect 26292 4780 26433 4808
rect 26292 4768 26298 4780
rect 26421 4777 26433 4780
rect 26467 4777 26479 4811
rect 26421 4771 26479 4777
rect 35618 4768 35624 4820
rect 35676 4808 35682 4820
rect 56870 4808 56876 4820
rect 35676 4780 56876 4808
rect 35676 4768 35682 4780
rect 56870 4768 56876 4780
rect 56928 4768 56934 4820
rect 1394 4700 1400 4752
rect 1452 4740 1458 4752
rect 1489 4743 1547 4749
rect 1489 4740 1501 4743
rect 1452 4712 1501 4740
rect 1452 4700 1458 4712
rect 1489 4709 1501 4712
rect 1535 4709 1547 4743
rect 37642 4740 37648 4752
rect 37603 4712 37648 4740
rect 1489 4703 1547 4709
rect 37642 4700 37648 4712
rect 37700 4700 37706 4752
rect 41230 4700 41236 4752
rect 41288 4740 41294 4752
rect 42613 4743 42671 4749
rect 42613 4740 42625 4743
rect 41288 4712 42625 4740
rect 41288 4700 41294 4712
rect 42613 4709 42625 4712
rect 42659 4709 42671 4743
rect 42613 4703 42671 4709
rect 56781 4743 56839 4749
rect 56781 4709 56793 4743
rect 56827 4740 56839 4743
rect 58066 4740 58072 4752
rect 56827 4712 58072 4740
rect 56827 4709 56839 4712
rect 56781 4703 56839 4709
rect 58066 4700 58072 4712
rect 58124 4700 58130 4752
rect 27430 4672 27436 4684
rect 27343 4644 27436 4672
rect 27430 4632 27436 4644
rect 27488 4672 27494 4684
rect 29917 4675 29975 4681
rect 29917 4672 29929 4675
rect 27488 4644 29929 4672
rect 27488 4632 27494 4644
rect 29917 4641 29929 4644
rect 29963 4641 29975 4675
rect 29917 4635 29975 4641
rect 40494 4632 40500 4684
rect 40552 4672 40558 4684
rect 40957 4675 41015 4681
rect 40957 4672 40969 4675
rect 40552 4644 40969 4672
rect 40552 4632 40558 4644
rect 40957 4641 40969 4644
rect 41003 4641 41015 4675
rect 40957 4635 41015 4641
rect 57425 4675 57483 4681
rect 57425 4641 57437 4675
rect 57471 4672 57483 4675
rect 57606 4672 57612 4684
rect 57471 4644 57612 4672
rect 57471 4641 57483 4644
rect 57425 4635 57483 4641
rect 57606 4632 57612 4644
rect 57664 4632 57670 4684
rect 28718 4564 28724 4616
rect 28776 4604 28782 4616
rect 29273 4607 29331 4613
rect 29273 4604 29285 4607
rect 28776 4576 29285 4604
rect 28776 4564 28782 4576
rect 29273 4573 29285 4576
rect 29319 4604 29331 4607
rect 38470 4604 38476 4616
rect 29319 4576 38476 4604
rect 29319 4573 29331 4576
rect 29273 4567 29331 4573
rect 38470 4564 38476 4576
rect 38528 4564 38534 4616
rect 41138 4564 41144 4616
rect 41196 4604 41202 4616
rect 41414 4604 41420 4616
rect 41196 4576 41420 4604
rect 41196 4564 41202 4576
rect 41414 4564 41420 4576
rect 41472 4564 41478 4616
rect 1673 4539 1731 4545
rect 1673 4505 1685 4539
rect 1719 4536 1731 4539
rect 10226 4536 10232 4548
rect 1719 4508 10232 4536
rect 1719 4505 1731 4508
rect 1673 4499 1731 4505
rect 10226 4496 10232 4508
rect 10284 4496 10290 4548
rect 27706 4496 27712 4548
rect 27764 4536 27770 4548
rect 38749 4539 38807 4545
rect 38749 4536 38761 4539
rect 27764 4508 38761 4536
rect 27764 4496 27770 4508
rect 38749 4505 38761 4508
rect 38795 4536 38807 4539
rect 39114 4536 39120 4548
rect 38795 4508 39120 4536
rect 38795 4505 38807 4508
rect 38749 4499 38807 4505
rect 39114 4496 39120 4508
rect 39172 4496 39178 4548
rect 39850 4496 39856 4548
rect 39908 4536 39914 4548
rect 41046 4536 41052 4548
rect 39908 4508 41052 4536
rect 39908 4496 39914 4508
rect 41046 4496 41052 4508
rect 41104 4496 41110 4548
rect 41322 4496 41328 4548
rect 41380 4536 41386 4548
rect 41380 4508 43300 4536
rect 41380 4496 41386 4508
rect 15841 4471 15899 4477
rect 15841 4437 15853 4471
rect 15887 4468 15899 4471
rect 16022 4468 16028 4480
rect 15887 4440 16028 4468
rect 15887 4437 15899 4440
rect 15841 4431 15899 4437
rect 16022 4428 16028 4440
rect 16080 4428 16086 4480
rect 16482 4468 16488 4480
rect 16443 4440 16488 4468
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 17497 4471 17555 4477
rect 17497 4437 17509 4471
rect 17543 4468 17555 4471
rect 17770 4468 17776 4480
rect 17543 4440 17776 4468
rect 17543 4437 17555 4440
rect 17497 4431 17555 4437
rect 17770 4428 17776 4440
rect 17828 4428 17834 4480
rect 20530 4428 20536 4480
rect 20588 4468 20594 4480
rect 27246 4468 27252 4480
rect 20588 4440 27252 4468
rect 20588 4428 20594 4440
rect 27246 4428 27252 4440
rect 27304 4428 27310 4480
rect 28721 4471 28779 4477
rect 28721 4437 28733 4471
rect 28767 4468 28779 4471
rect 28810 4468 28816 4480
rect 28767 4440 28816 4468
rect 28767 4437 28779 4440
rect 28721 4431 28779 4437
rect 28810 4428 28816 4440
rect 28868 4428 28874 4480
rect 29917 4471 29975 4477
rect 29917 4437 29929 4471
rect 29963 4468 29975 4471
rect 36354 4468 36360 4480
rect 29963 4440 36360 4468
rect 29963 4437 29975 4440
rect 29917 4431 29975 4437
rect 36354 4428 36360 4440
rect 36412 4428 36418 4480
rect 36814 4428 36820 4480
rect 36872 4468 36878 4480
rect 37093 4471 37151 4477
rect 37093 4468 37105 4471
rect 36872 4440 37105 4468
rect 36872 4428 36878 4440
rect 37093 4437 37105 4440
rect 37139 4437 37151 4471
rect 37093 4431 37151 4437
rect 39298 4428 39304 4480
rect 39356 4468 39362 4480
rect 39761 4471 39819 4477
rect 39761 4468 39773 4471
rect 39356 4440 39773 4468
rect 39356 4428 39362 4440
rect 39761 4437 39773 4440
rect 39807 4437 39819 4471
rect 41138 4468 41144 4480
rect 41099 4440 41144 4468
rect 39761 4431 39819 4437
rect 41138 4428 41144 4440
rect 41196 4428 41202 4480
rect 42153 4471 42211 4477
rect 42153 4437 42165 4471
rect 42199 4468 42211 4471
rect 42426 4468 42432 4480
rect 42199 4440 42432 4468
rect 42199 4437 42211 4440
rect 42153 4431 42211 4437
rect 42426 4428 42432 4440
rect 42484 4428 42490 4480
rect 43272 4477 43300 4508
rect 44082 4496 44088 4548
rect 44140 4536 44146 4548
rect 52362 4536 52368 4548
rect 44140 4508 52368 4536
rect 44140 4496 44146 4508
rect 52362 4496 52368 4508
rect 52420 4496 52426 4548
rect 57882 4536 57888 4548
rect 57843 4508 57888 4536
rect 57882 4496 57888 4508
rect 57940 4496 57946 4548
rect 43257 4471 43315 4477
rect 43257 4437 43269 4471
rect 43303 4468 43315 4471
rect 43809 4471 43867 4477
rect 43809 4468 43821 4471
rect 43303 4440 43821 4468
rect 43303 4437 43315 4440
rect 43257 4431 43315 4437
rect 43809 4437 43821 4440
rect 43855 4468 43867 4471
rect 44361 4471 44419 4477
rect 44361 4468 44373 4471
rect 43855 4440 44373 4468
rect 43855 4437 43867 4440
rect 43809 4431 43867 4437
rect 44361 4437 44373 4440
rect 44407 4468 44419 4471
rect 44634 4468 44640 4480
rect 44407 4440 44640 4468
rect 44407 4437 44419 4440
rect 44361 4431 44419 4437
rect 44634 4428 44640 4440
rect 44692 4428 44698 4480
rect 57238 4468 57244 4480
rect 57199 4440 57244 4468
rect 57238 4428 57244 4440
rect 57296 4428 57302 4480
rect 1104 4378 58880 4400
rect 1104 4326 10614 4378
rect 10666 4326 10678 4378
rect 10730 4326 10742 4378
rect 10794 4326 10806 4378
rect 10858 4326 29878 4378
rect 29930 4326 29942 4378
rect 29994 4326 30006 4378
rect 30058 4326 30070 4378
rect 30122 4326 49142 4378
rect 49194 4326 49206 4378
rect 49258 4326 49270 4378
rect 49322 4326 49334 4378
rect 49386 4326 58880 4378
rect 1104 4304 58880 4326
rect 3789 4267 3847 4273
rect 3789 4233 3801 4267
rect 3835 4264 3847 4267
rect 4246 4264 4252 4276
rect 3835 4236 4252 4264
rect 3835 4233 3847 4236
rect 3789 4227 3847 4233
rect 4246 4224 4252 4236
rect 4304 4224 4310 4276
rect 10318 4264 10324 4276
rect 10279 4236 10324 4264
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 19337 4267 19395 4273
rect 19337 4233 19349 4267
rect 19383 4264 19395 4267
rect 19426 4264 19432 4276
rect 19383 4236 19432 4264
rect 19383 4233 19395 4236
rect 19337 4227 19395 4233
rect 19426 4224 19432 4236
rect 19484 4224 19490 4276
rect 21542 4224 21548 4276
rect 21600 4264 21606 4276
rect 21818 4264 21824 4276
rect 21600 4236 21824 4264
rect 21600 4224 21606 4236
rect 21818 4224 21824 4236
rect 21876 4264 21882 4276
rect 22741 4267 22799 4273
rect 22741 4264 22753 4267
rect 21876 4236 22753 4264
rect 21876 4224 21882 4236
rect 22741 4233 22753 4236
rect 22787 4233 22799 4267
rect 22741 4227 22799 4233
rect 24458 4236 25820 4264
rect 15381 4199 15439 4205
rect 15381 4165 15393 4199
rect 15427 4196 15439 4199
rect 24458 4196 24486 4236
rect 25682 4196 25688 4208
rect 15427 4168 24486 4196
rect 24596 4168 25688 4196
rect 15427 4165 15439 4168
rect 15381 4159 15439 4165
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 24596 4128 24624 4168
rect 25682 4156 25688 4168
rect 25740 4156 25746 4208
rect 25792 4196 25820 4236
rect 25866 4224 25872 4276
rect 25924 4264 25930 4276
rect 26329 4267 26387 4273
rect 26329 4264 26341 4267
rect 25924 4236 26341 4264
rect 25924 4224 25930 4236
rect 26329 4233 26341 4236
rect 26375 4233 26387 4267
rect 28902 4264 28908 4276
rect 28863 4236 28908 4264
rect 26329 4227 26387 4233
rect 28902 4224 28908 4236
rect 28960 4224 28966 4276
rect 29454 4264 29460 4276
rect 29415 4236 29460 4264
rect 29454 4224 29460 4236
rect 29512 4224 29518 4276
rect 36998 4264 37004 4276
rect 36959 4236 37004 4264
rect 36998 4224 37004 4236
rect 37056 4224 37062 4276
rect 40865 4267 40923 4273
rect 40865 4233 40877 4267
rect 40911 4264 40923 4267
rect 43622 4264 43628 4276
rect 40911 4236 43628 4264
rect 40911 4233 40923 4236
rect 40865 4227 40923 4233
rect 43622 4224 43628 4236
rect 43680 4224 43686 4276
rect 43990 4224 43996 4276
rect 44048 4264 44054 4276
rect 57238 4264 57244 4276
rect 44048 4236 57244 4264
rect 44048 4224 44054 4236
rect 57238 4224 57244 4236
rect 57296 4224 57302 4276
rect 57977 4267 58035 4273
rect 57977 4233 57989 4267
rect 58023 4264 58035 4267
rect 58250 4264 58256 4276
rect 58023 4236 58256 4264
rect 58023 4233 58035 4236
rect 57977 4227 58035 4233
rect 58250 4224 58256 4236
rect 58308 4224 58314 4276
rect 26970 4196 26976 4208
rect 25792 4168 26976 4196
rect 26970 4156 26976 4168
rect 27028 4156 27034 4208
rect 28810 4156 28816 4208
rect 28868 4196 28874 4208
rect 57882 4196 57888 4208
rect 28868 4168 57888 4196
rect 28868 4156 28874 4168
rect 57882 4156 57888 4168
rect 57940 4156 57946 4208
rect 25774 4128 25780 4140
rect 24458 4100 24624 4128
rect 25056 4100 25780 4128
rect 1578 4060 1584 4072
rect 1539 4032 1584 4060
rect 1578 4020 1584 4032
rect 1636 4020 1642 4072
rect 1946 4020 1952 4072
rect 2004 4060 2010 4072
rect 2317 4063 2375 4069
rect 2317 4060 2329 4063
rect 2004 4032 2329 4060
rect 2004 4020 2010 4032
rect 2317 4029 2329 4032
rect 2363 4029 2375 4063
rect 15194 4060 15200 4072
rect 15155 4032 15200 4060
rect 2317 4023 2375 4029
rect 15194 4020 15200 4032
rect 15252 4060 15258 4072
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15252 4032 15853 4060
rect 15252 4020 15258 4032
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 17586 4020 17592 4072
rect 17644 4060 17650 4072
rect 17681 4063 17739 4069
rect 17681 4060 17693 4063
rect 17644 4032 17693 4060
rect 17644 4020 17650 4032
rect 17681 4029 17693 4032
rect 17727 4060 17739 4063
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 17727 4032 18153 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 18141 4029 18153 4032
rect 18187 4029 18199 4063
rect 18141 4023 18199 4029
rect 1302 3952 1308 4004
rect 1360 3992 1366 4004
rect 2133 3995 2191 4001
rect 2133 3992 2145 3995
rect 1360 3964 2145 3992
rect 1360 3952 1366 3964
rect 2133 3961 2145 3964
rect 2179 3961 2191 3995
rect 2133 3955 2191 3961
rect 16666 3952 16672 4004
rect 16724 3992 16730 4004
rect 17037 3995 17095 4001
rect 17037 3992 17049 3995
rect 16724 3964 17049 3992
rect 16724 3952 16730 3964
rect 17037 3961 17049 3964
rect 17083 3992 17095 3995
rect 24458 3992 24486 4100
rect 25056 4072 25084 4100
rect 25774 4088 25780 4100
rect 25832 4088 25838 4140
rect 27246 4088 27252 4140
rect 27304 4128 27310 4140
rect 27304 4100 44220 4128
rect 27304 4088 27310 4100
rect 25038 4060 25044 4072
rect 24999 4032 25044 4060
rect 25038 4020 25044 4032
rect 25096 4020 25102 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4029 25283 4063
rect 25682 4060 25688 4072
rect 25643 4032 25688 4060
rect 25225 4023 25283 4029
rect 17083 3964 24486 3992
rect 24581 3995 24639 4001
rect 17083 3961 17095 3964
rect 17037 3955 17095 3961
rect 24581 3961 24593 3995
rect 24627 3992 24639 3995
rect 25240 3992 25268 4023
rect 25682 4020 25688 4032
rect 25740 4020 25746 4072
rect 25866 4060 25872 4072
rect 25827 4032 25872 4060
rect 25866 4020 25872 4032
rect 25924 4020 25930 4072
rect 34606 4060 34612 4072
rect 33474 4032 34612 4060
rect 33474 3992 33502 4032
rect 34606 4020 34612 4032
rect 34664 4020 34670 4072
rect 36814 4060 36820 4072
rect 36775 4032 36820 4060
rect 36814 4020 36820 4032
rect 36872 4020 36878 4072
rect 37458 4060 37464 4072
rect 37292 4032 37464 4060
rect 24627 3964 33502 3992
rect 24627 3961 24639 3964
rect 24581 3955 24639 3961
rect 36078 3952 36084 4004
rect 36136 3992 36142 4004
rect 36173 3995 36231 4001
rect 36173 3992 36185 3995
rect 36136 3964 36185 3992
rect 36136 3952 36142 3964
rect 36173 3961 36185 3964
rect 36219 3992 36231 3995
rect 37292 3992 37320 4032
rect 37458 4020 37464 4032
rect 37516 4060 37522 4072
rect 39390 4060 39396 4072
rect 37516 4032 39396 4060
rect 37516 4020 37522 4032
rect 39390 4020 39396 4032
rect 39448 4020 39454 4072
rect 39850 4020 39856 4072
rect 39908 4060 39914 4072
rect 40037 4063 40095 4069
rect 40037 4060 40049 4063
rect 39908 4032 40049 4060
rect 39908 4020 39914 4032
rect 40037 4029 40049 4032
rect 40083 4029 40095 4063
rect 40037 4023 40095 4029
rect 40221 4063 40279 4069
rect 40221 4029 40233 4063
rect 40267 4060 40279 4063
rect 40865 4063 40923 4069
rect 40865 4060 40877 4063
rect 40267 4032 40877 4060
rect 40267 4029 40279 4032
rect 40221 4023 40279 4029
rect 40865 4029 40877 4032
rect 40911 4029 40923 4063
rect 40865 4023 40923 4029
rect 40957 4063 41015 4069
rect 40957 4029 40969 4063
rect 41003 4060 41015 4063
rect 41046 4060 41052 4072
rect 41003 4032 41052 4060
rect 41003 4029 41015 4032
rect 40957 4023 41015 4029
rect 41046 4020 41052 4032
rect 41104 4020 41110 4072
rect 41141 4063 41199 4069
rect 41141 4029 41153 4063
rect 41187 4060 41199 4063
rect 41414 4060 41420 4072
rect 41187 4032 41420 4060
rect 41187 4029 41199 4032
rect 41141 4023 41199 4029
rect 41414 4020 41420 4032
rect 41472 4060 41478 4072
rect 41693 4063 41751 4069
rect 41693 4060 41705 4063
rect 41472 4032 41705 4060
rect 41472 4020 41478 4032
rect 41693 4029 41705 4032
rect 41739 4029 41751 4063
rect 41693 4023 41751 4029
rect 41785 4063 41843 4069
rect 41785 4029 41797 4063
rect 41831 4029 41843 4063
rect 42426 4060 42432 4072
rect 42387 4032 42432 4060
rect 41785 4023 41843 4029
rect 36219 3964 37320 3992
rect 36219 3961 36231 3964
rect 36173 3955 36231 3961
rect 37366 3952 37372 4004
rect 37424 3992 37430 4004
rect 41800 3992 41828 4023
rect 42426 4020 42432 4032
rect 42484 4020 42490 4072
rect 43806 4020 43812 4072
rect 43864 4060 43870 4072
rect 44082 4060 44088 4072
rect 43864 4032 44088 4060
rect 43864 4020 43870 4032
rect 44082 4020 44088 4032
rect 44140 4020 44146 4072
rect 44192 4060 44220 4100
rect 44266 4088 44272 4140
rect 44324 4128 44330 4140
rect 45189 4131 45247 4137
rect 45189 4128 45201 4131
rect 44324 4100 45201 4128
rect 44324 4088 44330 4100
rect 45189 4097 45201 4100
rect 45235 4128 45247 4131
rect 48406 4128 48412 4140
rect 45235 4100 48412 4128
rect 45235 4097 45247 4100
rect 45189 4091 45247 4097
rect 48406 4088 48412 4100
rect 48464 4088 48470 4140
rect 55122 4128 55128 4140
rect 55083 4100 55128 4128
rect 55122 4088 55128 4100
rect 55180 4128 55186 4140
rect 57974 4128 57980 4140
rect 55180 4100 57980 4128
rect 55180 4088 55186 4100
rect 57974 4088 57980 4100
rect 58032 4088 58038 4140
rect 47118 4060 47124 4072
rect 44192 4032 47124 4060
rect 47118 4020 47124 4032
rect 47176 4020 47182 4072
rect 56321 4063 56379 4069
rect 56321 4029 56333 4063
rect 56367 4060 56379 4063
rect 57333 4063 57391 4069
rect 57333 4060 57345 4063
rect 56367 4032 57345 4060
rect 56367 4029 56379 4032
rect 56321 4023 56379 4029
rect 57333 4029 57345 4032
rect 57379 4060 57391 4063
rect 57790 4060 57796 4072
rect 57379 4032 57796 4060
rect 57379 4029 57391 4032
rect 57333 4023 57391 4029
rect 57790 4020 57796 4032
rect 57848 4020 57854 4072
rect 57882 4020 57888 4072
rect 57940 4060 57946 4072
rect 58161 4063 58219 4069
rect 58161 4060 58173 4063
rect 57940 4032 58173 4060
rect 57940 4020 57946 4032
rect 58161 4029 58173 4032
rect 58207 4029 58219 4063
rect 58161 4023 58219 4029
rect 45462 3992 45468 4004
rect 37424 3964 41736 3992
rect 41800 3964 45468 3992
rect 37424 3952 37430 3964
rect 3142 3924 3148 3936
rect 3103 3896 3148 3924
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 17402 3884 17408 3936
rect 17460 3924 17466 3936
rect 17497 3927 17555 3933
rect 17497 3924 17509 3927
rect 17460 3896 17509 3924
rect 17460 3884 17466 3896
rect 17497 3893 17509 3896
rect 17543 3893 17555 3927
rect 18690 3924 18696 3936
rect 18651 3896 18696 3924
rect 17497 3887 17555 3893
rect 18690 3884 18696 3896
rect 18748 3884 18754 3936
rect 21174 3924 21180 3936
rect 21135 3896 21180 3924
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 25130 3924 25136 3936
rect 25091 3896 25136 3924
rect 25130 3884 25136 3896
rect 25188 3884 25194 3936
rect 25777 3927 25835 3933
rect 25777 3893 25789 3927
rect 25823 3924 25835 3927
rect 25958 3924 25964 3936
rect 25823 3896 25964 3924
rect 25823 3893 25835 3896
rect 25777 3887 25835 3893
rect 25958 3884 25964 3896
rect 26016 3884 26022 3936
rect 27614 3924 27620 3936
rect 27575 3896 27620 3924
rect 27614 3884 27620 3896
rect 27672 3884 27678 3936
rect 28074 3884 28080 3936
rect 28132 3924 28138 3936
rect 28169 3927 28227 3933
rect 28169 3924 28181 3927
rect 28132 3896 28181 3924
rect 28132 3884 28138 3896
rect 28169 3893 28181 3896
rect 28215 3893 28227 3927
rect 28169 3887 28227 3893
rect 34974 3884 34980 3936
rect 35032 3924 35038 3936
rect 35529 3927 35587 3933
rect 35529 3924 35541 3927
rect 35032 3896 35541 3924
rect 35032 3884 35038 3896
rect 35529 3893 35541 3896
rect 35575 3893 35587 3927
rect 35529 3887 35587 3893
rect 38194 3884 38200 3936
rect 38252 3924 38258 3936
rect 38289 3927 38347 3933
rect 38289 3924 38301 3927
rect 38252 3896 38301 3924
rect 38252 3884 38258 3896
rect 38289 3893 38301 3896
rect 38335 3893 38347 3927
rect 38289 3887 38347 3893
rect 38654 3884 38660 3936
rect 38712 3924 38718 3936
rect 38933 3927 38991 3933
rect 38933 3924 38945 3927
rect 38712 3896 38945 3924
rect 38712 3884 38718 3896
rect 38933 3893 38945 3896
rect 38979 3893 38991 3927
rect 38933 3887 38991 3893
rect 39390 3884 39396 3936
rect 39448 3924 39454 3936
rect 39485 3927 39543 3933
rect 39485 3924 39497 3927
rect 39448 3896 39497 3924
rect 39448 3884 39454 3896
rect 39485 3893 39497 3896
rect 39531 3893 39543 3927
rect 40126 3924 40132 3936
rect 40087 3896 40132 3924
rect 39485 3887 39543 3893
rect 40126 3884 40132 3896
rect 40184 3884 40190 3936
rect 41049 3927 41107 3933
rect 41049 3893 41061 3927
rect 41095 3924 41107 3927
rect 41598 3924 41604 3936
rect 41095 3896 41604 3924
rect 41095 3893 41107 3896
rect 41049 3887 41107 3893
rect 41598 3884 41604 3896
rect 41656 3884 41662 3936
rect 41708 3924 41736 3964
rect 45462 3952 45468 3964
rect 45520 3952 45526 4004
rect 45554 3952 45560 4004
rect 45612 3992 45618 4004
rect 45741 3995 45799 4001
rect 45741 3992 45753 3995
rect 45612 3964 45753 3992
rect 45612 3952 45618 3964
rect 45741 3961 45753 3964
rect 45787 3992 45799 3995
rect 51074 3992 51080 4004
rect 45787 3964 51080 3992
rect 45787 3961 45799 3964
rect 45741 3955 45799 3961
rect 51074 3952 51080 3964
rect 51132 3952 51138 4004
rect 56873 3995 56931 4001
rect 56873 3961 56885 3995
rect 56919 3992 56931 3995
rect 57900 3992 57928 4020
rect 56919 3964 57928 3992
rect 56919 3961 56931 3964
rect 56873 3955 56931 3961
rect 42245 3927 42303 3933
rect 42245 3924 42257 3927
rect 41708 3896 42257 3924
rect 42245 3893 42257 3896
rect 42291 3893 42303 3927
rect 43438 3924 43444 3936
rect 43399 3896 43444 3924
rect 42245 3887 42303 3893
rect 43438 3884 43444 3896
rect 43496 3884 43502 3936
rect 44542 3924 44548 3936
rect 44503 3896 44548 3924
rect 44542 3884 44548 3896
rect 44600 3884 44606 3936
rect 44634 3884 44640 3936
rect 44692 3924 44698 3936
rect 46290 3924 46296 3936
rect 44692 3896 46296 3924
rect 44692 3884 44698 3896
rect 46290 3884 46296 3896
rect 46348 3884 46354 3936
rect 46845 3927 46903 3933
rect 46845 3893 46857 3927
rect 46891 3924 46903 3927
rect 47302 3924 47308 3936
rect 46891 3896 47308 3924
rect 46891 3893 46903 3896
rect 46845 3887 46903 3893
rect 47302 3884 47308 3896
rect 47360 3884 47366 3936
rect 47578 3924 47584 3936
rect 47539 3896 47584 3924
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 55582 3884 55588 3936
rect 55640 3924 55646 3936
rect 55677 3927 55735 3933
rect 55677 3924 55689 3927
rect 55640 3896 55689 3924
rect 55640 3884 55646 3896
rect 55677 3893 55689 3896
rect 55723 3893 55735 3927
rect 57514 3924 57520 3936
rect 57475 3896 57520 3924
rect 55677 3887 55735 3893
rect 57514 3884 57520 3896
rect 57572 3884 57578 3936
rect 1104 3834 58880 3856
rect 1104 3782 20246 3834
rect 20298 3782 20310 3834
rect 20362 3782 20374 3834
rect 20426 3782 20438 3834
rect 20490 3782 39510 3834
rect 39562 3782 39574 3834
rect 39626 3782 39638 3834
rect 39690 3782 39702 3834
rect 39754 3782 58880 3834
rect 1104 3760 58880 3782
rect 11514 3720 11520 3732
rect 11475 3692 11520 3720
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 14366 3720 14372 3732
rect 14327 3692 14372 3720
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 15470 3680 15476 3732
rect 15528 3720 15534 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15528 3692 15577 3720
rect 15528 3680 15534 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 22554 3720 22560 3732
rect 22515 3692 22560 3720
rect 15565 3683 15623 3689
rect 22554 3680 22560 3692
rect 22612 3680 22618 3732
rect 25774 3720 25780 3732
rect 25735 3692 25780 3720
rect 25774 3680 25780 3692
rect 25832 3680 25838 3732
rect 30466 3720 30472 3732
rect 30427 3692 30472 3720
rect 30466 3680 30472 3692
rect 30524 3680 30530 3732
rect 31202 3680 31208 3732
rect 31260 3720 31266 3732
rect 31665 3723 31723 3729
rect 31665 3720 31677 3723
rect 31260 3692 31677 3720
rect 31260 3680 31266 3692
rect 31665 3689 31677 3692
rect 31711 3689 31723 3723
rect 32398 3720 32404 3732
rect 32359 3692 32404 3720
rect 31665 3683 31723 3689
rect 32398 3680 32404 3692
rect 32456 3680 32462 3732
rect 34790 3680 34796 3732
rect 34848 3720 34854 3732
rect 35713 3723 35771 3729
rect 35713 3720 35725 3723
rect 34848 3692 35725 3720
rect 34848 3680 34854 3692
rect 35713 3689 35725 3692
rect 35759 3689 35771 3723
rect 35713 3683 35771 3689
rect 38746 3680 38752 3732
rect 38804 3720 38810 3732
rect 38841 3723 38899 3729
rect 38841 3720 38853 3723
rect 38804 3692 38853 3720
rect 38804 3680 38810 3692
rect 38841 3689 38853 3692
rect 38887 3689 38899 3723
rect 38841 3683 38899 3689
rect 41414 3680 41420 3732
rect 41472 3720 41478 3732
rect 42426 3720 42432 3732
rect 41472 3692 42432 3720
rect 41472 3680 41478 3692
rect 42426 3680 42432 3692
rect 42484 3680 42490 3732
rect 43622 3680 43628 3732
rect 43680 3720 43686 3732
rect 43901 3723 43959 3729
rect 43901 3720 43913 3723
rect 43680 3692 43913 3720
rect 43680 3680 43686 3692
rect 43901 3689 43913 3692
rect 43947 3689 43959 3723
rect 43901 3683 43959 3689
rect 2038 3612 2044 3664
rect 2096 3652 2102 3664
rect 2317 3655 2375 3661
rect 2317 3652 2329 3655
rect 2096 3624 2329 3652
rect 2096 3612 2102 3624
rect 2317 3621 2329 3624
rect 2363 3621 2375 3655
rect 2317 3615 2375 3621
rect 3053 3655 3111 3661
rect 3053 3621 3065 3655
rect 3099 3652 3111 3655
rect 4246 3652 4252 3664
rect 3099 3624 4252 3652
rect 3099 3621 3111 3624
rect 3053 3615 3111 3621
rect 4246 3612 4252 3624
rect 4304 3612 4310 3664
rect 11054 3652 11060 3664
rect 6426 3624 11060 3652
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 1627 3556 4445 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 4433 3553 4445 3556
rect 4479 3584 4491 3587
rect 6426 3584 6454 3624
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 4479 3556 6454 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 9214 3544 9220 3596
rect 9272 3584 9278 3596
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 9272 3556 9505 3584
rect 9272 3544 9278 3556
rect 9493 3553 9505 3556
rect 9539 3584 9551 3587
rect 10137 3587 10195 3593
rect 10137 3584 10149 3587
rect 9539 3556 10149 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 10137 3553 10149 3556
rect 10183 3553 10195 3587
rect 14384 3584 14412 3680
rect 16482 3652 16488 3664
rect 16316 3624 16488 3652
rect 14921 3587 14979 3593
rect 14921 3584 14933 3587
rect 14384 3556 14933 3584
rect 10137 3547 10195 3553
rect 14921 3553 14933 3556
rect 14967 3553 14979 3587
rect 14921 3547 14979 3553
rect 15105 3587 15163 3593
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15378 3584 15384 3596
rect 15151 3556 15384 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15378 3544 15384 3556
rect 15436 3584 15442 3596
rect 16316 3593 16344 3624
rect 16482 3612 16488 3624
rect 16540 3652 16546 3664
rect 47857 3655 47915 3661
rect 47857 3652 47869 3655
rect 16540 3624 47869 3652
rect 16540 3612 16546 3624
rect 47857 3621 47869 3624
rect 47903 3621 47915 3655
rect 57974 3652 57980 3664
rect 57935 3624 57980 3652
rect 47857 3615 47915 3621
rect 57974 3612 57980 3624
rect 58032 3612 58038 3664
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 15436 3556 16221 3584
rect 15436 3544 15442 3556
rect 16209 3553 16221 3556
rect 16255 3553 16267 3587
rect 16209 3547 16267 3553
rect 16301 3587 16359 3593
rect 16301 3553 16313 3587
rect 16347 3553 16359 3587
rect 16758 3584 16764 3596
rect 16719 3556 16764 3584
rect 16301 3547 16359 3553
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 17402 3584 17408 3596
rect 17363 3556 17408 3584
rect 17402 3544 17408 3556
rect 17460 3544 17466 3596
rect 18414 3584 18420 3596
rect 18327 3556 18420 3584
rect 18414 3544 18420 3556
rect 18472 3584 18478 3596
rect 18690 3584 18696 3596
rect 18472 3556 18696 3584
rect 18472 3544 18478 3556
rect 18690 3544 18696 3556
rect 18748 3544 18754 3596
rect 21174 3544 21180 3596
rect 21232 3584 21238 3596
rect 21232 3556 22232 3584
rect 21232 3544 21238 3556
rect 22204 3528 22232 3556
rect 22646 3544 22652 3596
rect 22704 3584 22710 3596
rect 22741 3587 22799 3593
rect 22741 3584 22753 3587
rect 22704 3556 22753 3584
rect 22704 3544 22710 3556
rect 22741 3553 22753 3556
rect 22787 3584 22799 3587
rect 23201 3587 23259 3593
rect 23201 3584 23213 3587
rect 22787 3556 23213 3584
rect 22787 3553 22799 3556
rect 22741 3547 22799 3553
rect 23201 3553 23213 3556
rect 23247 3553 23259 3587
rect 23201 3547 23259 3553
rect 25225 3587 25283 3593
rect 25225 3553 25237 3587
rect 25271 3584 25283 3587
rect 25869 3587 25927 3593
rect 25869 3584 25881 3587
rect 25271 3556 25881 3584
rect 25271 3553 25283 3556
rect 25225 3547 25283 3553
rect 25869 3553 25881 3556
rect 25915 3584 25927 3587
rect 26142 3584 26148 3596
rect 25915 3556 26148 3584
rect 25915 3553 25927 3556
rect 25869 3547 25927 3553
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 27341 3587 27399 3593
rect 27341 3553 27353 3587
rect 27387 3584 27399 3587
rect 27798 3584 27804 3596
rect 27387 3556 27804 3584
rect 27387 3553 27399 3556
rect 27341 3547 27399 3553
rect 27798 3544 27804 3556
rect 27856 3544 27862 3596
rect 27893 3587 27951 3593
rect 27893 3553 27905 3587
rect 27939 3584 27951 3587
rect 28074 3584 28080 3596
rect 27939 3556 28080 3584
rect 27939 3553 27951 3556
rect 27893 3547 27951 3553
rect 28074 3544 28080 3556
rect 28132 3544 28138 3596
rect 28718 3584 28724 3596
rect 28679 3556 28724 3584
rect 28718 3544 28724 3556
rect 28776 3544 28782 3596
rect 29273 3587 29331 3593
rect 29273 3553 29285 3587
rect 29319 3553 29331 3587
rect 29273 3547 29331 3553
rect 21910 3516 21916 3528
rect 11578 3488 21916 3516
rect 474 3408 480 3460
rect 532 3448 538 3460
rect 2869 3451 2927 3457
rect 2869 3448 2881 3451
rect 532 3420 2881 3448
rect 532 3408 538 3420
rect 2869 3417 2881 3420
rect 2915 3417 2927 3451
rect 2869 3411 2927 3417
rect 9677 3451 9735 3457
rect 9677 3417 9689 3451
rect 9723 3448 9735 3451
rect 11578 3448 11606 3488
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 22186 3476 22192 3528
rect 22244 3516 22250 3528
rect 27614 3516 27620 3528
rect 22244 3488 27620 3516
rect 22244 3476 22250 3488
rect 27614 3476 27620 3488
rect 27672 3476 27678 3528
rect 29288 3516 29316 3547
rect 30190 3544 30196 3596
rect 30248 3584 30254 3596
rect 30653 3587 30711 3593
rect 30653 3584 30665 3587
rect 30248 3556 30665 3584
rect 30248 3544 30254 3556
rect 30653 3553 30665 3556
rect 30699 3584 30711 3587
rect 31113 3587 31171 3593
rect 31113 3584 31125 3587
rect 30699 3556 31125 3584
rect 30699 3553 30711 3556
rect 30653 3547 30711 3553
rect 31113 3553 31125 3556
rect 31159 3553 31171 3587
rect 32214 3584 32220 3596
rect 32175 3556 32220 3584
rect 31113 3547 31171 3553
rect 32214 3544 32220 3556
rect 32272 3584 32278 3596
rect 32861 3587 32919 3593
rect 32861 3584 32873 3587
rect 32272 3556 32873 3584
rect 32272 3544 32278 3556
rect 32861 3553 32873 3556
rect 32907 3553 32919 3587
rect 34054 3584 34060 3596
rect 34015 3556 34060 3584
rect 32861 3547 32919 3553
rect 34054 3544 34060 3556
rect 34112 3584 34118 3596
rect 34701 3587 34759 3593
rect 34701 3584 34713 3587
rect 34112 3556 34713 3584
rect 34112 3544 34118 3556
rect 34701 3553 34713 3556
rect 34747 3553 34759 3587
rect 34701 3547 34759 3553
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 35897 3587 35955 3593
rect 35897 3584 35909 3587
rect 35032 3556 35909 3584
rect 35032 3544 35038 3556
rect 35897 3553 35909 3556
rect 35943 3553 35955 3587
rect 35897 3547 35955 3553
rect 36541 3587 36599 3593
rect 36541 3553 36553 3587
rect 36587 3584 36599 3587
rect 36630 3584 36636 3596
rect 36587 3556 36636 3584
rect 36587 3553 36599 3556
rect 36541 3547 36599 3553
rect 36630 3544 36636 3556
rect 36688 3544 36694 3596
rect 37277 3587 37335 3593
rect 37277 3553 37289 3587
rect 37323 3584 37335 3587
rect 37366 3584 37372 3596
rect 37323 3556 37372 3584
rect 37323 3553 37335 3556
rect 37277 3547 37335 3553
rect 37366 3544 37372 3556
rect 37424 3544 37430 3596
rect 38013 3587 38071 3593
rect 38013 3553 38025 3587
rect 38059 3584 38071 3587
rect 38194 3584 38200 3596
rect 38059 3556 38200 3584
rect 38059 3553 38071 3556
rect 38013 3547 38071 3553
rect 38194 3544 38200 3556
rect 38252 3544 38258 3596
rect 38654 3584 38660 3596
rect 38615 3556 38660 3584
rect 38654 3544 38660 3556
rect 38712 3544 38718 3596
rect 39761 3587 39819 3593
rect 39761 3553 39773 3587
rect 39807 3584 39819 3587
rect 40126 3584 40132 3596
rect 39807 3556 40132 3584
rect 39807 3553 39819 3556
rect 39761 3547 39819 3553
rect 40126 3544 40132 3556
rect 40184 3544 40190 3596
rect 41138 3584 41144 3596
rect 41099 3556 41144 3584
rect 41138 3544 41144 3556
rect 41196 3544 41202 3596
rect 41598 3544 41604 3596
rect 41656 3584 41662 3596
rect 42061 3587 42119 3593
rect 42061 3584 42073 3587
rect 41656 3556 42073 3584
rect 41656 3544 41662 3556
rect 42061 3553 42073 3556
rect 42107 3553 42119 3587
rect 42061 3547 42119 3553
rect 43349 3587 43407 3593
rect 43349 3553 43361 3587
rect 43395 3584 43407 3587
rect 43438 3584 43444 3596
rect 43395 3556 43444 3584
rect 43395 3553 43407 3556
rect 43349 3547 43407 3553
rect 43438 3544 43444 3556
rect 43496 3544 43502 3596
rect 43990 3584 43996 3596
rect 43951 3556 43996 3584
rect 43990 3544 43996 3556
rect 44048 3544 44054 3596
rect 44637 3587 44695 3593
rect 44637 3553 44649 3587
rect 44683 3553 44695 3587
rect 44637 3547 44695 3553
rect 48041 3587 48099 3593
rect 48041 3553 48053 3587
rect 48087 3553 48099 3587
rect 48041 3547 48099 3553
rect 28092 3488 29316 3516
rect 9723 3420 11606 3448
rect 16945 3451 17003 3457
rect 9723 3417 9735 3420
rect 9677 3411 9735 3417
rect 16945 3417 16957 3451
rect 16991 3448 17003 3451
rect 18138 3448 18144 3460
rect 16991 3420 18144 3448
rect 16991 3417 17003 3420
rect 16945 3411 17003 3417
rect 18138 3408 18144 3420
rect 18196 3408 18202 3460
rect 19426 3408 19432 3460
rect 19484 3448 19490 3460
rect 26326 3448 26332 3460
rect 19484 3420 26332 3448
rect 19484 3408 19490 3420
rect 26326 3408 26332 3420
rect 26384 3448 26390 3460
rect 26605 3451 26663 3457
rect 26605 3448 26617 3451
rect 26384 3420 26617 3448
rect 26384 3408 26390 3420
rect 26605 3417 26617 3420
rect 26651 3417 26663 3451
rect 27154 3448 27160 3460
rect 27115 3420 27160 3448
rect 26605 3411 26663 3417
rect 27154 3408 27160 3420
rect 27212 3408 27218 3460
rect 28092 3457 28120 3488
rect 43714 3476 43720 3528
rect 43772 3516 43778 3528
rect 44652 3516 44680 3547
rect 45097 3519 45155 3525
rect 45097 3516 45109 3519
rect 43772 3488 45109 3516
rect 43772 3476 43778 3488
rect 45097 3485 45109 3488
rect 45143 3485 45155 3519
rect 45097 3479 45155 3485
rect 45204 3488 47670 3516
rect 28077 3451 28135 3457
rect 28077 3417 28089 3451
rect 28123 3417 28135 3451
rect 36354 3448 36360 3460
rect 36315 3420 36360 3448
rect 28077 3411 28135 3417
rect 36354 3408 36360 3420
rect 36412 3408 36418 3460
rect 39390 3408 39396 3460
rect 39448 3448 39454 3460
rect 39577 3451 39635 3457
rect 39577 3448 39589 3451
rect 39448 3420 39589 3448
rect 39448 3408 39454 3420
rect 39577 3417 39589 3420
rect 39623 3417 39635 3451
rect 41874 3448 41880 3460
rect 41835 3420 41880 3448
rect 39577 3411 39635 3417
rect 41874 3408 41880 3420
rect 41932 3408 41938 3460
rect 43990 3408 43996 3460
rect 44048 3448 44054 3460
rect 45204 3448 45232 3488
rect 44048 3420 45232 3448
rect 47642 3448 47670 3488
rect 47854 3476 47860 3528
rect 47912 3516 47918 3528
rect 48056 3516 48084 3547
rect 57054 3544 57060 3596
rect 57112 3584 57118 3596
rect 57238 3584 57244 3596
rect 57112 3556 57244 3584
rect 57112 3544 57118 3556
rect 57238 3544 57244 3556
rect 57296 3544 57302 3596
rect 48593 3519 48651 3525
rect 48593 3516 48605 3519
rect 47912 3488 48605 3516
rect 47912 3476 47918 3488
rect 48593 3485 48605 3488
rect 48639 3485 48651 3519
rect 48593 3479 48651 3485
rect 55769 3519 55827 3525
rect 55769 3485 55781 3519
rect 55815 3516 55827 3519
rect 58066 3516 58072 3528
rect 55815 3488 58072 3516
rect 55815 3485 55827 3488
rect 55769 3479 55827 3485
rect 58066 3476 58072 3488
rect 58124 3476 58130 3528
rect 54202 3448 54208 3460
rect 47642 3420 54208 3448
rect 44048 3408 44054 3420
rect 54202 3408 54208 3420
rect 54260 3448 54266 3460
rect 54297 3451 54355 3457
rect 54297 3448 54309 3451
rect 54260 3420 54309 3448
rect 54260 3408 54266 3420
rect 54297 3417 54309 3420
rect 54343 3417 54355 3451
rect 57422 3448 57428 3460
rect 57383 3420 57428 3448
rect 54297 3411 54355 3417
rect 57422 3408 57428 3420
rect 57480 3408 57486 3460
rect 58161 3451 58219 3457
rect 58161 3417 58173 3451
rect 58207 3448 58219 3451
rect 58894 3448 58900 3460
rect 58207 3420 58900 3448
rect 58207 3417 58219 3420
rect 58161 3411 58219 3417
rect 58894 3408 58900 3420
rect 58952 3408 58958 3460
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 2225 3383 2283 3389
rect 2225 3349 2237 3383
rect 2271 3380 2283 3383
rect 2590 3380 2596 3392
rect 2271 3352 2596 3380
rect 2271 3349 2283 3352
rect 2225 3343 2283 3349
rect 2590 3340 2596 3352
rect 2648 3340 2654 3392
rect 3234 3340 3240 3392
rect 3292 3380 3298 3392
rect 3881 3383 3939 3389
rect 3881 3380 3893 3383
rect 3292 3352 3893 3380
rect 3292 3340 3298 3352
rect 3881 3349 3893 3352
rect 3927 3349 3939 3383
rect 3881 3343 3939 3349
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 6512 3352 6653 3380
rect 6512 3340 6518 3352
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 6641 3343 6699 3349
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10560 3352 10977 3380
rect 10560 3340 10566 3352
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 13262 3380 13268 3392
rect 13223 3352 13268 3380
rect 10965 3343 11023 3349
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 14366 3340 14372 3392
rect 14424 3380 14430 3392
rect 15105 3383 15163 3389
rect 15105 3380 15117 3383
rect 14424 3352 15117 3380
rect 14424 3340 14430 3352
rect 15105 3349 15117 3352
rect 15151 3349 15163 3383
rect 17494 3380 17500 3392
rect 17455 3352 17500 3380
rect 15105 3343 15163 3349
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 18598 3380 18604 3392
rect 18559 3352 18604 3380
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 19610 3380 19616 3392
rect 19571 3352 19616 3380
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 20257 3383 20315 3389
rect 20257 3349 20269 3383
rect 20303 3380 20315 3383
rect 20530 3380 20536 3392
rect 20303 3352 20536 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 20993 3383 21051 3389
rect 20993 3380 21005 3383
rect 20772 3352 21005 3380
rect 20772 3340 20778 3352
rect 20993 3349 21005 3352
rect 21039 3349 21051 3383
rect 22002 3380 22008 3392
rect 21963 3352 22008 3380
rect 20993 3343 21051 3349
rect 22002 3340 22008 3352
rect 22060 3340 22066 3392
rect 24302 3380 24308 3392
rect 24263 3352 24308 3380
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 28626 3380 28632 3392
rect 28587 3352 28632 3380
rect 28626 3340 28632 3352
rect 28684 3340 28690 3392
rect 29365 3383 29423 3389
rect 29365 3349 29377 3383
rect 29411 3380 29423 3383
rect 29730 3380 29736 3392
rect 29411 3352 29736 3380
rect 29411 3349 29423 3352
rect 29365 3343 29423 3349
rect 29730 3340 29736 3352
rect 29788 3340 29794 3392
rect 34241 3383 34299 3389
rect 34241 3349 34253 3383
rect 34287 3380 34299 3383
rect 34606 3380 34612 3392
rect 34287 3352 34612 3380
rect 34287 3349 34299 3352
rect 34241 3343 34299 3349
rect 34606 3340 34612 3352
rect 34664 3340 34670 3392
rect 36446 3340 36452 3392
rect 36504 3380 36510 3392
rect 37185 3383 37243 3389
rect 37185 3380 37197 3383
rect 36504 3352 37197 3380
rect 36504 3340 36510 3352
rect 37185 3349 37197 3352
rect 37231 3349 37243 3383
rect 37185 3343 37243 3349
rect 38197 3383 38255 3389
rect 38197 3349 38209 3383
rect 38243 3380 38255 3383
rect 38286 3380 38292 3392
rect 38243 3352 38292 3380
rect 38243 3349 38255 3352
rect 38197 3343 38255 3349
rect 38286 3340 38292 3352
rect 38344 3340 38350 3392
rect 40586 3340 40592 3392
rect 40644 3380 40650 3392
rect 41049 3383 41107 3389
rect 41049 3380 41061 3383
rect 40644 3352 41061 3380
rect 40644 3340 40650 3352
rect 41049 3349 41061 3352
rect 41095 3380 41107 3383
rect 41782 3380 41788 3392
rect 41095 3352 41788 3380
rect 41095 3349 41107 3352
rect 41049 3343 41107 3349
rect 41782 3340 41788 3352
rect 41840 3340 41846 3392
rect 42705 3383 42763 3389
rect 42705 3349 42717 3383
rect 42751 3380 42763 3383
rect 42794 3380 42800 3392
rect 42751 3352 42800 3380
rect 42751 3349 42763 3352
rect 42705 3343 42763 3349
rect 42794 3340 42800 3352
rect 42852 3340 42858 3392
rect 43162 3380 43168 3392
rect 43123 3352 43168 3380
rect 43162 3340 43168 3352
rect 43220 3340 43226 3392
rect 44082 3340 44088 3392
rect 44140 3380 44146 3392
rect 44453 3383 44511 3389
rect 44453 3380 44465 3383
rect 44140 3352 44465 3380
rect 44140 3340 44146 3352
rect 44453 3349 44465 3352
rect 44499 3349 44511 3383
rect 45830 3380 45836 3392
rect 45791 3352 45836 3380
rect 44453 3343 44511 3349
rect 45830 3340 45836 3352
rect 45888 3340 45894 3392
rect 46014 3340 46020 3392
rect 46072 3380 46078 3392
rect 46385 3383 46443 3389
rect 46385 3380 46397 3383
rect 46072 3352 46397 3380
rect 46072 3340 46078 3352
rect 46385 3349 46397 3352
rect 46431 3349 46443 3383
rect 46385 3343 46443 3349
rect 47026 3340 47032 3392
rect 47084 3380 47090 3392
rect 47305 3383 47363 3389
rect 47305 3380 47317 3383
rect 47084 3352 47317 3380
rect 47084 3340 47090 3352
rect 47305 3349 47317 3352
rect 47351 3349 47363 3383
rect 49602 3380 49608 3392
rect 49563 3352 49608 3380
rect 47305 3343 47363 3349
rect 49602 3340 49608 3352
rect 49660 3340 49666 3392
rect 50062 3380 50068 3392
rect 50023 3352 50068 3380
rect 50062 3340 50068 3352
rect 50120 3340 50126 3392
rect 52089 3383 52147 3389
rect 52089 3349 52101 3383
rect 52135 3380 52147 3383
rect 52362 3380 52368 3392
rect 52135 3352 52368 3380
rect 52135 3349 52147 3352
rect 52089 3343 52147 3349
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 52546 3380 52552 3392
rect 52507 3352 52552 3380
rect 52546 3340 52552 3352
rect 52604 3340 52610 3392
rect 53190 3380 53196 3392
rect 53151 3352 53196 3380
rect 53190 3340 53196 3352
rect 53248 3340 53254 3392
rect 53374 3340 53380 3392
rect 53432 3380 53438 3392
rect 53745 3383 53803 3389
rect 53745 3380 53757 3383
rect 53432 3352 53757 3380
rect 53432 3340 53438 3352
rect 53745 3349 53757 3352
rect 53791 3349 53803 3383
rect 53745 3343 53803 3349
rect 55217 3383 55275 3389
rect 55217 3349 55229 3383
rect 55263 3380 55275 3383
rect 55674 3380 55680 3392
rect 55263 3352 55680 3380
rect 55263 3349 55275 3352
rect 55217 3343 55275 3349
rect 55674 3340 55680 3352
rect 55732 3340 55738 3392
rect 56318 3380 56324 3392
rect 56279 3352 56324 3380
rect 56318 3340 56324 3352
rect 56376 3340 56382 3392
rect 1104 3290 58880 3312
rect 1104 3238 10614 3290
rect 10666 3238 10678 3290
rect 10730 3238 10742 3290
rect 10794 3238 10806 3290
rect 10858 3238 29878 3290
rect 29930 3238 29942 3290
rect 29994 3238 30006 3290
rect 30058 3238 30070 3290
rect 30122 3238 49142 3290
rect 49194 3238 49206 3290
rect 49258 3238 49270 3290
rect 49322 3238 49334 3290
rect 49386 3238 58880 3290
rect 1104 3216 58880 3238
rect 7006 3176 7012 3188
rect 6967 3148 7012 3176
rect 7006 3136 7012 3148
rect 7064 3136 7070 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 8757 3179 8815 3185
rect 8757 3176 8769 3179
rect 8720 3148 8769 3176
rect 8720 3136 8726 3148
rect 8757 3145 8769 3148
rect 8803 3145 8815 3179
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 8757 3139 8815 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 13722 3176 13728 3188
rect 13683 3148 13728 3176
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 15381 3179 15439 3185
rect 15381 3176 15393 3179
rect 14240 3148 15393 3176
rect 14240 3136 14246 3148
rect 15381 3145 15393 3148
rect 15427 3145 15439 3179
rect 15381 3139 15439 3145
rect 16758 3136 16764 3188
rect 16816 3176 16822 3188
rect 17034 3176 17040 3188
rect 16816 3148 17040 3176
rect 16816 3136 16822 3148
rect 17034 3136 17040 3148
rect 17092 3136 17098 3188
rect 19794 3176 19800 3188
rect 19755 3148 19800 3176
rect 19794 3136 19800 3148
rect 19852 3136 19858 3188
rect 27798 3176 27804 3188
rect 27759 3148 27804 3176
rect 27798 3136 27804 3148
rect 27856 3136 27862 3188
rect 29362 3136 29368 3188
rect 29420 3176 29426 3188
rect 47029 3179 47087 3185
rect 29420 3148 46980 3176
rect 29420 3136 29426 3148
rect 35066 3108 35072 3120
rect 4172 3080 35072 3108
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 1412 3012 3525 3040
rect 1412 2984 1440 3012
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 1394 2972 1400 2984
rect 1355 2944 1400 2972
rect 1394 2932 1400 2944
rect 1452 2932 1458 2984
rect 2133 2975 2191 2981
rect 2133 2941 2145 2975
rect 2179 2972 2191 2975
rect 2406 2972 2412 2984
rect 2179 2944 2412 2972
rect 2179 2941 2191 2944
rect 2133 2935 2191 2941
rect 2406 2932 2412 2944
rect 2464 2932 2470 2984
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3142 2972 3148 2984
rect 3007 2944 3148 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 3142 2932 3148 2944
rect 3200 2972 3206 2984
rect 4172 2972 4200 3080
rect 35066 3068 35072 3080
rect 35124 3068 35130 3120
rect 36538 3108 36544 3120
rect 35360 3080 36544 3108
rect 35360 3052 35388 3080
rect 36538 3068 36544 3080
rect 36596 3068 36602 3120
rect 37826 3068 37832 3120
rect 37884 3108 37890 3120
rect 38378 3108 38384 3120
rect 37884 3080 38384 3108
rect 37884 3068 37890 3080
rect 38378 3068 38384 3080
rect 38436 3068 38442 3120
rect 41598 3108 41604 3120
rect 39224 3080 41604 3108
rect 16206 3040 16212 3052
rect 4356 3012 16212 3040
rect 4356 2981 4384 3012
rect 16206 3000 16212 3012
rect 16264 3000 16270 3052
rect 19426 3040 19432 3052
rect 19076 3012 19432 3040
rect 3200 2944 4200 2972
rect 4341 2975 4399 2981
rect 3200 2932 3206 2944
rect 4341 2941 4353 2975
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 6454 2932 6460 2984
rect 6512 2972 6518 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6512 2944 6837 2972
rect 6512 2932 6518 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 8941 2975 8999 2981
rect 8941 2972 8953 2975
rect 8812 2944 8953 2972
rect 8812 2932 8818 2944
rect 8941 2941 8953 2944
rect 8987 2941 8999 2975
rect 8941 2935 8999 2941
rect 9674 2932 9680 2984
rect 9732 2972 9738 2984
rect 9861 2975 9919 2981
rect 9861 2972 9873 2975
rect 9732 2944 9873 2972
rect 9732 2932 9738 2944
rect 9861 2941 9873 2944
rect 9907 2972 9919 2975
rect 10321 2975 10379 2981
rect 10321 2972 10333 2975
rect 9907 2944 10333 2972
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 10321 2941 10333 2944
rect 10367 2941 10379 2975
rect 10321 2935 10379 2941
rect 11057 2975 11115 2981
rect 11057 2941 11069 2975
rect 11103 2972 11115 2975
rect 11514 2972 11520 2984
rect 11103 2944 11520 2972
rect 11103 2941 11115 2944
rect 11057 2935 11115 2941
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 13078 2972 13084 2984
rect 12991 2944 13084 2972
rect 13078 2932 13084 2944
rect 13136 2972 13142 2984
rect 13262 2972 13268 2984
rect 13136 2944 13268 2972
rect 13136 2932 13142 2944
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 15378 2972 15384 2984
rect 15339 2944 15384 2972
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15528 2944 15577 2972
rect 15528 2932 15534 2944
rect 15565 2941 15577 2944
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 16301 2975 16359 2981
rect 16301 2941 16313 2975
rect 16347 2972 16359 2975
rect 16850 2972 16856 2984
rect 16347 2944 16856 2972
rect 16347 2941 16359 2944
rect 16301 2935 16359 2941
rect 16850 2932 16856 2944
rect 16908 2932 16914 2984
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 19076 2981 19104 3012
rect 19426 3000 19432 3012
rect 19484 3000 19490 3052
rect 27614 3000 27620 3052
rect 27672 3040 27678 3052
rect 28353 3043 28411 3049
rect 28353 3040 28365 3043
rect 27672 3012 28365 3040
rect 27672 3000 27678 3012
rect 28353 3009 28365 3012
rect 28399 3009 28411 3043
rect 28353 3003 28411 3009
rect 29638 3000 29644 3052
rect 29696 3040 29702 3052
rect 29917 3043 29975 3049
rect 29917 3040 29929 3043
rect 29696 3012 29929 3040
rect 29696 3000 29702 3012
rect 29917 3009 29929 3012
rect 29963 3009 29975 3043
rect 29917 3003 29975 3009
rect 34701 3043 34759 3049
rect 34701 3009 34713 3043
rect 34747 3040 34759 3043
rect 35342 3040 35348 3052
rect 34747 3012 35348 3040
rect 34747 3009 34759 3012
rect 34701 3003 34759 3009
rect 35342 3000 35348 3012
rect 35400 3000 35406 3052
rect 36170 3040 36176 3052
rect 36131 3012 36176 3040
rect 36170 3000 36176 3012
rect 36228 3000 36234 3052
rect 39224 3040 39252 3080
rect 41598 3068 41604 3080
rect 41656 3068 41662 3120
rect 41693 3111 41751 3117
rect 41693 3077 41705 3111
rect 41739 3077 41751 3111
rect 42334 3108 42340 3120
rect 42295 3080 42340 3108
rect 41693 3071 41751 3077
rect 37660 3012 39252 3040
rect 39301 3043 39359 3049
rect 37660 2984 37688 3012
rect 39301 3009 39313 3043
rect 39347 3040 39359 3043
rect 40034 3040 40040 3052
rect 39347 3012 40040 3040
rect 39347 3009 39359 3012
rect 39301 3003 39359 3009
rect 40034 3000 40040 3012
rect 40092 3000 40098 3052
rect 41046 3040 41052 3052
rect 41007 3012 41052 3040
rect 41046 3000 41052 3012
rect 41104 3000 41110 3052
rect 41230 3040 41236 3052
rect 41191 3012 41236 3040
rect 41230 3000 41236 3012
rect 41288 3000 41294 3052
rect 41506 3040 41512 3052
rect 41340 3012 41512 3040
rect 17957 2975 18015 2981
rect 17957 2972 17969 2975
rect 17552 2944 17969 2972
rect 17552 2932 17558 2944
rect 17957 2941 17969 2944
rect 18003 2941 18015 2975
rect 17957 2935 18015 2941
rect 19061 2975 19119 2981
rect 19061 2941 19073 2975
rect 19107 2941 19119 2975
rect 19061 2935 19119 2941
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 19610 2972 19616 2984
rect 19392 2944 19616 2972
rect 19392 2932 19398 2944
rect 19610 2932 19616 2944
rect 19668 2932 19674 2984
rect 20714 2972 20720 2984
rect 20675 2944 20720 2972
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 22094 2932 22100 2984
rect 22152 2972 22158 2984
rect 22741 2975 22799 2981
rect 22741 2972 22753 2975
rect 22152 2944 22753 2972
rect 22152 2932 22158 2944
rect 22741 2941 22753 2944
rect 22787 2941 22799 2975
rect 22741 2935 22799 2941
rect 23661 2975 23719 2981
rect 23661 2941 23673 2975
rect 23707 2941 23719 2975
rect 23661 2935 23719 2941
rect 2314 2904 2320 2916
rect 2275 2876 2320 2904
rect 2314 2864 2320 2876
rect 2372 2864 2378 2916
rect 2774 2904 2780 2916
rect 2735 2876 2780 2904
rect 2774 2864 2780 2876
rect 2832 2864 2838 2916
rect 4154 2904 4160 2916
rect 3436 2876 4016 2904
rect 4115 2876 4160 2904
rect 1581 2839 1639 2845
rect 1581 2805 1593 2839
rect 1627 2836 1639 2839
rect 3436 2836 3464 2876
rect 1627 2808 3464 2836
rect 3988 2836 4016 2876
rect 4154 2864 4160 2876
rect 4212 2864 4218 2916
rect 4614 2864 4620 2916
rect 4672 2904 4678 2916
rect 4893 2907 4951 2913
rect 4893 2904 4905 2907
rect 4672 2876 4905 2904
rect 4672 2864 4678 2876
rect 4893 2873 4905 2876
rect 4939 2873 4951 2907
rect 4893 2867 4951 2873
rect 5077 2907 5135 2913
rect 5077 2873 5089 2907
rect 5123 2904 5135 2907
rect 5718 2904 5724 2916
rect 5123 2876 5724 2904
rect 5123 2873 5135 2876
rect 5077 2867 5135 2873
rect 5718 2864 5724 2876
rect 5776 2864 5782 2916
rect 12158 2904 12164 2916
rect 6426 2876 12164 2904
rect 6426 2836 6454 2876
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 12894 2904 12900 2916
rect 12855 2876 12900 2904
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 14274 2904 14280 2916
rect 14235 2876 14280 2904
rect 14274 2864 14280 2876
rect 14332 2864 14338 2916
rect 14458 2904 14464 2916
rect 14419 2876 14464 2904
rect 14458 2864 14464 2876
rect 14516 2864 14522 2916
rect 16114 2904 16120 2916
rect 16075 2876 16120 2904
rect 16114 2864 16120 2876
rect 16172 2864 16178 2916
rect 23676 2904 23704 2935
rect 24302 2932 24308 2984
rect 24360 2972 24366 2984
rect 24397 2975 24455 2981
rect 24397 2972 24409 2975
rect 24360 2944 24409 2972
rect 24360 2932 24366 2944
rect 24397 2941 24409 2944
rect 24443 2941 24455 2975
rect 25130 2972 25136 2984
rect 25091 2944 25136 2972
rect 24397 2935 24455 2941
rect 25130 2932 25136 2944
rect 25188 2932 25194 2984
rect 25958 2972 25964 2984
rect 25919 2944 25964 2972
rect 25958 2932 25964 2944
rect 26016 2932 26022 2984
rect 26234 2932 26240 2984
rect 26292 2972 26298 2984
rect 26697 2975 26755 2981
rect 26697 2972 26709 2975
rect 26292 2944 26709 2972
rect 26292 2932 26298 2944
rect 26697 2941 26709 2944
rect 26743 2941 26755 2975
rect 26697 2935 26755 2941
rect 26970 2932 26976 2984
rect 27028 2972 27034 2984
rect 28169 2975 28227 2981
rect 28169 2972 28181 2975
rect 27028 2944 28181 2972
rect 27028 2932 27034 2944
rect 28169 2941 28181 2944
rect 28215 2941 28227 2975
rect 28169 2935 28227 2941
rect 28261 2975 28319 2981
rect 28261 2941 28273 2975
rect 28307 2972 28319 2975
rect 28810 2972 28816 2984
rect 28307 2944 28816 2972
rect 28307 2941 28319 2944
rect 28261 2935 28319 2941
rect 28810 2932 28816 2944
rect 28868 2932 28874 2984
rect 28902 2932 28908 2984
rect 28960 2972 28966 2984
rect 29181 2975 29239 2981
rect 29181 2972 29193 2975
rect 28960 2944 29193 2972
rect 28960 2932 28966 2944
rect 29181 2941 29193 2944
rect 29227 2941 29239 2975
rect 29181 2935 29239 2941
rect 29730 2932 29736 2984
rect 29788 2972 29794 2984
rect 29825 2975 29883 2981
rect 29825 2972 29837 2975
rect 29788 2944 29837 2972
rect 29788 2932 29794 2944
rect 29825 2941 29837 2944
rect 29871 2941 29883 2975
rect 29825 2935 29883 2941
rect 31113 2975 31171 2981
rect 31113 2941 31125 2975
rect 31159 2972 31171 2975
rect 31202 2972 31208 2984
rect 31159 2944 31208 2972
rect 31159 2941 31171 2944
rect 31113 2935 31171 2941
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 31938 2972 31944 2984
rect 31899 2944 31944 2972
rect 31938 2932 31944 2944
rect 31996 2932 32002 2984
rect 33137 2975 33195 2981
rect 33137 2941 33149 2975
rect 33183 2972 33195 2975
rect 33594 2972 33600 2984
rect 33183 2944 33600 2972
rect 33183 2941 33195 2944
rect 33137 2935 33195 2941
rect 33594 2932 33600 2944
rect 33652 2932 33658 2984
rect 34606 2972 34612 2984
rect 34567 2944 34612 2972
rect 34606 2932 34612 2944
rect 34664 2932 34670 2984
rect 36446 2972 36452 2984
rect 36407 2944 36452 2972
rect 36446 2932 36452 2944
rect 36504 2932 36510 2984
rect 37093 2975 37151 2981
rect 37093 2941 37105 2975
rect 37139 2972 37151 2975
rect 37642 2972 37648 2984
rect 37139 2944 37648 2972
rect 37139 2941 37151 2944
rect 37093 2935 37151 2941
rect 37642 2932 37648 2944
rect 37700 2932 37706 2984
rect 38286 2972 38292 2984
rect 38247 2944 38292 2972
rect 38286 2932 38292 2944
rect 38344 2932 38350 2984
rect 39482 2932 39488 2984
rect 39540 2972 39546 2984
rect 39945 2975 40003 2981
rect 39945 2972 39957 2975
rect 39540 2944 39957 2972
rect 39540 2932 39546 2944
rect 39945 2941 39957 2944
rect 39991 2972 40003 2975
rect 40313 2975 40371 2981
rect 39991 2944 40264 2972
rect 39991 2941 40003 2944
rect 39945 2935 40003 2941
rect 20916 2876 23704 2904
rect 24581 2907 24639 2913
rect 3988 2808 6454 2836
rect 1627 2805 1639 2808
rect 1581 2799 1639 2805
rect 7374 2796 7380 2848
rect 7432 2836 7438 2848
rect 7745 2839 7803 2845
rect 7745 2836 7757 2839
rect 7432 2808 7757 2836
rect 7432 2796 7438 2808
rect 7745 2805 7757 2808
rect 7791 2805 7803 2839
rect 10962 2836 10968 2848
rect 10923 2808 10968 2836
rect 7745 2799 7803 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 12069 2839 12127 2845
rect 12069 2836 12081 2839
rect 12032 2808 12081 2836
rect 12032 2796 12038 2808
rect 12069 2805 12081 2808
rect 12115 2805 12127 2839
rect 19058 2836 19064 2848
rect 19019 2808 19064 2836
rect 12069 2799 12127 2805
rect 19058 2796 19064 2808
rect 19116 2796 19122 2848
rect 20916 2845 20944 2876
rect 24581 2873 24593 2907
rect 24627 2904 24639 2907
rect 24854 2904 24860 2916
rect 24627 2876 24860 2904
rect 24627 2873 24639 2876
rect 24581 2867 24639 2873
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 25314 2904 25320 2916
rect 25275 2876 25320 2904
rect 25314 2864 25320 2876
rect 25372 2864 25378 2916
rect 25774 2904 25780 2916
rect 25735 2876 25780 2904
rect 25774 2864 25780 2876
rect 25832 2864 25838 2916
rect 30374 2864 30380 2916
rect 30432 2904 30438 2916
rect 30929 2907 30987 2913
rect 30929 2904 30941 2907
rect 30432 2876 30941 2904
rect 30432 2864 30438 2876
rect 30929 2873 30941 2876
rect 30975 2873 30987 2907
rect 31754 2904 31760 2916
rect 31715 2876 31760 2904
rect 30929 2867 30987 2873
rect 31754 2864 31760 2876
rect 31812 2864 31818 2916
rect 34698 2864 34704 2916
rect 34756 2904 34762 2916
rect 35253 2907 35311 2913
rect 35253 2904 35265 2907
rect 34756 2876 35265 2904
rect 34756 2864 34762 2876
rect 35253 2873 35265 2876
rect 35299 2904 35311 2907
rect 36262 2904 36268 2916
rect 35299 2876 36268 2904
rect 35299 2873 35311 2876
rect 35253 2867 35311 2873
rect 36262 2864 36268 2876
rect 36320 2864 36326 2916
rect 39117 2907 39175 2913
rect 39117 2873 39129 2907
rect 39163 2904 39175 2907
rect 40126 2904 40132 2916
rect 39163 2876 40132 2904
rect 39163 2873 39175 2876
rect 39117 2867 39175 2873
rect 40126 2864 40132 2876
rect 40184 2864 40190 2916
rect 20901 2839 20959 2845
rect 20901 2805 20913 2839
rect 20947 2805 20959 2839
rect 20901 2799 20959 2805
rect 21637 2839 21695 2845
rect 21637 2805 21649 2839
rect 21683 2836 21695 2839
rect 22094 2836 22100 2848
rect 21683 2808 22100 2836
rect 21683 2805 21695 2808
rect 21637 2799 21695 2805
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 22554 2836 22560 2848
rect 22515 2808 22560 2836
rect 22554 2796 22560 2808
rect 22612 2796 22618 2848
rect 23753 2839 23811 2845
rect 23753 2805 23765 2839
rect 23799 2836 23811 2839
rect 25866 2836 25872 2848
rect 23799 2808 25872 2836
rect 23799 2805 23811 2808
rect 23753 2799 23811 2805
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 26786 2836 26792 2848
rect 26747 2808 26792 2836
rect 26786 2796 26792 2808
rect 26844 2796 26850 2848
rect 33778 2836 33784 2848
rect 33739 2808 33784 2836
rect 33778 2796 33784 2808
rect 33836 2796 33842 2848
rect 39942 2796 39948 2848
rect 40000 2836 40006 2848
rect 40037 2839 40095 2845
rect 40037 2836 40049 2839
rect 40000 2808 40049 2836
rect 40000 2796 40006 2808
rect 40037 2805 40049 2808
rect 40083 2805 40095 2839
rect 40236 2836 40264 2944
rect 40313 2941 40325 2975
rect 40359 2972 40371 2975
rect 40586 2972 40592 2984
rect 40359 2944 40592 2972
rect 40359 2941 40371 2944
rect 40313 2935 40371 2941
rect 40586 2932 40592 2944
rect 40644 2932 40650 2984
rect 41340 2981 41368 3012
rect 41506 3000 41512 3012
rect 41564 3000 41570 3052
rect 41708 3040 41736 3071
rect 42334 3068 42340 3080
rect 42392 3068 42398 3120
rect 43622 3108 43628 3120
rect 43583 3080 43628 3108
rect 43622 3068 43628 3080
rect 43680 3068 43686 3120
rect 45462 3108 45468 3120
rect 45423 3080 45468 3108
rect 45462 3068 45468 3080
rect 45520 3068 45526 3120
rect 46952 3108 46980 3148
rect 47029 3145 47041 3179
rect 47075 3176 47087 3179
rect 47118 3176 47124 3188
rect 47075 3148 47124 3176
rect 47075 3145 47087 3148
rect 47029 3139 47087 3145
rect 47118 3136 47124 3148
rect 47176 3136 47182 3188
rect 53098 3176 53104 3188
rect 47642 3148 52960 3176
rect 53059 3148 53104 3176
rect 47642 3108 47670 3148
rect 49694 3108 49700 3120
rect 46952 3080 47670 3108
rect 49655 3080 49700 3108
rect 49694 3068 49700 3080
rect 49752 3068 49758 3120
rect 50798 3068 50804 3120
rect 50856 3108 50862 3120
rect 52932 3108 52960 3148
rect 53098 3136 53104 3148
rect 53156 3136 53162 3188
rect 56410 3176 56416 3188
rect 55876 3148 56416 3176
rect 55582 3108 55588 3120
rect 50856 3080 52868 3108
rect 52932 3080 55588 3108
rect 50856 3068 50862 3080
rect 44082 3040 44088 3052
rect 41708 3012 42518 3040
rect 44043 3012 44088 3040
rect 41325 2975 41383 2981
rect 41325 2941 41337 2975
rect 41371 2941 41383 2975
rect 42490 2972 42518 3012
rect 44082 3000 44088 3012
rect 44140 3000 44146 3052
rect 52840 3040 52868 3080
rect 55582 3068 55588 3080
rect 55640 3068 55646 3120
rect 55876 3040 55904 3148
rect 56410 3136 56416 3148
rect 56468 3176 56474 3188
rect 56468 3148 56686 3176
rect 56468 3136 56474 3148
rect 55953 3111 56011 3117
rect 55953 3077 55965 3111
rect 55999 3077 56011 3111
rect 56658 3108 56686 3148
rect 57146 3136 57152 3188
rect 57204 3176 57210 3188
rect 57241 3179 57299 3185
rect 57241 3176 57253 3179
rect 57204 3148 57253 3176
rect 57204 3136 57210 3148
rect 57241 3145 57253 3148
rect 57287 3145 57299 3179
rect 57241 3139 57299 3145
rect 56658 3080 57836 3108
rect 55953 3071 56011 3077
rect 44192 3012 51764 3040
rect 52840 3012 55904 3040
rect 55968 3040 55996 3071
rect 57808 3049 57836 3080
rect 57793 3043 57851 3049
rect 55968 3012 57744 3040
rect 44192 2972 44220 3012
rect 42490 2944 44220 2972
rect 41325 2935 41383 2941
rect 45094 2932 45100 2984
rect 45152 2972 45158 2984
rect 45649 2975 45707 2981
rect 45649 2972 45661 2975
rect 45152 2944 45661 2972
rect 45152 2932 45158 2944
rect 45649 2941 45661 2944
rect 45695 2972 45707 2975
rect 45830 2972 45836 2984
rect 45695 2944 45836 2972
rect 45695 2941 45707 2944
rect 45649 2935 45707 2941
rect 45830 2932 45836 2944
rect 45888 2932 45894 2984
rect 46293 2975 46351 2981
rect 46293 2941 46305 2975
rect 46339 2972 46351 2975
rect 46934 2972 46940 2984
rect 46339 2944 46940 2972
rect 46339 2941 46351 2944
rect 46293 2935 46351 2941
rect 46934 2932 46940 2944
rect 46992 2932 46998 2984
rect 47026 2932 47032 2984
rect 47084 2972 47090 2984
rect 47121 2975 47179 2981
rect 47121 2972 47133 2975
rect 47084 2944 47133 2972
rect 47084 2932 47090 2944
rect 47121 2941 47133 2944
rect 47167 2941 47179 2975
rect 47121 2935 47179 2941
rect 47578 2932 47584 2984
rect 47636 2972 47642 2984
rect 47673 2975 47731 2981
rect 47673 2972 47685 2975
rect 47636 2944 47685 2972
rect 47636 2932 47642 2944
rect 47673 2941 47685 2944
rect 47719 2941 47731 2975
rect 47673 2935 47731 2941
rect 47857 2975 47915 2981
rect 47857 2941 47869 2975
rect 47903 2972 47915 2975
rect 47903 2944 49648 2972
rect 47903 2941 47915 2944
rect 47857 2935 47915 2941
rect 41230 2864 41236 2916
rect 41288 2904 41294 2916
rect 42058 2904 42064 2916
rect 41288 2876 42064 2904
rect 41288 2864 41294 2876
rect 42058 2864 42064 2876
rect 42116 2864 42122 2916
rect 42521 2907 42579 2913
rect 42521 2873 42533 2907
rect 42567 2904 42579 2907
rect 42794 2904 42800 2916
rect 42567 2876 42800 2904
rect 42567 2873 42579 2876
rect 42521 2867 42579 2873
rect 42794 2864 42800 2876
rect 42852 2864 42858 2916
rect 44174 2904 44180 2916
rect 44135 2876 44180 2904
rect 44174 2864 44180 2876
rect 44232 2864 44238 2916
rect 44634 2864 44640 2916
rect 44692 2904 44698 2916
rect 44729 2907 44787 2913
rect 44729 2904 44741 2907
rect 44692 2876 44741 2904
rect 44692 2864 44698 2876
rect 44729 2873 44741 2876
rect 44775 2873 44787 2907
rect 44910 2904 44916 2916
rect 44871 2876 44916 2904
rect 44729 2867 44787 2873
rect 44910 2864 44916 2876
rect 44968 2864 44974 2916
rect 46474 2904 46480 2916
rect 46435 2876 46480 2904
rect 46474 2864 46480 2876
rect 46532 2864 46538 2916
rect 43990 2836 43996 2848
rect 40236 2808 43996 2836
rect 40037 2799 40095 2805
rect 43990 2796 43996 2808
rect 44048 2796 44054 2848
rect 44085 2839 44143 2845
rect 44085 2805 44097 2839
rect 44131 2836 44143 2839
rect 44266 2836 44272 2848
rect 44131 2808 44272 2836
rect 44131 2805 44143 2808
rect 44085 2799 44143 2805
rect 44266 2796 44272 2808
rect 44324 2796 44330 2848
rect 44358 2796 44364 2848
rect 44416 2836 44422 2848
rect 47596 2836 47624 2932
rect 48314 2864 48320 2916
rect 48372 2904 48378 2916
rect 48777 2907 48835 2913
rect 48777 2904 48789 2907
rect 48372 2876 48789 2904
rect 48372 2864 48378 2876
rect 48777 2873 48789 2876
rect 48823 2873 48835 2907
rect 48777 2867 48835 2873
rect 48961 2907 49019 2913
rect 48961 2873 48973 2907
rect 49007 2873 49019 2907
rect 48961 2867 49019 2873
rect 44416 2808 47624 2836
rect 47765 2839 47823 2845
rect 44416 2796 44422 2808
rect 47765 2805 47777 2839
rect 47811 2836 47823 2839
rect 48976 2836 49004 2867
rect 47811 2808 49004 2836
rect 49620 2836 49648 2944
rect 49694 2932 49700 2984
rect 49752 2972 49758 2984
rect 49881 2975 49939 2981
rect 49881 2972 49893 2975
rect 49752 2944 49893 2972
rect 49752 2932 49758 2944
rect 49881 2941 49893 2944
rect 49927 2972 49939 2975
rect 50062 2972 50068 2984
rect 49927 2944 50068 2972
rect 49927 2941 49939 2944
rect 49881 2935 49939 2941
rect 50062 2932 50068 2944
rect 50120 2932 50126 2984
rect 51736 2981 51764 3012
rect 51721 2975 51779 2981
rect 51721 2941 51733 2975
rect 51767 2941 51779 2975
rect 51721 2935 51779 2941
rect 52457 2975 52515 2981
rect 52457 2941 52469 2975
rect 52503 2972 52515 2975
rect 52546 2972 52552 2984
rect 52503 2944 52552 2972
rect 52503 2941 52515 2944
rect 52457 2935 52515 2941
rect 52546 2932 52552 2944
rect 52604 2932 52610 2984
rect 52914 2972 52920 2984
rect 52827 2944 52920 2972
rect 52914 2932 52920 2944
rect 52972 2972 52978 2984
rect 53190 2972 53196 2984
rect 52972 2944 53196 2972
rect 52972 2932 52978 2944
rect 53190 2932 53196 2944
rect 53248 2932 53254 2984
rect 54018 2972 54024 2984
rect 53931 2944 54024 2972
rect 54018 2932 54024 2944
rect 54076 2932 54082 2984
rect 54202 2972 54208 2984
rect 54163 2944 54208 2972
rect 54202 2932 54208 2944
rect 54260 2932 54266 2984
rect 54938 2972 54944 2984
rect 54899 2944 54944 2972
rect 54938 2932 54944 2944
rect 54996 2932 55002 2984
rect 55769 2975 55827 2981
rect 55769 2941 55781 2975
rect 55815 2972 55827 2975
rect 56318 2972 56324 2984
rect 55815 2944 56324 2972
rect 55815 2941 55827 2944
rect 55769 2935 55827 2941
rect 56318 2932 56324 2944
rect 56376 2932 56382 2984
rect 57514 2972 57520 2984
rect 57475 2944 57520 2972
rect 57514 2932 57520 2944
rect 57572 2932 57578 2984
rect 50154 2864 50160 2916
rect 50212 2904 50218 2916
rect 50433 2907 50491 2913
rect 50433 2904 50445 2907
rect 50212 2876 50445 2904
rect 50212 2864 50218 2876
rect 50433 2873 50445 2876
rect 50479 2873 50491 2907
rect 50614 2904 50620 2916
rect 50575 2876 50620 2904
rect 50433 2867 50491 2873
rect 50614 2864 50620 2876
rect 50672 2864 50678 2916
rect 51534 2904 51540 2916
rect 51495 2876 51540 2904
rect 51534 2864 51540 2876
rect 51592 2864 51598 2916
rect 54036 2904 54064 2932
rect 54754 2904 54760 2916
rect 52012 2876 54064 2904
rect 54715 2876 54760 2904
rect 52012 2836 52040 2876
rect 54754 2864 54760 2876
rect 54812 2864 54818 2916
rect 56502 2904 56508 2916
rect 56463 2876 56508 2904
rect 56502 2864 56508 2876
rect 56560 2864 56566 2916
rect 57716 2913 57744 3012
rect 57793 3009 57805 3043
rect 57839 3009 57851 3043
rect 57793 3003 57851 3009
rect 57701 2907 57759 2913
rect 57701 2873 57713 2907
rect 57747 2873 57759 2907
rect 57701 2867 57759 2873
rect 52270 2836 52276 2848
rect 49620 2808 52040 2836
rect 52231 2808 52276 2836
rect 47811 2805 47823 2808
rect 47765 2799 47823 2805
rect 52270 2796 52276 2808
rect 52328 2796 52334 2848
rect 54110 2836 54116 2848
rect 54071 2808 54116 2836
rect 54110 2796 54116 2808
rect 54168 2796 54174 2848
rect 56594 2836 56600 2848
rect 56555 2808 56600 2836
rect 56594 2796 56600 2808
rect 56652 2796 56658 2848
rect 1104 2746 58880 2768
rect 1104 2694 20246 2746
rect 20298 2694 20310 2746
rect 20362 2694 20374 2746
rect 20426 2694 20438 2746
rect 20490 2694 39510 2746
rect 39562 2694 39574 2746
rect 39626 2694 39638 2746
rect 39690 2694 39702 2746
rect 39754 2694 58880 2746
rect 1104 2672 58880 2694
rect 8754 2592 8760 2644
rect 8812 2632 8818 2644
rect 12434 2632 12440 2644
rect 8812 2604 9260 2632
rect 8812 2592 8818 2604
rect 1670 2564 1676 2576
rect 1631 2536 1676 2564
rect 1670 2524 1676 2536
rect 1728 2524 1734 2576
rect 8294 2564 8300 2576
rect 8255 2536 8300 2564
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 9232 2573 9260 2604
rect 10428 2604 12440 2632
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2533 9275 2567
rect 9217 2527 9275 2533
rect 9953 2567 10011 2573
rect 9953 2533 9965 2567
rect 9999 2564 10011 2567
rect 10318 2564 10324 2576
rect 9999 2536 10324 2564
rect 9999 2533 10011 2536
rect 9953 2527 10011 2533
rect 10318 2524 10324 2536
rect 10376 2524 10382 2576
rect 934 2456 940 2508
rect 992 2496 998 2508
rect 2041 2499 2099 2505
rect 2041 2496 2053 2499
rect 992 2468 2053 2496
rect 992 2456 998 2468
rect 2041 2465 2053 2468
rect 2087 2465 2099 2499
rect 2041 2459 2099 2465
rect 3145 2499 3203 2505
rect 3145 2465 3157 2499
rect 3191 2496 3203 2499
rect 3234 2496 3240 2508
rect 3191 2468 3240 2496
rect 3191 2465 3203 2468
rect 3145 2459 3203 2465
rect 2056 2428 2084 2459
rect 3234 2456 3240 2468
rect 3292 2456 3298 2508
rect 4893 2499 4951 2505
rect 4893 2465 4905 2499
rect 4939 2465 4951 2499
rect 4893 2459 4951 2465
rect 3881 2431 3939 2437
rect 3881 2428 3893 2431
rect 2056 2400 3893 2428
rect 3881 2397 3893 2400
rect 3927 2397 3939 2431
rect 4908 2428 4936 2459
rect 5534 2456 5540 2508
rect 5592 2496 5598 2508
rect 5629 2499 5687 2505
rect 5629 2496 5641 2499
rect 5592 2468 5641 2496
rect 5592 2456 5598 2468
rect 5629 2465 5641 2468
rect 5675 2496 5687 2499
rect 6549 2499 6607 2505
rect 6549 2496 6561 2499
rect 5675 2468 6561 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 6549 2465 6561 2468
rect 6595 2465 6607 2499
rect 6549 2459 6607 2465
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 7432 2468 7481 2496
rect 7432 2456 7438 2468
rect 7469 2465 7481 2468
rect 7515 2465 7527 2499
rect 7469 2459 7527 2465
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 10428 2496 10456 2604
rect 12434 2592 12440 2604
rect 12492 2592 12498 2644
rect 14366 2632 14372 2644
rect 13648 2604 14372 2632
rect 13648 2564 13676 2604
rect 14366 2592 14372 2604
rect 14424 2592 14430 2644
rect 14458 2592 14464 2644
rect 14516 2632 14522 2644
rect 14921 2635 14979 2641
rect 14921 2632 14933 2635
rect 14516 2604 14933 2632
rect 14516 2592 14522 2604
rect 14921 2601 14933 2604
rect 14967 2601 14979 2635
rect 15286 2632 15292 2644
rect 15247 2604 15292 2632
rect 14921 2595 14979 2601
rect 15286 2592 15292 2604
rect 15344 2592 15350 2644
rect 22002 2632 22008 2644
rect 21836 2604 22008 2632
rect 13814 2564 13820 2576
rect 10796 2536 13676 2564
rect 13775 2536 13820 2564
rect 10183 2468 10456 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 10689 2499 10747 2505
rect 10689 2496 10701 2499
rect 10560 2468 10701 2496
rect 10560 2456 10566 2468
rect 10689 2465 10701 2468
rect 10735 2465 10747 2499
rect 10689 2459 10747 2465
rect 10796 2428 10824 2536
rect 13814 2524 13820 2536
rect 13872 2524 13878 2576
rect 15381 2567 15439 2573
rect 15381 2533 15393 2567
rect 15427 2564 15439 2567
rect 16022 2564 16028 2576
rect 15427 2536 16028 2564
rect 15427 2533 15439 2536
rect 15381 2527 15439 2533
rect 16022 2524 16028 2536
rect 16080 2524 16086 2576
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 16301 2567 16359 2573
rect 16301 2564 16313 2567
rect 16264 2536 16313 2564
rect 16264 2524 16270 2536
rect 16301 2533 16313 2536
rect 16347 2533 16359 2567
rect 17494 2564 17500 2576
rect 16301 2527 16359 2533
rect 16500 2536 17500 2564
rect 11974 2456 11980 2508
rect 12032 2496 12038 2508
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 12032 2468 12357 2496
rect 12032 2456 12038 2468
rect 12345 2465 12357 2468
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 14182 2496 14188 2508
rect 13127 2468 14188 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 14182 2456 14188 2468
rect 14240 2456 14246 2508
rect 16500 2505 16528 2536
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 18138 2564 18144 2576
rect 18099 2536 18144 2564
rect 18138 2524 18144 2536
rect 18196 2524 18202 2576
rect 19061 2567 19119 2573
rect 19061 2533 19073 2567
rect 19107 2564 19119 2567
rect 19886 2564 19892 2576
rect 19107 2536 19892 2564
rect 19107 2533 19119 2536
rect 19061 2527 19119 2533
rect 19886 2524 19892 2536
rect 19944 2524 19950 2576
rect 20441 2567 20499 2573
rect 20441 2533 20453 2567
rect 20487 2564 20499 2567
rect 20622 2564 20628 2576
rect 20487 2536 20628 2564
rect 20487 2533 20499 2536
rect 20441 2527 20499 2533
rect 20622 2524 20628 2536
rect 20680 2524 20686 2576
rect 21836 2573 21864 2604
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 23474 2592 23480 2644
rect 23532 2632 23538 2644
rect 29362 2632 29368 2644
rect 23532 2604 24486 2632
rect 29323 2604 29368 2632
rect 23532 2592 23538 2604
rect 21821 2567 21879 2573
rect 21821 2533 21833 2567
rect 21867 2533 21879 2567
rect 21821 2527 21879 2533
rect 21910 2524 21916 2576
rect 21968 2564 21974 2576
rect 23109 2567 23167 2573
rect 23109 2564 23121 2567
rect 21968 2536 23121 2564
rect 21968 2524 21974 2536
rect 23109 2533 23121 2536
rect 23155 2533 23167 2567
rect 24458 2564 24486 2604
rect 29362 2592 29368 2604
rect 29420 2592 29426 2644
rect 33134 2592 33140 2644
rect 33192 2632 33198 2644
rect 33689 2635 33747 2641
rect 33689 2632 33701 2635
rect 33192 2604 33701 2632
rect 33192 2592 33198 2604
rect 33689 2601 33701 2604
rect 33735 2601 33747 2635
rect 35066 2632 35072 2644
rect 35027 2604 35072 2632
rect 33689 2595 33747 2601
rect 35066 2592 35072 2604
rect 35124 2592 35130 2644
rect 37366 2632 37372 2644
rect 37327 2604 37372 2632
rect 37366 2592 37372 2604
rect 37424 2592 37430 2644
rect 39945 2635 40003 2641
rect 39945 2601 39957 2635
rect 39991 2632 40003 2635
rect 40126 2632 40132 2644
rect 39991 2604 40132 2632
rect 39991 2601 40003 2604
rect 39945 2595 40003 2601
rect 40126 2592 40132 2604
rect 40184 2592 40190 2644
rect 41598 2592 41604 2644
rect 41656 2632 41662 2644
rect 43070 2632 43076 2644
rect 41656 2604 43076 2632
rect 41656 2592 41662 2604
rect 43070 2592 43076 2604
rect 43128 2592 43134 2644
rect 43162 2592 43168 2644
rect 43220 2632 43226 2644
rect 43220 2604 43265 2632
rect 43220 2592 43226 2604
rect 43346 2592 43352 2644
rect 43404 2632 43410 2644
rect 43993 2635 44051 2641
rect 43993 2632 44005 2635
rect 43404 2604 44005 2632
rect 43404 2592 43410 2604
rect 43993 2601 44005 2604
rect 44039 2632 44051 2635
rect 44358 2632 44364 2644
rect 44039 2604 44364 2632
rect 44039 2601 44051 2604
rect 43993 2595 44051 2601
rect 44358 2592 44364 2604
rect 44416 2592 44422 2644
rect 44545 2635 44603 2641
rect 44545 2601 44557 2635
rect 44591 2632 44603 2635
rect 44910 2632 44916 2644
rect 44591 2604 44916 2632
rect 44591 2601 44603 2604
rect 44545 2595 44603 2601
rect 44910 2592 44916 2604
rect 44968 2592 44974 2644
rect 46934 2632 46940 2644
rect 46895 2604 46940 2632
rect 46934 2592 46940 2604
rect 46992 2592 46998 2644
rect 49602 2592 49608 2644
rect 49660 2632 49666 2644
rect 50798 2632 50804 2644
rect 49660 2604 50804 2632
rect 49660 2592 49666 2604
rect 50798 2592 50804 2604
rect 50856 2592 50862 2644
rect 51074 2592 51080 2644
rect 51132 2632 51138 2644
rect 52365 2635 52423 2641
rect 52365 2632 52377 2635
rect 51132 2604 52377 2632
rect 51132 2592 51138 2604
rect 52365 2601 52377 2604
rect 52411 2601 52423 2635
rect 52365 2595 52423 2601
rect 26973 2567 27031 2573
rect 26973 2564 26985 2567
rect 24458 2536 26985 2564
rect 23109 2527 23167 2533
rect 26973 2533 26985 2536
rect 27019 2533 27031 2567
rect 26973 2527 27031 2533
rect 27157 2567 27215 2573
rect 27157 2533 27169 2567
rect 27203 2564 27215 2567
rect 27430 2564 27436 2576
rect 27203 2536 27436 2564
rect 27203 2533 27215 2536
rect 27157 2527 27215 2533
rect 27430 2524 27436 2536
rect 27488 2524 27494 2576
rect 28534 2524 28540 2576
rect 28592 2564 28598 2576
rect 28629 2567 28687 2573
rect 28629 2564 28641 2567
rect 28592 2536 28641 2564
rect 28592 2524 28598 2536
rect 28629 2533 28641 2536
rect 28675 2533 28687 2567
rect 30561 2567 30619 2573
rect 30561 2564 30573 2567
rect 28629 2527 28687 2533
rect 29288 2536 30573 2564
rect 16485 2499 16543 2505
rect 16485 2465 16497 2499
rect 16531 2465 16543 2499
rect 16666 2496 16672 2508
rect 16627 2468 16672 2496
rect 16485 2459 16543 2465
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 20530 2496 20536 2508
rect 18156 2468 20536 2496
rect 4908 2400 10824 2428
rect 3881 2391 3939 2397
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 18156 2437 18184 2468
rect 20530 2456 20536 2468
rect 20588 2456 20594 2508
rect 21637 2499 21695 2505
rect 21637 2465 21649 2499
rect 21683 2496 21695 2499
rect 22554 2496 22560 2508
rect 21683 2468 22560 2496
rect 21683 2465 21695 2468
rect 21637 2459 21695 2465
rect 22554 2456 22560 2468
rect 22612 2456 22618 2508
rect 24121 2499 24179 2505
rect 24121 2465 24133 2499
rect 24167 2496 24179 2499
rect 24167 2468 24486 2496
rect 24167 2465 24179 2468
rect 24121 2459 24179 2465
rect 15565 2431 15623 2437
rect 15565 2428 15577 2431
rect 13780 2400 15577 2428
rect 13780 2388 13786 2400
rect 15565 2397 15577 2400
rect 15611 2428 15623 2431
rect 18141 2431 18199 2437
rect 15611 2400 17816 2428
rect 15611 2397 15623 2400
rect 15565 2391 15623 2397
rect 17788 2372 17816 2400
rect 18141 2397 18153 2431
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 21913 2431 21971 2437
rect 21913 2428 21925 2431
rect 18279 2400 21925 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 21913 2397 21925 2400
rect 21959 2428 21971 2431
rect 22186 2428 22192 2440
rect 21959 2400 22192 2428
rect 21959 2397 21971 2400
rect 21913 2391 21971 2397
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 5994 2360 6000 2372
rect 5123 2332 6000 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 5994 2320 6000 2332
rect 6052 2320 6058 2372
rect 7834 2320 7840 2372
rect 7892 2360 7898 2372
rect 8113 2363 8171 2369
rect 8113 2360 8125 2363
rect 7892 2332 8125 2360
rect 7892 2320 7898 2332
rect 8113 2329 8125 2332
rect 8159 2329 8171 2363
rect 8113 2323 8171 2329
rect 13265 2363 13323 2369
rect 13265 2329 13277 2363
rect 13311 2360 13323 2363
rect 15654 2360 15660 2372
rect 13311 2332 15660 2360
rect 13311 2329 13323 2332
rect 13265 2323 13323 2329
rect 15654 2320 15660 2332
rect 15712 2320 15718 2372
rect 17770 2320 17776 2372
rect 17828 2360 17834 2372
rect 18248 2360 18276 2391
rect 22186 2388 22192 2400
rect 22244 2388 22250 2440
rect 18874 2360 18880 2372
rect 17828 2332 18276 2360
rect 18835 2332 18880 2360
rect 17828 2320 17834 2332
rect 18874 2320 18880 2332
rect 18932 2320 18938 2372
rect 20254 2360 20260 2372
rect 20215 2332 20260 2360
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 21634 2320 21640 2372
rect 21692 2360 21698 2372
rect 22925 2363 22983 2369
rect 22925 2360 22937 2363
rect 21692 2332 22937 2360
rect 21692 2320 21698 2332
rect 22925 2329 22937 2332
rect 22971 2329 22983 2363
rect 23934 2360 23940 2372
rect 23895 2332 23940 2360
rect 22925 2323 22983 2329
rect 23934 2320 23940 2332
rect 23992 2320 23998 2372
rect 24458 2360 24486 2468
rect 25866 2456 25872 2508
rect 25924 2496 25930 2508
rect 25961 2499 26019 2505
rect 25961 2496 25973 2499
rect 25924 2468 25973 2496
rect 25924 2456 25930 2468
rect 25961 2465 25973 2468
rect 26007 2465 26019 2499
rect 26326 2496 26332 2508
rect 26287 2468 26332 2496
rect 25961 2459 26019 2465
rect 26326 2456 26332 2468
rect 26384 2456 26390 2508
rect 28445 2499 28503 2505
rect 28445 2465 28457 2499
rect 28491 2496 28503 2499
rect 28994 2496 29000 2508
rect 28491 2468 29000 2496
rect 28491 2465 28503 2468
rect 28445 2459 28503 2465
rect 28994 2456 29000 2468
rect 29052 2496 29058 2508
rect 29288 2496 29316 2536
rect 30561 2533 30573 2536
rect 30607 2533 30619 2567
rect 31478 2564 31484 2576
rect 31439 2536 31484 2564
rect 30561 2527 30619 2533
rect 31478 2524 31484 2536
rect 31536 2524 31542 2576
rect 48317 2567 48375 2573
rect 48317 2564 48329 2567
rect 31588 2536 48329 2564
rect 29052 2468 29316 2496
rect 29365 2499 29423 2505
rect 29052 2456 29058 2468
rect 29365 2465 29377 2499
rect 29411 2496 29423 2499
rect 29454 2496 29460 2508
rect 29411 2468 29460 2496
rect 29411 2465 29423 2468
rect 29365 2459 29423 2465
rect 29454 2456 29460 2468
rect 29512 2456 29518 2508
rect 29641 2499 29699 2505
rect 29641 2465 29653 2499
rect 29687 2496 29699 2499
rect 29730 2496 29736 2508
rect 29687 2468 29736 2496
rect 29687 2465 29699 2468
rect 29641 2459 29699 2465
rect 29730 2456 29736 2468
rect 29788 2456 29794 2508
rect 26050 2428 26056 2440
rect 26011 2400 26056 2428
rect 26050 2388 26056 2400
rect 26108 2388 26114 2440
rect 26142 2388 26148 2440
rect 26200 2428 26206 2440
rect 31588 2428 31616 2536
rect 48317 2533 48329 2536
rect 48363 2533 48375 2567
rect 50617 2567 50675 2573
rect 48317 2527 48375 2533
rect 48516 2536 49740 2564
rect 32493 2499 32551 2505
rect 32493 2465 32505 2499
rect 32539 2465 32551 2499
rect 32493 2459 32551 2465
rect 26200 2400 31616 2428
rect 26200 2388 26206 2400
rect 25317 2363 25375 2369
rect 25317 2360 25329 2363
rect 24458 2332 25329 2360
rect 25317 2329 25329 2332
rect 25363 2360 25375 2363
rect 28258 2360 28264 2372
rect 25363 2332 28264 2360
rect 25363 2329 25375 2332
rect 25317 2323 25375 2329
rect 28258 2320 28264 2332
rect 28316 2320 28322 2372
rect 31294 2360 31300 2372
rect 31255 2332 31300 2360
rect 31294 2320 31300 2332
rect 31352 2320 31358 2372
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 3786 2292 3792 2304
rect 3283 2264 3792 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 5718 2292 5724 2304
rect 5679 2264 5724 2292
rect 5718 2252 5724 2264
rect 5776 2252 5782 2304
rect 7558 2292 7564 2304
rect 7519 2264 7564 2292
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 10781 2295 10839 2301
rect 10781 2261 10793 2295
rect 10827 2292 10839 2295
rect 12342 2292 12348 2304
rect 10827 2264 12348 2292
rect 10827 2261 10839 2264
rect 10781 2255 10839 2261
rect 12342 2252 12348 2264
rect 12400 2252 12406 2304
rect 12437 2295 12495 2301
rect 12437 2261 12449 2295
rect 12483 2292 12495 2295
rect 13722 2292 13728 2304
rect 12483 2264 13728 2292
rect 12483 2261 12495 2264
rect 12437 2255 12495 2261
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 13814 2252 13820 2304
rect 13872 2292 13878 2304
rect 13909 2295 13967 2301
rect 13909 2292 13921 2295
rect 13872 2264 13921 2292
rect 13872 2252 13878 2264
rect 13909 2261 13921 2264
rect 13955 2261 13967 2295
rect 17678 2292 17684 2304
rect 17639 2264 17684 2292
rect 13909 2255 13967 2261
rect 17678 2252 17684 2264
rect 17736 2252 17742 2304
rect 21358 2292 21364 2304
rect 21319 2264 21364 2292
rect 21358 2252 21364 2264
rect 21416 2252 21422 2304
rect 32508 2292 32536 2459
rect 33226 2456 33232 2508
rect 33284 2496 33290 2508
rect 33781 2499 33839 2505
rect 33781 2496 33793 2499
rect 33284 2468 33793 2496
rect 33284 2456 33290 2468
rect 33781 2465 33793 2468
rect 33827 2465 33839 2499
rect 33781 2459 33839 2465
rect 34885 2499 34943 2505
rect 34885 2465 34897 2499
rect 34931 2465 34943 2499
rect 34885 2459 34943 2465
rect 35345 2499 35403 2505
rect 35345 2465 35357 2499
rect 35391 2496 35403 2499
rect 36078 2496 36084 2508
rect 35391 2468 36084 2496
rect 35391 2465 35403 2468
rect 35345 2459 35403 2465
rect 34900 2428 34928 2459
rect 36078 2456 36084 2468
rect 36136 2456 36142 2508
rect 36262 2496 36268 2508
rect 36223 2468 36268 2496
rect 36262 2456 36268 2468
rect 36320 2456 36326 2508
rect 36538 2496 36544 2508
rect 36499 2468 36544 2496
rect 36538 2456 36544 2468
rect 36596 2456 36602 2508
rect 37553 2499 37611 2505
rect 37553 2465 37565 2499
rect 37599 2465 37611 2499
rect 37553 2459 37611 2465
rect 37568 2428 37596 2459
rect 37826 2456 37832 2508
rect 37884 2496 37890 2508
rect 39114 2496 39120 2508
rect 37884 2468 37929 2496
rect 39075 2468 39120 2496
rect 37884 2456 37890 2468
rect 39114 2456 39120 2468
rect 39172 2456 39178 2508
rect 39298 2456 39304 2508
rect 39356 2496 39362 2508
rect 39758 2496 39764 2508
rect 39356 2468 39764 2496
rect 39356 2456 39362 2468
rect 39758 2456 39764 2468
rect 39816 2496 39822 2508
rect 40313 2499 40371 2505
rect 40313 2496 40325 2499
rect 39816 2468 40325 2496
rect 39816 2456 39822 2468
rect 40313 2465 40325 2468
rect 40359 2465 40371 2499
rect 40313 2459 40371 2465
rect 40402 2456 40408 2508
rect 40460 2496 40466 2508
rect 41598 2496 41604 2508
rect 40460 2468 40505 2496
rect 41559 2468 41604 2496
rect 40460 2456 40466 2468
rect 41598 2456 41604 2468
rect 41656 2456 41662 2508
rect 41782 2496 41788 2508
rect 41743 2468 41788 2496
rect 41782 2456 41788 2468
rect 41840 2456 41846 2508
rect 43257 2499 43315 2505
rect 43257 2496 43269 2499
rect 42490 2468 43269 2496
rect 39850 2428 39856 2440
rect 34900 2400 36492 2428
rect 37568 2400 39856 2428
rect 36464 2372 36492 2400
rect 39850 2388 39856 2400
rect 39908 2388 39914 2440
rect 40589 2431 40647 2437
rect 40589 2397 40601 2431
rect 40635 2428 40647 2431
rect 41230 2428 41236 2440
rect 40635 2400 41236 2428
rect 40635 2397 40647 2400
rect 40589 2391 40647 2397
rect 41230 2388 41236 2400
rect 41288 2388 41294 2440
rect 41800 2400 42012 2428
rect 32677 2363 32735 2369
rect 32677 2329 32689 2363
rect 32723 2360 32735 2363
rect 35434 2360 35440 2372
rect 32723 2332 35440 2360
rect 32723 2329 32735 2332
rect 32677 2323 32735 2329
rect 35434 2320 35440 2332
rect 35492 2320 35498 2372
rect 36446 2320 36452 2372
rect 36504 2320 36510 2372
rect 36541 2363 36599 2369
rect 36541 2329 36553 2363
rect 36587 2360 36599 2363
rect 41800 2360 41828 2400
rect 36587 2332 41828 2360
rect 41877 2363 41935 2369
rect 36587 2329 36599 2332
rect 36541 2323 36599 2329
rect 41877 2329 41889 2363
rect 41923 2329 41935 2363
rect 41984 2360 42012 2400
rect 42058 2388 42064 2440
rect 42116 2428 42122 2440
rect 42490 2428 42518 2468
rect 43257 2465 43269 2468
rect 43303 2496 43315 2499
rect 43303 2468 44220 2496
rect 43303 2465 43315 2468
rect 43257 2459 43315 2465
rect 44192 2440 44220 2468
rect 44542 2456 44548 2508
rect 44600 2496 44606 2508
rect 44910 2496 44916 2508
rect 44600 2468 44916 2496
rect 44600 2456 44606 2468
rect 44910 2456 44916 2468
rect 44968 2456 44974 2508
rect 45005 2499 45063 2505
rect 45005 2465 45017 2499
rect 45051 2496 45063 2499
rect 45554 2496 45560 2508
rect 45051 2468 45560 2496
rect 45051 2465 45063 2468
rect 45005 2459 45063 2465
rect 45554 2456 45560 2468
rect 45612 2456 45618 2508
rect 45738 2496 45744 2508
rect 45699 2468 45744 2496
rect 45738 2456 45744 2468
rect 45796 2456 45802 2508
rect 45925 2499 45983 2505
rect 45925 2465 45937 2499
rect 45971 2496 45983 2499
rect 46014 2496 46020 2508
rect 45971 2468 46020 2496
rect 45971 2465 45983 2468
rect 45925 2459 45983 2465
rect 46014 2456 46020 2468
rect 46072 2456 46078 2508
rect 47302 2496 47308 2508
rect 47263 2468 47308 2496
rect 47302 2456 47308 2468
rect 47360 2456 47366 2508
rect 48406 2496 48412 2508
rect 47504 2468 48412 2496
rect 42116 2400 42518 2428
rect 43165 2431 43223 2437
rect 42116 2388 42122 2400
rect 43165 2397 43177 2431
rect 43211 2428 43223 2431
rect 43806 2428 43812 2440
rect 43211 2400 43812 2428
rect 43211 2397 43223 2400
rect 43165 2391 43223 2397
rect 43806 2388 43812 2400
rect 43864 2388 43870 2440
rect 44174 2388 44180 2440
rect 44232 2428 44238 2440
rect 45189 2431 45247 2437
rect 45189 2428 45201 2431
rect 44232 2400 45201 2428
rect 44232 2388 44238 2400
rect 45189 2397 45201 2400
rect 45235 2397 45247 2431
rect 47394 2428 47400 2440
rect 47355 2400 47400 2428
rect 45189 2391 45247 2397
rect 47394 2388 47400 2400
rect 47452 2388 47458 2440
rect 47504 2360 47532 2468
rect 48406 2456 48412 2468
rect 48464 2456 48470 2508
rect 47581 2431 47639 2437
rect 47581 2397 47593 2431
rect 47627 2397 47639 2431
rect 48516 2428 48544 2536
rect 48593 2499 48651 2505
rect 48593 2465 48605 2499
rect 48639 2496 48651 2499
rect 49510 2496 49516 2508
rect 48639 2468 49516 2496
rect 48639 2465 48651 2468
rect 48593 2459 48651 2465
rect 49510 2456 49516 2468
rect 49568 2456 49574 2508
rect 47581 2391 47639 2397
rect 48240 2400 48544 2428
rect 49712 2428 49740 2536
rect 50617 2533 50629 2567
rect 50663 2564 50675 2567
rect 52270 2564 52276 2576
rect 50663 2536 52276 2564
rect 50663 2533 50675 2536
rect 50617 2527 50675 2533
rect 52270 2524 52276 2536
rect 52328 2524 52334 2576
rect 54110 2524 54116 2576
rect 54168 2564 54174 2576
rect 55125 2567 55183 2573
rect 55125 2564 55137 2567
rect 54168 2536 55137 2564
rect 54168 2524 54174 2536
rect 55125 2533 55137 2536
rect 55171 2533 55183 2567
rect 55125 2527 55183 2533
rect 55582 2524 55588 2576
rect 55640 2564 55646 2576
rect 56597 2567 56655 2573
rect 56597 2564 56609 2567
rect 55640 2536 56609 2564
rect 55640 2524 55646 2536
rect 56597 2533 56609 2536
rect 56643 2533 56655 2567
rect 56597 2527 56655 2533
rect 50522 2496 50528 2508
rect 50483 2468 50528 2496
rect 50522 2456 50528 2468
rect 50580 2456 50586 2508
rect 52362 2456 52368 2508
rect 52420 2496 52426 2508
rect 52457 2499 52515 2505
rect 52457 2496 52469 2499
rect 52420 2468 52469 2496
rect 52420 2456 52426 2468
rect 52457 2465 52469 2468
rect 52503 2465 52515 2499
rect 52457 2459 52515 2465
rect 53374 2456 53380 2508
rect 53432 2496 53438 2508
rect 53561 2499 53619 2505
rect 53561 2496 53573 2499
rect 53432 2468 53573 2496
rect 53432 2456 53438 2468
rect 53561 2465 53573 2468
rect 53607 2465 53619 2499
rect 53561 2459 53619 2465
rect 55674 2456 55680 2508
rect 55732 2496 55738 2508
rect 55861 2499 55919 2505
rect 55861 2496 55873 2499
rect 55732 2468 55873 2496
rect 55732 2456 55738 2468
rect 55861 2465 55873 2468
rect 55907 2465 55919 2499
rect 57698 2496 57704 2508
rect 57659 2468 57704 2496
rect 55861 2459 55919 2465
rect 57698 2456 57704 2468
rect 57756 2456 57762 2508
rect 58066 2496 58072 2508
rect 57979 2468 58072 2496
rect 58066 2456 58072 2468
rect 58124 2496 58130 2508
rect 59354 2496 59360 2508
rect 58124 2468 59360 2496
rect 58124 2456 58130 2468
rect 59354 2456 59360 2468
rect 59412 2456 59418 2508
rect 50709 2431 50767 2437
rect 50709 2428 50721 2431
rect 49712 2400 50721 2428
rect 41984 2332 45048 2360
rect 41877 2323 41935 2329
rect 35342 2292 35348 2304
rect 32508 2264 35348 2292
rect 35342 2252 35348 2264
rect 35400 2252 35406 2304
rect 37274 2252 37280 2304
rect 37332 2292 37338 2304
rect 39025 2295 39083 2301
rect 39025 2292 39037 2295
rect 37332 2264 39037 2292
rect 37332 2252 37338 2264
rect 39025 2261 39037 2264
rect 39071 2261 39083 2295
rect 41892 2292 41920 2323
rect 42518 2292 42524 2304
rect 41892 2264 42524 2292
rect 39025 2255 39083 2261
rect 42518 2252 42524 2264
rect 42576 2252 42582 2304
rect 42702 2292 42708 2304
rect 42663 2264 42708 2292
rect 42702 2252 42708 2264
rect 42760 2252 42766 2304
rect 45020 2292 45048 2332
rect 45204 2332 47532 2360
rect 45204 2292 45232 2332
rect 45020 2264 45232 2292
rect 46290 2252 46296 2304
rect 46348 2292 46354 2304
rect 47596 2292 47624 2391
rect 48240 2292 48268 2400
rect 50709 2397 50721 2400
rect 50755 2428 50767 2431
rect 50798 2428 50804 2440
rect 50755 2400 50804 2428
rect 50755 2397 50767 2400
rect 50709 2391 50767 2397
rect 50798 2388 50804 2400
rect 50856 2388 50862 2440
rect 48317 2363 48375 2369
rect 48317 2329 48329 2363
rect 48363 2360 48375 2363
rect 48363 2332 53604 2360
rect 48363 2329 48375 2332
rect 48317 2323 48375 2329
rect 48498 2292 48504 2304
rect 46348 2264 48268 2292
rect 48459 2264 48504 2292
rect 46348 2252 46354 2264
rect 48498 2252 48504 2264
rect 48556 2252 48562 2304
rect 49329 2295 49387 2301
rect 49329 2261 49341 2295
rect 49375 2292 49387 2295
rect 49510 2292 49516 2304
rect 49375 2264 49516 2292
rect 49375 2261 49387 2264
rect 49329 2255 49387 2261
rect 49510 2252 49516 2264
rect 49568 2252 49574 2304
rect 50157 2295 50215 2301
rect 50157 2261 50169 2295
rect 50203 2292 50215 2295
rect 50614 2292 50620 2304
rect 50203 2264 50620 2292
rect 50203 2261 50215 2264
rect 50157 2255 50215 2261
rect 50614 2252 50620 2264
rect 50672 2252 50678 2304
rect 53466 2292 53472 2304
rect 53427 2264 53472 2292
rect 53466 2252 53472 2264
rect 53524 2252 53530 2304
rect 53576 2292 53604 2332
rect 54294 2320 54300 2372
rect 54352 2360 54358 2372
rect 54941 2363 54999 2369
rect 54941 2360 54953 2363
rect 54352 2332 54953 2360
rect 54352 2320 54358 2332
rect 54941 2329 54953 2332
rect 54987 2329 54999 2363
rect 54941 2323 54999 2329
rect 56134 2320 56140 2372
rect 56192 2360 56198 2372
rect 56413 2363 56471 2369
rect 56413 2360 56425 2363
rect 56192 2332 56425 2360
rect 56192 2320 56198 2332
rect 56413 2329 56425 2332
rect 56459 2329 56471 2363
rect 56413 2323 56471 2329
rect 55769 2295 55827 2301
rect 55769 2292 55781 2295
rect 53576 2264 55781 2292
rect 55769 2261 55781 2264
rect 55815 2261 55827 2295
rect 55769 2255 55827 2261
rect 55858 2252 55864 2304
rect 55916 2292 55922 2304
rect 57238 2292 57244 2304
rect 55916 2264 57244 2292
rect 55916 2252 55922 2264
rect 57238 2252 57244 2264
rect 57296 2252 57302 2304
rect 1104 2202 58880 2224
rect 1104 2150 10614 2202
rect 10666 2150 10678 2202
rect 10730 2150 10742 2202
rect 10794 2150 10806 2202
rect 10858 2150 29878 2202
rect 29930 2150 29942 2202
rect 29994 2150 30006 2202
rect 30058 2150 30070 2202
rect 30122 2150 49142 2202
rect 49194 2150 49206 2202
rect 49258 2150 49270 2202
rect 49322 2150 49334 2202
rect 49386 2150 58880 2202
rect 1104 2128 58880 2150
rect 13078 2048 13084 2100
rect 13136 2088 13142 2100
rect 37366 2088 37372 2100
rect 13136 2060 37372 2088
rect 13136 2048 13142 2060
rect 37366 2048 37372 2060
rect 37424 2048 37430 2100
rect 40310 2048 40316 2100
rect 40368 2088 40374 2100
rect 48498 2088 48504 2100
rect 40368 2060 48504 2088
rect 40368 2048 40374 2060
rect 48498 2048 48504 2060
rect 48556 2048 48562 2100
rect 24302 1980 24308 2032
rect 24360 2020 24366 2032
rect 42702 2020 42708 2032
rect 24360 1992 42708 2020
rect 24360 1980 24366 1992
rect 42702 1980 42708 1992
rect 42760 1980 42766 2032
rect 47394 1980 47400 2032
rect 47452 2020 47458 2032
rect 56686 2020 56692 2032
rect 47452 1992 56692 2020
rect 47452 1980 47458 1992
rect 56686 1980 56692 1992
rect 56744 1980 56750 2032
rect 1854 1912 1860 1964
rect 1912 1952 1918 1964
rect 17678 1952 17684 1964
rect 1912 1924 17684 1952
rect 1912 1912 1918 1924
rect 17678 1912 17684 1924
rect 17736 1912 17742 1964
rect 18598 1912 18604 1964
rect 18656 1952 18662 1964
rect 41506 1952 41512 1964
rect 18656 1924 41512 1952
rect 18656 1912 18662 1924
rect 41506 1912 41512 1924
rect 41564 1912 41570 1964
rect 42518 1912 42524 1964
rect 42576 1952 42582 1964
rect 48317 1955 48375 1961
rect 48317 1952 48329 1955
rect 42576 1924 48329 1952
rect 42576 1912 42582 1924
rect 48317 1921 48329 1924
rect 48363 1921 48375 1955
rect 48317 1915 48375 1921
rect 48406 1912 48412 1964
rect 48464 1952 48470 1964
rect 55858 1952 55864 1964
rect 48464 1924 55864 1952
rect 48464 1912 48470 1924
rect 55858 1912 55864 1924
rect 55916 1912 55922 1964
rect 14918 1844 14924 1896
rect 14976 1884 14982 1896
rect 21358 1884 21364 1896
rect 14976 1856 21364 1884
rect 14976 1844 14982 1856
rect 21358 1844 21364 1856
rect 21416 1844 21422 1896
rect 22002 1844 22008 1896
rect 22060 1884 22066 1896
rect 53466 1884 53472 1896
rect 22060 1856 53472 1884
rect 22060 1844 22066 1856
rect 53466 1844 53472 1856
rect 53524 1844 53530 1896
rect 12342 1776 12348 1828
rect 12400 1816 12406 1828
rect 20070 1816 20076 1828
rect 12400 1788 20076 1816
rect 12400 1776 12406 1788
rect 20070 1776 20076 1788
rect 20128 1776 20134 1828
rect 26050 1776 26056 1828
rect 26108 1816 26114 1828
rect 52362 1816 52368 1828
rect 26108 1788 52368 1816
rect 26108 1776 26114 1788
rect 52362 1776 52368 1788
rect 52420 1776 52426 1828
rect 5718 1708 5724 1760
rect 5776 1748 5782 1760
rect 47302 1748 47308 1760
rect 5776 1720 47308 1748
rect 5776 1708 5782 1720
rect 47302 1708 47308 1720
rect 47360 1708 47366 1760
rect 48317 1751 48375 1757
rect 48317 1717 48329 1751
rect 48363 1748 48375 1751
rect 56502 1748 56508 1760
rect 48363 1720 56508 1748
rect 48363 1717 48375 1720
rect 48317 1711 48375 1717
rect 56502 1708 56508 1720
rect 56560 1708 56566 1760
rect 3786 1640 3792 1692
rect 3844 1680 3850 1692
rect 28350 1680 28356 1692
rect 3844 1652 28356 1680
rect 3844 1640 3850 1652
rect 28350 1640 28356 1652
rect 28408 1640 28414 1692
rect 33778 1640 33784 1692
rect 33836 1680 33842 1692
rect 50522 1680 50528 1692
rect 33836 1652 50528 1680
rect 33836 1640 33842 1652
rect 50522 1640 50528 1652
rect 50580 1640 50586 1692
rect 7558 1572 7564 1624
rect 7616 1612 7622 1624
rect 39758 1612 39764 1624
rect 7616 1584 39764 1612
rect 7616 1572 7622 1584
rect 39758 1572 39764 1584
rect 39816 1572 39822 1624
rect 13722 1504 13728 1556
rect 13780 1544 13786 1556
rect 44910 1544 44916 1556
rect 13780 1516 44916 1544
rect 13780 1504 13786 1516
rect 44910 1504 44916 1516
rect 44968 1504 44974 1556
<< via1 >>
rect 17040 28092 17092 28144
rect 18604 28092 18656 28144
rect 18972 28092 19024 28144
rect 37464 28092 37516 28144
rect 16488 28024 16540 28076
rect 24308 28024 24360 28076
rect 5724 27956 5776 28008
rect 17408 27956 17460 28008
rect 20628 27956 20680 28008
rect 29736 27956 29788 28008
rect 8024 27888 8076 27940
rect 34336 28024 34388 28076
rect 33968 27956 34020 28008
rect 45376 27956 45428 28008
rect 30196 27888 30248 27940
rect 34612 27888 34664 27940
rect 9404 27820 9456 27872
rect 47032 27820 47084 27872
rect 20246 27718 20298 27770
rect 20310 27718 20362 27770
rect 20374 27718 20426 27770
rect 20438 27718 20490 27770
rect 39510 27718 39562 27770
rect 39574 27718 39626 27770
rect 39638 27718 39690 27770
rect 39702 27718 39754 27770
rect 3240 27616 3292 27668
rect 8024 27659 8076 27668
rect 8024 27625 8033 27659
rect 8033 27625 8067 27659
rect 8067 27625 8076 27659
rect 8024 27616 8076 27625
rect 8116 27616 8168 27668
rect 13820 27659 13872 27668
rect 2780 27548 2832 27600
rect 5540 27591 5592 27600
rect 5540 27557 5549 27591
rect 5549 27557 5583 27591
rect 5583 27557 5592 27591
rect 5540 27548 5592 27557
rect 5724 27591 5776 27600
rect 5724 27557 5733 27591
rect 5733 27557 5767 27591
rect 5767 27557 5776 27591
rect 5724 27548 5776 27557
rect 7840 27548 7892 27600
rect 9680 27591 9732 27600
rect 9680 27557 9689 27591
rect 9689 27557 9723 27591
rect 9723 27557 9732 27591
rect 9680 27548 9732 27557
rect 10600 27591 10652 27600
rect 10600 27557 10609 27591
rect 10609 27557 10643 27591
rect 10643 27557 10652 27591
rect 10600 27548 10652 27557
rect 11980 27591 12032 27600
rect 11980 27557 11989 27591
rect 11989 27557 12023 27591
rect 12023 27557 12032 27591
rect 11980 27548 12032 27557
rect 12440 27591 12492 27600
rect 12440 27557 12449 27591
rect 12449 27557 12483 27591
rect 12483 27557 12492 27591
rect 12440 27548 12492 27557
rect 13820 27625 13829 27659
rect 13829 27625 13863 27659
rect 13863 27625 13872 27659
rect 13820 27616 13872 27625
rect 14740 27548 14792 27600
rect 16120 27548 16172 27600
rect 16488 27591 16540 27600
rect 16488 27557 16497 27591
rect 16497 27557 16531 27591
rect 16531 27557 16540 27591
rect 16488 27548 16540 27557
rect 17960 27548 18012 27600
rect 19340 27591 19392 27600
rect 19340 27557 19349 27591
rect 19349 27557 19383 27591
rect 19383 27557 19392 27591
rect 19340 27548 19392 27557
rect 20628 27591 20680 27600
rect 20628 27557 20637 27591
rect 20637 27557 20671 27591
rect 20671 27557 20680 27591
rect 20628 27548 20680 27557
rect 940 27480 992 27532
rect 2228 27480 2280 27532
rect 3240 27523 3292 27532
rect 3240 27489 3249 27523
rect 3249 27489 3283 27523
rect 3283 27489 3292 27523
rect 3240 27480 3292 27489
rect 3884 27480 3936 27532
rect 5172 27480 5224 27532
rect 4896 27455 4948 27464
rect 4896 27421 4905 27455
rect 4905 27421 4939 27455
rect 4939 27421 4948 27455
rect 4896 27412 4948 27421
rect 6920 27387 6972 27396
rect 1768 27276 1820 27328
rect 4436 27276 4488 27328
rect 6920 27353 6929 27387
rect 6929 27353 6963 27387
rect 6963 27353 6972 27387
rect 6920 27344 6972 27353
rect 10416 27480 10468 27532
rect 13544 27480 13596 27532
rect 15016 27480 15068 27532
rect 15844 27480 15896 27532
rect 17684 27523 17736 27532
rect 17684 27489 17693 27523
rect 17693 27489 17727 27523
rect 17727 27489 17736 27523
rect 17684 27480 17736 27489
rect 17868 27523 17920 27532
rect 17868 27489 17877 27523
rect 17877 27489 17911 27523
rect 17911 27489 17920 27523
rect 17868 27480 17920 27489
rect 18604 27523 18656 27532
rect 18604 27489 18613 27523
rect 18613 27489 18647 27523
rect 18647 27489 18656 27523
rect 18604 27480 18656 27489
rect 19800 27480 19852 27532
rect 20260 27523 20312 27532
rect 20260 27489 20269 27523
rect 20269 27489 20303 27523
rect 20303 27489 20312 27523
rect 20260 27480 20312 27489
rect 20444 27523 20496 27532
rect 20444 27489 20453 27523
rect 20453 27489 20487 27523
rect 20487 27489 20496 27523
rect 20444 27480 20496 27489
rect 20536 27480 20588 27532
rect 17040 27412 17092 27464
rect 17408 27412 17460 27464
rect 20720 27412 20772 27464
rect 25872 27616 25924 27668
rect 29920 27659 29972 27668
rect 29920 27625 29929 27659
rect 29929 27625 29963 27659
rect 29963 27625 29972 27659
rect 29920 27616 29972 27625
rect 31484 27616 31536 27668
rect 37832 27616 37884 27668
rect 23940 27591 23992 27600
rect 23940 27557 23949 27591
rect 23949 27557 23983 27591
rect 23983 27557 23992 27591
rect 23940 27548 23992 27557
rect 24492 27548 24544 27600
rect 22100 27480 22152 27532
rect 23756 27480 23808 27532
rect 24124 27523 24176 27532
rect 24124 27489 24133 27523
rect 24133 27489 24167 27523
rect 24167 27489 24176 27523
rect 24124 27480 24176 27489
rect 26976 27480 27028 27532
rect 27252 27412 27304 27464
rect 28540 27548 28592 27600
rect 29736 27548 29788 27600
rect 32220 27591 32272 27600
rect 29368 27480 29420 27532
rect 32220 27557 32229 27591
rect 32229 27557 32263 27591
rect 32263 27557 32272 27591
rect 32220 27548 32272 27557
rect 33968 27591 34020 27600
rect 33968 27557 33977 27591
rect 33977 27557 34011 27591
rect 34011 27557 34020 27591
rect 33968 27548 34020 27557
rect 34152 27591 34204 27600
rect 34152 27557 34161 27591
rect 34161 27557 34195 27591
rect 34195 27557 34204 27591
rect 34152 27548 34204 27557
rect 35440 27548 35492 27600
rect 37280 27548 37332 27600
rect 37556 27591 37608 27600
rect 37556 27557 37578 27591
rect 37578 27557 37608 27591
rect 37556 27548 37608 27557
rect 38016 27548 38068 27600
rect 40132 27548 40184 27600
rect 43260 27616 43312 27668
rect 47032 27659 47084 27668
rect 47032 27625 47041 27659
rect 47041 27625 47075 27659
rect 47075 27625 47084 27659
rect 47032 27616 47084 27625
rect 52920 27616 52972 27668
rect 54760 27616 54812 27668
rect 42800 27548 42852 27600
rect 43812 27548 43864 27600
rect 45560 27548 45612 27600
rect 46480 27548 46532 27600
rect 46940 27548 46992 27600
rect 48320 27548 48372 27600
rect 48964 27548 49016 27600
rect 51540 27548 51592 27600
rect 52000 27548 52052 27600
rect 53380 27548 53432 27600
rect 54300 27548 54352 27600
rect 55220 27548 55272 27600
rect 57980 27548 58032 27600
rect 31484 27412 31536 27464
rect 9864 27276 9916 27328
rect 17132 27276 17184 27328
rect 17500 27276 17552 27328
rect 25780 27276 25832 27328
rect 30288 27344 30340 27396
rect 33600 27480 33652 27532
rect 34428 27480 34480 27532
rect 36636 27480 36688 27532
rect 33508 27412 33560 27464
rect 39304 27523 39356 27532
rect 39304 27489 39313 27523
rect 39313 27489 39347 27523
rect 39347 27489 39356 27523
rect 39304 27480 39356 27489
rect 40224 27480 40276 27532
rect 41420 27480 41472 27532
rect 43536 27480 43588 27532
rect 44088 27480 44140 27532
rect 45836 27523 45888 27532
rect 28724 27319 28776 27328
rect 28724 27285 28733 27319
rect 28733 27285 28767 27319
rect 28767 27285 28776 27319
rect 28724 27276 28776 27285
rect 29184 27276 29236 27328
rect 36820 27344 36872 27396
rect 39028 27387 39080 27396
rect 39028 27353 39037 27387
rect 39037 27353 39071 27387
rect 39071 27353 39080 27387
rect 39028 27344 39080 27353
rect 39764 27412 39816 27464
rect 45836 27489 45845 27523
rect 45845 27489 45879 27523
rect 45879 27489 45888 27523
rect 45836 27480 45888 27489
rect 49516 27480 49568 27532
rect 50436 27523 50488 27532
rect 50436 27489 50445 27523
rect 50445 27489 50479 27523
rect 50479 27489 50488 27523
rect 50436 27480 50488 27489
rect 54392 27480 54444 27532
rect 56048 27480 56100 27532
rect 30472 27276 30524 27328
rect 31208 27276 31260 27328
rect 34888 27319 34940 27328
rect 34888 27285 34897 27319
rect 34897 27285 34931 27319
rect 34931 27285 34940 27319
rect 34888 27276 34940 27285
rect 38476 27276 38528 27328
rect 39120 27276 39172 27328
rect 55128 27344 55180 27396
rect 41788 27319 41840 27328
rect 41788 27285 41797 27319
rect 41797 27285 41831 27319
rect 41831 27285 41840 27319
rect 41788 27276 41840 27285
rect 48412 27319 48464 27328
rect 48412 27285 48421 27319
rect 48421 27285 48455 27319
rect 48455 27285 48464 27319
rect 48412 27276 48464 27285
rect 51172 27319 51224 27328
rect 51172 27285 51181 27319
rect 51181 27285 51215 27319
rect 51215 27285 51224 27319
rect 51172 27276 51224 27285
rect 52368 27319 52420 27328
rect 52368 27285 52377 27319
rect 52377 27285 52411 27319
rect 52411 27285 52420 27319
rect 52368 27276 52420 27285
rect 53472 27319 53524 27328
rect 53472 27285 53481 27319
rect 53481 27285 53515 27319
rect 53515 27285 53524 27319
rect 53472 27276 53524 27285
rect 57612 27276 57664 27328
rect 10614 27174 10666 27226
rect 10678 27174 10730 27226
rect 10742 27174 10794 27226
rect 10806 27174 10858 27226
rect 29878 27174 29930 27226
rect 29942 27174 29994 27226
rect 30006 27174 30058 27226
rect 30070 27174 30122 27226
rect 49142 27174 49194 27226
rect 49206 27174 49258 27226
rect 49270 27174 49322 27226
rect 49334 27174 49386 27226
rect 19984 27072 20036 27124
rect 20536 27072 20588 27124
rect 24124 27072 24176 27124
rect 25872 27072 25924 27124
rect 30196 27072 30248 27124
rect 30288 27072 30340 27124
rect 1400 27004 1452 27056
rect 3884 27004 3936 27056
rect 4252 27047 4304 27056
rect 4252 27013 4261 27047
rect 4261 27013 4295 27047
rect 4295 27013 4304 27047
rect 4252 27004 4304 27013
rect 6000 27004 6052 27056
rect 6920 27004 6972 27056
rect 5724 26936 5776 26988
rect 6460 26936 6512 26988
rect 1492 26911 1544 26920
rect 1492 26877 1501 26911
rect 1501 26877 1535 26911
rect 1535 26877 1544 26911
rect 1492 26868 1544 26877
rect 2872 26911 2924 26920
rect 2872 26877 2881 26911
rect 2881 26877 2915 26911
rect 2915 26877 2924 26911
rect 2872 26868 2924 26877
rect 4620 26868 4672 26920
rect 8116 26936 8168 26988
rect 8852 26936 8904 26988
rect 11244 26936 11296 26988
rect 16948 27004 17000 27056
rect 17684 27004 17736 27056
rect 17960 27047 18012 27056
rect 17960 27013 17969 27047
rect 17969 27013 18003 27047
rect 18003 27013 18012 27047
rect 17960 27004 18012 27013
rect 22284 27004 22336 27056
rect 22560 27047 22612 27056
rect 22560 27013 22569 27047
rect 22569 27013 22603 27047
rect 22603 27013 22612 27047
rect 22560 27004 22612 27013
rect 7380 26868 7432 26920
rect 8760 26868 8812 26920
rect 9404 26911 9456 26920
rect 9404 26877 9413 26911
rect 9413 26877 9447 26911
rect 9447 26877 9456 26911
rect 9404 26868 9456 26877
rect 10324 26868 10376 26920
rect 1676 26843 1728 26852
rect 1676 26809 1685 26843
rect 1685 26809 1719 26843
rect 1719 26809 1728 26843
rect 1676 26800 1728 26809
rect 3332 26800 3384 26852
rect 4896 26800 4948 26852
rect 7932 26800 7984 26852
rect 11980 26868 12032 26920
rect 12900 26911 12952 26920
rect 12900 26877 12909 26911
rect 12909 26877 12943 26911
rect 12943 26877 12952 26911
rect 12900 26868 12952 26877
rect 14280 26911 14332 26920
rect 14280 26877 14289 26911
rect 14289 26877 14323 26911
rect 14323 26877 14332 26911
rect 14280 26868 14332 26877
rect 15660 26868 15712 26920
rect 16396 26911 16448 26920
rect 16396 26877 16405 26911
rect 16405 26877 16439 26911
rect 16439 26877 16448 26911
rect 16396 26868 16448 26877
rect 16764 26868 16816 26920
rect 24308 26936 24360 26988
rect 27160 27004 27212 27056
rect 29000 27047 29052 27056
rect 29000 27013 29009 27047
rect 29009 27013 29043 27047
rect 29043 27013 29052 27047
rect 29000 27004 29052 27013
rect 29552 27047 29604 27056
rect 29552 27013 29561 27047
rect 29561 27013 29595 27047
rect 29595 27013 29604 27047
rect 29552 27004 29604 27013
rect 30840 27047 30892 27056
rect 30840 27013 30849 27047
rect 30849 27013 30883 27047
rect 30883 27013 30892 27047
rect 30840 27004 30892 27013
rect 29460 26936 29512 26988
rect 17500 26843 17552 26852
rect 8024 26732 8076 26784
rect 9680 26732 9732 26784
rect 11060 26775 11112 26784
rect 11060 26741 11069 26775
rect 11069 26741 11103 26775
rect 11103 26741 11112 26775
rect 11060 26732 11112 26741
rect 12256 26775 12308 26784
rect 12256 26741 12265 26775
rect 12265 26741 12299 26775
rect 12299 26741 12308 26775
rect 12256 26732 12308 26741
rect 12900 26732 12952 26784
rect 14464 26775 14516 26784
rect 14464 26741 14473 26775
rect 14473 26741 14507 26775
rect 14507 26741 14516 26775
rect 14464 26732 14516 26741
rect 15568 26775 15620 26784
rect 15568 26741 15577 26775
rect 15577 26741 15611 26775
rect 15611 26741 15620 26775
rect 15568 26732 15620 26741
rect 17500 26809 17509 26843
rect 17509 26809 17543 26843
rect 17543 26809 17552 26843
rect 17500 26800 17552 26809
rect 17684 26843 17736 26852
rect 17684 26809 17693 26843
rect 17693 26809 17727 26843
rect 17727 26809 17736 26843
rect 17684 26800 17736 26809
rect 18052 26800 18104 26852
rect 19064 26800 19116 26852
rect 20444 26868 20496 26920
rect 21088 26911 21140 26920
rect 21088 26877 21097 26911
rect 21097 26877 21131 26911
rect 21131 26877 21140 26911
rect 21088 26868 21140 26877
rect 22836 26868 22888 26920
rect 20260 26800 20312 26852
rect 22744 26843 22796 26852
rect 22744 26809 22753 26843
rect 22753 26809 22787 26843
rect 22787 26809 22796 26843
rect 22744 26800 22796 26809
rect 23204 26800 23256 26852
rect 23572 26868 23624 26920
rect 25320 26911 25372 26920
rect 25320 26877 25329 26911
rect 25329 26877 25363 26911
rect 25363 26877 25372 26911
rect 25320 26868 25372 26877
rect 26332 26868 26384 26920
rect 26884 26868 26936 26920
rect 28080 26911 28132 26920
rect 26608 26800 26660 26852
rect 27252 26800 27304 26852
rect 28080 26877 28089 26911
rect 28089 26877 28123 26911
rect 28123 26877 28132 26911
rect 28080 26868 28132 26877
rect 30472 26936 30524 26988
rect 28172 26843 28224 26852
rect 28172 26809 28181 26843
rect 28181 26809 28215 26843
rect 28215 26809 28224 26843
rect 28172 26800 28224 26809
rect 28356 26800 28408 26852
rect 33416 26936 33468 26988
rect 31760 26868 31812 26920
rect 31024 26843 31076 26852
rect 31024 26809 31033 26843
rect 31033 26809 31067 26843
rect 31067 26809 31076 26843
rect 31024 26800 31076 26809
rect 32588 26800 32640 26852
rect 33876 26868 33928 26920
rect 34704 26911 34756 26920
rect 34704 26877 34713 26911
rect 34713 26877 34747 26911
rect 34747 26877 34756 26911
rect 34704 26868 34756 26877
rect 19616 26732 19668 26784
rect 20720 26732 20772 26784
rect 20996 26775 21048 26784
rect 20996 26741 21005 26775
rect 21005 26741 21039 26775
rect 21039 26741 21048 26775
rect 20996 26732 21048 26741
rect 23572 26732 23624 26784
rect 25964 26732 26016 26784
rect 30932 26732 30984 26784
rect 33324 26732 33376 26784
rect 33508 26732 33560 26784
rect 34520 26775 34572 26784
rect 34520 26741 34529 26775
rect 34529 26741 34563 26775
rect 34563 26741 34572 26775
rect 34520 26732 34572 26741
rect 48320 27072 48372 27124
rect 52000 27072 52052 27124
rect 53380 27072 53432 27124
rect 39304 27004 39356 27056
rect 39856 27004 39908 27056
rect 41880 27047 41932 27056
rect 41880 27013 41889 27047
rect 41889 27013 41923 27047
rect 41923 27013 41932 27047
rect 41880 27004 41932 27013
rect 44088 27047 44140 27056
rect 44088 27013 44097 27047
rect 44097 27013 44131 27047
rect 44131 27013 44140 27047
rect 44088 27004 44140 27013
rect 44640 27047 44692 27056
rect 44640 27013 44649 27047
rect 44649 27013 44683 27047
rect 44683 27013 44692 27047
rect 44640 27004 44692 27013
rect 45376 27047 45428 27056
rect 45376 27013 45385 27047
rect 45385 27013 45419 27047
rect 45419 27013 45428 27047
rect 45376 27004 45428 27013
rect 47860 27047 47912 27056
rect 47860 27013 47869 27047
rect 47869 27013 47903 27047
rect 47903 27013 47912 27047
rect 47860 27004 47912 27013
rect 49700 27047 49752 27056
rect 49700 27013 49709 27047
rect 49709 27013 49743 27047
rect 49743 27013 49752 27047
rect 49700 27004 49752 27013
rect 50160 27047 50212 27056
rect 50160 27013 50169 27047
rect 50169 27013 50203 27047
rect 50203 27013 50212 27047
rect 50160 27004 50212 27013
rect 51080 27047 51132 27056
rect 51080 27013 51089 27047
rect 51089 27013 51123 27047
rect 51123 27013 51132 27047
rect 51080 27004 51132 27013
rect 56140 27047 56192 27056
rect 56140 27013 56149 27047
rect 56149 27013 56183 27047
rect 56183 27013 56192 27047
rect 56140 27004 56192 27013
rect 57520 27004 57572 27056
rect 41696 26936 41748 26988
rect 35808 26911 35860 26920
rect 35808 26877 35817 26911
rect 35817 26877 35851 26911
rect 35851 26877 35860 26911
rect 35808 26868 35860 26877
rect 36728 26911 36780 26920
rect 36728 26877 36737 26911
rect 36737 26877 36771 26911
rect 36771 26877 36780 26911
rect 36728 26868 36780 26877
rect 38660 26868 38712 26920
rect 39856 26911 39908 26920
rect 39856 26877 39865 26911
rect 39865 26877 39899 26911
rect 39899 26877 39908 26911
rect 39856 26868 39908 26877
rect 40040 26868 40092 26920
rect 40960 26868 41012 26920
rect 36268 26800 36320 26852
rect 40592 26843 40644 26852
rect 36176 26732 36228 26784
rect 40592 26809 40601 26843
rect 40601 26809 40635 26843
rect 40635 26809 40644 26843
rect 40592 26800 40644 26809
rect 41880 26868 41932 26920
rect 45100 26868 45152 26920
rect 54392 26911 54444 26920
rect 54392 26877 54401 26911
rect 54401 26877 54435 26911
rect 54435 26877 54444 26911
rect 54392 26868 54444 26877
rect 59360 26936 59412 26988
rect 42340 26800 42392 26852
rect 44456 26800 44508 26852
rect 47768 26800 47820 26852
rect 49976 26800 50028 26852
rect 41328 26775 41380 26784
rect 41328 26741 41337 26775
rect 41337 26741 41371 26775
rect 41371 26741 41380 26775
rect 41328 26732 41380 26741
rect 47860 26732 47912 26784
rect 54668 26800 54720 26852
rect 58072 26911 58124 26920
rect 58072 26877 58081 26911
rect 58081 26877 58115 26911
rect 58115 26877 58124 26911
rect 58072 26868 58124 26877
rect 55496 26775 55548 26784
rect 55496 26741 55505 26775
rect 55505 26741 55539 26775
rect 55539 26741 55548 26775
rect 55496 26732 55548 26741
rect 55680 26732 55732 26784
rect 57704 26800 57756 26852
rect 20246 26630 20298 26682
rect 20310 26630 20362 26682
rect 20374 26630 20426 26682
rect 20438 26630 20490 26682
rect 39510 26630 39562 26682
rect 39574 26630 39626 26682
rect 39638 26630 39690 26682
rect 39702 26630 39754 26682
rect 2596 26528 2648 26580
rect 4620 26528 4672 26580
rect 5724 26571 5776 26580
rect 5724 26537 5733 26571
rect 5733 26537 5767 26571
rect 5767 26537 5776 26571
rect 5724 26528 5776 26537
rect 7380 26571 7432 26580
rect 7380 26537 7389 26571
rect 7389 26537 7423 26571
rect 7423 26537 7432 26571
rect 7380 26528 7432 26537
rect 8116 26528 8168 26580
rect 8760 26528 8812 26580
rect 9772 26528 9824 26580
rect 10324 26571 10376 26580
rect 10324 26537 10333 26571
rect 10333 26537 10367 26571
rect 10367 26537 10376 26571
rect 10324 26528 10376 26537
rect 15660 26528 15712 26580
rect 17040 26571 17092 26580
rect 17040 26537 17049 26571
rect 17049 26537 17083 26571
rect 17083 26537 17092 26571
rect 17040 26528 17092 26537
rect 17132 26528 17184 26580
rect 17776 26528 17828 26580
rect 18972 26528 19024 26580
rect 1584 26503 1636 26512
rect 1584 26469 1593 26503
rect 1593 26469 1627 26503
rect 1627 26469 1636 26503
rect 1584 26460 1636 26469
rect 2228 26460 2280 26512
rect 4160 26460 4212 26512
rect 4436 26503 4488 26512
rect 4436 26469 4445 26503
rect 4445 26469 4479 26503
rect 4479 26469 4488 26503
rect 4436 26460 4488 26469
rect 4528 26460 4580 26512
rect 7932 26460 7984 26512
rect 9220 26460 9272 26512
rect 9680 26503 9732 26512
rect 9680 26469 9689 26503
rect 9689 26469 9723 26503
rect 9723 26469 9732 26503
rect 9680 26460 9732 26469
rect 11244 26460 11296 26512
rect 2320 26435 2372 26444
rect 2320 26401 2329 26435
rect 2329 26401 2363 26435
rect 2363 26401 2372 26435
rect 2320 26392 2372 26401
rect 10232 26435 10284 26444
rect 10232 26401 10241 26435
rect 10241 26401 10275 26435
rect 10275 26401 10284 26435
rect 10232 26392 10284 26401
rect 11152 26392 11204 26444
rect 14464 26460 14516 26512
rect 20076 26460 20128 26512
rect 20720 26528 20772 26580
rect 21180 26503 21232 26512
rect 16764 26392 16816 26444
rect 16948 26435 17000 26444
rect 16948 26401 16957 26435
rect 16957 26401 16991 26435
rect 16991 26401 17000 26435
rect 16948 26392 17000 26401
rect 4436 26256 4488 26308
rect 14188 26256 14240 26308
rect 17776 26392 17828 26444
rect 18880 26435 18932 26444
rect 17868 26324 17920 26376
rect 18880 26401 18889 26435
rect 18889 26401 18923 26435
rect 18923 26401 18932 26435
rect 18880 26392 18932 26401
rect 21180 26469 21189 26503
rect 21189 26469 21223 26503
rect 21223 26469 21232 26503
rect 21180 26460 21232 26469
rect 23480 26528 23532 26580
rect 27988 26528 28040 26580
rect 28080 26528 28132 26580
rect 31760 26528 31812 26580
rect 34152 26571 34204 26580
rect 34152 26537 34161 26571
rect 34161 26537 34195 26571
rect 34195 26537 34204 26571
rect 34152 26528 34204 26537
rect 35808 26571 35860 26580
rect 35808 26537 35817 26571
rect 35817 26537 35851 26571
rect 35851 26537 35860 26571
rect 35808 26528 35860 26537
rect 36268 26528 36320 26580
rect 41420 26528 41472 26580
rect 41696 26528 41748 26580
rect 47400 26528 47452 26580
rect 51540 26571 51592 26580
rect 51540 26537 51549 26571
rect 51549 26537 51583 26571
rect 51583 26537 51592 26571
rect 54668 26571 54720 26580
rect 51540 26528 51592 26537
rect 54668 26537 54677 26571
rect 54677 26537 54711 26571
rect 54711 26537 54720 26571
rect 54668 26528 54720 26537
rect 58072 26528 58124 26580
rect 26332 26460 26384 26512
rect 27620 26503 27672 26512
rect 27620 26469 27629 26503
rect 27629 26469 27663 26503
rect 27663 26469 27672 26503
rect 27620 26460 27672 26469
rect 33140 26503 33192 26512
rect 33140 26469 33149 26503
rect 33149 26469 33183 26503
rect 33183 26469 33192 26503
rect 33140 26460 33192 26469
rect 33324 26503 33376 26512
rect 33324 26469 33333 26503
rect 33333 26469 33367 26503
rect 33367 26469 33376 26503
rect 33324 26460 33376 26469
rect 38752 26503 38804 26512
rect 38752 26469 38761 26503
rect 38761 26469 38795 26503
rect 38795 26469 38804 26503
rect 38752 26460 38804 26469
rect 39396 26460 39448 26512
rect 39856 26460 39908 26512
rect 41880 26460 41932 26512
rect 55128 26503 55180 26512
rect 55128 26469 55137 26503
rect 55137 26469 55171 26503
rect 55171 26469 55180 26503
rect 55128 26460 55180 26469
rect 56600 26460 56652 26512
rect 58164 26503 58216 26512
rect 58164 26469 58173 26503
rect 58173 26469 58207 26503
rect 58207 26469 58216 26503
rect 58164 26460 58216 26469
rect 22284 26435 22336 26444
rect 22284 26401 22293 26435
rect 22293 26401 22327 26435
rect 22327 26401 22336 26435
rect 22284 26392 22336 26401
rect 26700 26392 26752 26444
rect 27804 26435 27856 26444
rect 27804 26401 27813 26435
rect 27813 26401 27847 26435
rect 27847 26401 27856 26435
rect 27804 26392 27856 26401
rect 30380 26392 30432 26444
rect 34060 26392 34112 26444
rect 34336 26392 34388 26444
rect 35716 26435 35768 26444
rect 35716 26401 35725 26435
rect 35725 26401 35759 26435
rect 35759 26401 35768 26435
rect 35716 26392 35768 26401
rect 36360 26392 36412 26444
rect 37280 26392 37332 26444
rect 37464 26392 37516 26444
rect 38200 26392 38252 26444
rect 38568 26392 38620 26444
rect 40500 26392 40552 26444
rect 41144 26435 41196 26444
rect 41144 26401 41153 26435
rect 41153 26401 41187 26435
rect 41187 26401 41196 26435
rect 41144 26392 41196 26401
rect 55036 26392 55088 26444
rect 56968 26392 57020 26444
rect 38660 26367 38712 26376
rect 19892 26256 19944 26308
rect 24492 26256 24544 26308
rect 37648 26299 37700 26308
rect 6368 26231 6420 26240
rect 6368 26197 6377 26231
rect 6377 26197 6411 26231
rect 6411 26197 6420 26231
rect 6368 26188 6420 26197
rect 11520 26188 11572 26240
rect 13544 26231 13596 26240
rect 13544 26197 13553 26231
rect 13553 26197 13587 26231
rect 13587 26197 13596 26231
rect 13544 26188 13596 26197
rect 15016 26188 15068 26240
rect 16948 26188 17000 26240
rect 18052 26188 18104 26240
rect 19524 26188 19576 26240
rect 22836 26188 22888 26240
rect 23204 26231 23256 26240
rect 23204 26197 23213 26231
rect 23213 26197 23247 26231
rect 23247 26197 23256 26231
rect 23204 26188 23256 26197
rect 26884 26188 26936 26240
rect 32588 26231 32640 26240
rect 32588 26197 32597 26231
rect 32597 26197 32631 26231
rect 32631 26197 32640 26231
rect 32588 26188 32640 26197
rect 34704 26231 34756 26240
rect 34704 26197 34713 26231
rect 34713 26197 34747 26231
rect 34747 26197 34756 26231
rect 34704 26188 34756 26197
rect 37648 26265 37657 26299
rect 37657 26265 37691 26299
rect 37691 26265 37700 26299
rect 37648 26256 37700 26265
rect 38660 26333 38669 26367
rect 38669 26333 38703 26367
rect 38703 26333 38712 26367
rect 38660 26324 38712 26333
rect 40592 26324 40644 26376
rect 57244 26324 57296 26376
rect 49424 26299 49476 26308
rect 49424 26265 49433 26299
rect 49433 26265 49467 26299
rect 49467 26265 49476 26299
rect 49424 26256 49476 26265
rect 38844 26188 38896 26240
rect 42340 26231 42392 26240
rect 42340 26197 42349 26231
rect 42349 26197 42383 26231
rect 42383 26197 42392 26231
rect 42340 26188 42392 26197
rect 44456 26231 44508 26240
rect 44456 26197 44465 26231
rect 44465 26197 44499 26231
rect 44499 26197 44508 26231
rect 44456 26188 44508 26197
rect 45836 26231 45888 26240
rect 45836 26197 45845 26231
rect 45845 26197 45879 26231
rect 45879 26197 45888 26231
rect 45836 26188 45888 26197
rect 49976 26231 50028 26240
rect 49976 26197 49985 26231
rect 49985 26197 50019 26231
rect 50019 26197 50028 26231
rect 49976 26188 50028 26197
rect 10614 26086 10666 26138
rect 10678 26086 10730 26138
rect 10742 26086 10794 26138
rect 10806 26086 10858 26138
rect 29878 26086 29930 26138
rect 29942 26086 29994 26138
rect 30006 26086 30058 26138
rect 30070 26086 30122 26138
rect 49142 26086 49194 26138
rect 49206 26086 49258 26138
rect 49270 26086 49322 26138
rect 49334 26086 49386 26138
rect 2320 25984 2372 26036
rect 3240 25984 3292 26036
rect 3516 25984 3568 26036
rect 4436 25984 4488 26036
rect 5172 25959 5224 25968
rect 5172 25925 5181 25959
rect 5181 25925 5215 25959
rect 5215 25925 5224 25959
rect 5172 25916 5224 25925
rect 1400 25891 1452 25900
rect 1400 25857 1409 25891
rect 1409 25857 1443 25891
rect 1443 25857 1452 25891
rect 1400 25848 1452 25857
rect 6368 25848 6420 25900
rect 8852 25916 8904 25968
rect 10232 25916 10284 25968
rect 11244 25916 11296 25968
rect 12900 25916 12952 25968
rect 16396 25916 16448 25968
rect 17684 25916 17736 25968
rect 18604 25916 18656 25968
rect 18972 25916 19024 25968
rect 2504 25780 2556 25832
rect 4896 25780 4948 25832
rect 9772 25823 9824 25832
rect 9772 25789 9787 25823
rect 9787 25789 9821 25823
rect 9821 25789 9824 25823
rect 9772 25780 9824 25789
rect 16948 25848 17000 25900
rect 17592 25780 17644 25832
rect 23204 25984 23256 26036
rect 33876 25984 33928 26036
rect 34060 25984 34112 26036
rect 34428 26027 34480 26036
rect 34428 25993 34437 26027
rect 34437 25993 34471 26027
rect 34471 25993 34480 26027
rect 34428 25984 34480 25993
rect 36360 25984 36412 26036
rect 37832 25984 37884 26036
rect 38476 26027 38528 26036
rect 38476 25993 38485 26027
rect 38485 25993 38519 26027
rect 38519 25993 38528 26027
rect 38476 25984 38528 25993
rect 38568 25984 38620 26036
rect 40132 25984 40184 26036
rect 40316 26027 40368 26036
rect 40316 25993 40325 26027
rect 40325 25993 40359 26027
rect 40359 25993 40368 26027
rect 40316 25984 40368 25993
rect 40960 26027 41012 26036
rect 40960 25993 40969 26027
rect 40969 25993 41003 26027
rect 41003 25993 41012 26027
rect 40960 25984 41012 25993
rect 41144 25984 41196 26036
rect 41604 25984 41656 26036
rect 55496 25984 55548 26036
rect 57244 26027 57296 26036
rect 57244 25993 57253 26027
rect 57253 25993 57287 26027
rect 57287 25993 57296 26027
rect 57244 25984 57296 25993
rect 19524 25916 19576 25968
rect 19616 25848 19668 25900
rect 32312 25916 32364 25968
rect 50436 25916 50488 25968
rect 55036 25959 55088 25968
rect 55036 25925 55045 25959
rect 55045 25925 55079 25959
rect 55079 25925 55088 25959
rect 55036 25916 55088 25925
rect 57980 25916 58032 25968
rect 20536 25780 20588 25832
rect 21088 25780 21140 25832
rect 23756 25780 23808 25832
rect 26332 25823 26384 25832
rect 26332 25789 26341 25823
rect 26341 25789 26375 25823
rect 26375 25789 26384 25823
rect 26332 25780 26384 25789
rect 26792 25823 26844 25832
rect 26792 25789 26801 25823
rect 26801 25789 26835 25823
rect 26835 25789 26844 25823
rect 26792 25780 26844 25789
rect 29460 25780 29512 25832
rect 33324 25823 33376 25832
rect 5724 25712 5776 25764
rect 30932 25712 30984 25764
rect 33324 25789 33333 25823
rect 33333 25789 33367 25823
rect 33367 25789 33376 25823
rect 33324 25780 33376 25789
rect 34980 25780 35032 25832
rect 36820 25780 36872 25832
rect 33508 25712 33560 25764
rect 37648 25848 37700 25900
rect 56048 25848 56100 25900
rect 58072 25848 58124 25900
rect 37556 25780 37608 25832
rect 37740 25780 37792 25832
rect 38660 25780 38712 25832
rect 39856 25823 39908 25832
rect 39856 25789 39865 25823
rect 39865 25789 39899 25823
rect 39899 25789 39908 25823
rect 39856 25780 39908 25789
rect 39948 25780 40000 25832
rect 41604 25780 41656 25832
rect 38016 25712 38068 25764
rect 38568 25712 38620 25764
rect 56692 25712 56744 25764
rect 9864 25687 9916 25696
rect 9864 25653 9873 25687
rect 9873 25653 9907 25687
rect 9907 25653 9916 25687
rect 9864 25644 9916 25653
rect 23664 25644 23716 25696
rect 57428 25644 57480 25696
rect 20246 25542 20298 25594
rect 20310 25542 20362 25594
rect 20374 25542 20426 25594
rect 20438 25542 20490 25594
rect 39510 25542 39562 25594
rect 39574 25542 39626 25594
rect 39638 25542 39690 25594
rect 39702 25542 39754 25594
rect 3332 25440 3384 25492
rect 9404 25440 9456 25492
rect 16764 25440 16816 25492
rect 17592 25440 17644 25492
rect 12256 25372 12308 25424
rect 32588 25440 32640 25492
rect 33876 25440 33928 25492
rect 35716 25440 35768 25492
rect 37464 25440 37516 25492
rect 38752 25440 38804 25492
rect 57428 25483 57480 25492
rect 57428 25449 57437 25483
rect 57437 25449 57471 25483
rect 57471 25449 57480 25483
rect 57428 25440 57480 25449
rect 17960 25372 18012 25424
rect 56876 25372 56928 25424
rect 58440 25372 58492 25424
rect 1400 25211 1452 25220
rect 1400 25177 1409 25211
rect 1409 25177 1443 25211
rect 1443 25177 1452 25211
rect 1400 25168 1452 25177
rect 16764 25304 16816 25356
rect 37740 25304 37792 25356
rect 33508 25279 33560 25288
rect 33508 25245 33517 25279
rect 33517 25245 33551 25279
rect 33551 25245 33560 25279
rect 33508 25236 33560 25245
rect 23664 25168 23716 25220
rect 36176 25211 36228 25220
rect 36176 25177 36185 25211
rect 36185 25177 36219 25211
rect 36219 25177 36228 25211
rect 36176 25168 36228 25177
rect 37464 25168 37516 25220
rect 36452 25100 36504 25152
rect 36728 25100 36780 25152
rect 37924 25236 37976 25288
rect 38568 25304 38620 25356
rect 39304 25304 39356 25356
rect 39396 25304 39448 25356
rect 57244 25347 57296 25356
rect 57244 25313 57253 25347
rect 57253 25313 57287 25347
rect 57287 25313 57296 25347
rect 57244 25304 57296 25313
rect 39120 25279 39172 25288
rect 39120 25245 39129 25279
rect 39129 25245 39163 25279
rect 39163 25245 39172 25279
rect 39120 25236 39172 25245
rect 47860 25168 47912 25220
rect 39396 25100 39448 25152
rect 55680 25143 55732 25152
rect 55680 25109 55689 25143
rect 55689 25109 55723 25143
rect 55723 25109 55732 25143
rect 55680 25100 55732 25109
rect 10614 24998 10666 25050
rect 10678 24998 10730 25050
rect 10742 24998 10794 25050
rect 10806 24998 10858 25050
rect 29878 24998 29930 25050
rect 29942 24998 29994 25050
rect 30006 24998 30058 25050
rect 30070 24998 30122 25050
rect 49142 24998 49194 25050
rect 49206 24998 49258 25050
rect 49270 24998 49322 25050
rect 49334 24998 49386 25050
rect 1492 24939 1544 24948
rect 1492 24905 1501 24939
rect 1501 24905 1535 24939
rect 1535 24905 1544 24939
rect 1492 24896 1544 24905
rect 1584 24896 1636 24948
rect 34336 24896 34388 24948
rect 29644 24828 29696 24880
rect 38016 24871 38068 24880
rect 38016 24837 38025 24871
rect 38025 24837 38059 24871
rect 38059 24837 38068 24871
rect 38016 24828 38068 24837
rect 38476 24828 38528 24880
rect 39948 24828 40000 24880
rect 54392 24896 54444 24948
rect 56692 24896 56744 24948
rect 56784 24896 56836 24948
rect 56968 24939 57020 24948
rect 56968 24905 56977 24939
rect 56977 24905 57011 24939
rect 57011 24905 57020 24939
rect 56968 24896 57020 24905
rect 55680 24828 55732 24880
rect 39396 24760 39448 24812
rect 23572 24735 23624 24744
rect 23572 24701 23581 24735
rect 23581 24701 23615 24735
rect 23615 24701 23624 24735
rect 23572 24692 23624 24701
rect 32312 24692 32364 24744
rect 57888 24692 57940 24744
rect 39856 24624 39908 24676
rect 23480 24599 23532 24608
rect 23480 24565 23489 24599
rect 23489 24565 23523 24599
rect 23523 24565 23532 24599
rect 23480 24556 23532 24565
rect 28908 24599 28960 24608
rect 28908 24565 28917 24599
rect 28917 24565 28951 24599
rect 28951 24565 28960 24599
rect 28908 24556 28960 24565
rect 36728 24599 36780 24608
rect 36728 24565 36737 24599
rect 36737 24565 36771 24599
rect 36771 24565 36780 24599
rect 36728 24556 36780 24565
rect 37280 24599 37332 24608
rect 37280 24565 37289 24599
rect 37289 24565 37323 24599
rect 37323 24565 37332 24599
rect 37280 24556 37332 24565
rect 20246 24454 20298 24506
rect 20310 24454 20362 24506
rect 20374 24454 20426 24506
rect 20438 24454 20490 24506
rect 39510 24454 39562 24506
rect 39574 24454 39626 24506
rect 39638 24454 39690 24506
rect 39702 24454 39754 24506
rect 37556 24352 37608 24404
rect 56876 24395 56928 24404
rect 56876 24361 56885 24395
rect 56885 24361 56919 24395
rect 56919 24361 56928 24395
rect 56876 24352 56928 24361
rect 23112 24216 23164 24268
rect 27436 24216 27488 24268
rect 28448 24216 28500 24268
rect 28908 24216 28960 24268
rect 37740 24259 37792 24268
rect 37740 24225 37749 24259
rect 37749 24225 37783 24259
rect 37783 24225 37792 24259
rect 37740 24216 37792 24225
rect 23480 24148 23532 24200
rect 38476 24191 38528 24200
rect 38476 24157 38485 24191
rect 38485 24157 38519 24191
rect 38519 24157 38528 24191
rect 38476 24148 38528 24157
rect 39212 24216 39264 24268
rect 39304 24148 39356 24200
rect 3516 24080 3568 24132
rect 28356 24123 28408 24132
rect 28356 24089 28365 24123
rect 28365 24089 28399 24123
rect 28399 24089 28408 24123
rect 28356 24080 28408 24089
rect 57888 24216 57940 24268
rect 57796 24148 57848 24200
rect 40684 24055 40736 24064
rect 40684 24021 40693 24055
rect 40693 24021 40727 24055
rect 40727 24021 40736 24055
rect 40684 24012 40736 24021
rect 57980 24055 58032 24064
rect 57980 24021 57989 24055
rect 57989 24021 58023 24055
rect 58023 24021 58032 24055
rect 57980 24012 58032 24021
rect 10614 23910 10666 23962
rect 10678 23910 10730 23962
rect 10742 23910 10794 23962
rect 10806 23910 10858 23962
rect 29878 23910 29930 23962
rect 29942 23910 29994 23962
rect 30006 23910 30058 23962
rect 30070 23910 30122 23962
rect 49142 23910 49194 23962
rect 49206 23910 49258 23962
rect 49270 23910 49322 23962
rect 49334 23910 49386 23962
rect 1492 23851 1544 23860
rect 1492 23817 1501 23851
rect 1501 23817 1535 23851
rect 1535 23817 1544 23851
rect 1492 23808 1544 23817
rect 22744 23808 22796 23860
rect 39212 23851 39264 23860
rect 39212 23817 39221 23851
rect 39221 23817 39255 23851
rect 39255 23817 39264 23851
rect 39212 23808 39264 23817
rect 40684 23808 40736 23860
rect 57980 23808 58032 23860
rect 37740 23740 37792 23792
rect 23480 23672 23532 23724
rect 22560 23647 22612 23656
rect 22560 23613 22569 23647
rect 22569 23613 22603 23647
rect 22603 23613 22612 23647
rect 22560 23604 22612 23613
rect 22744 23647 22796 23656
rect 22744 23613 22753 23647
rect 22753 23613 22787 23647
rect 22787 23613 22796 23647
rect 28448 23672 28500 23724
rect 22744 23604 22796 23613
rect 28540 23647 28592 23656
rect 2136 23511 2188 23520
rect 2136 23477 2145 23511
rect 2145 23477 2179 23511
rect 2179 23477 2188 23511
rect 2136 23468 2188 23477
rect 28540 23613 28549 23647
rect 28549 23613 28583 23647
rect 28583 23613 28592 23647
rect 28540 23604 28592 23613
rect 58164 23647 58216 23656
rect 58164 23613 58173 23647
rect 58173 23613 58207 23647
rect 58207 23613 58216 23647
rect 58164 23604 58216 23613
rect 26240 23536 26292 23588
rect 35900 23536 35952 23588
rect 27436 23468 27488 23520
rect 28264 23511 28316 23520
rect 28264 23477 28273 23511
rect 28273 23477 28307 23511
rect 28307 23477 28316 23511
rect 28264 23468 28316 23477
rect 36728 23468 36780 23520
rect 39948 23468 40000 23520
rect 57796 23468 57848 23520
rect 20246 23366 20298 23418
rect 20310 23366 20362 23418
rect 20374 23366 20426 23418
rect 20438 23366 20490 23418
rect 39510 23366 39562 23418
rect 39574 23366 39626 23418
rect 39638 23366 39690 23418
rect 39702 23366 39754 23418
rect 23112 23264 23164 23316
rect 28540 23264 28592 23316
rect 27436 23239 27488 23248
rect 27436 23205 27445 23239
rect 27445 23205 27479 23239
rect 27479 23205 27488 23239
rect 27436 23196 27488 23205
rect 27620 23239 27672 23248
rect 27620 23205 27629 23239
rect 27629 23205 27663 23239
rect 27663 23205 27672 23239
rect 27620 23196 27672 23205
rect 1400 23171 1452 23180
rect 1400 23137 1409 23171
rect 1409 23137 1443 23171
rect 1443 23137 1452 23171
rect 1400 23128 1452 23137
rect 4160 23128 4212 23180
rect 21180 23128 21232 23180
rect 23112 23128 23164 23180
rect 4896 23103 4948 23112
rect 4896 23069 4905 23103
rect 4905 23069 4939 23103
rect 4939 23069 4948 23103
rect 4896 23060 4948 23069
rect 21548 23035 21600 23044
rect 21548 23001 21557 23035
rect 21557 23001 21591 23035
rect 21591 23001 21600 23035
rect 21548 22992 21600 23001
rect 52460 22992 52512 23044
rect 1676 22924 1728 22976
rect 10614 22822 10666 22874
rect 10678 22822 10730 22874
rect 10742 22822 10794 22874
rect 10806 22822 10858 22874
rect 29878 22822 29930 22874
rect 29942 22822 29994 22874
rect 30006 22822 30058 22874
rect 30070 22822 30122 22874
rect 49142 22822 49194 22874
rect 49206 22822 49258 22874
rect 49270 22822 49322 22874
rect 49334 22822 49386 22874
rect 4160 22763 4212 22772
rect 4160 22729 4169 22763
rect 4169 22729 4203 22763
rect 4203 22729 4212 22763
rect 4160 22720 4212 22729
rect 34612 22720 34664 22772
rect 21180 22559 21232 22568
rect 21180 22525 21189 22559
rect 21189 22525 21223 22559
rect 21223 22525 21232 22559
rect 21180 22516 21232 22525
rect 22744 22516 22796 22568
rect 25964 22516 26016 22568
rect 40224 22720 40276 22772
rect 35992 22516 36044 22568
rect 36544 22516 36596 22568
rect 58164 22559 58216 22568
rect 58164 22525 58173 22559
rect 58173 22525 58207 22559
rect 58207 22525 58216 22559
rect 58164 22516 58216 22525
rect 1400 22491 1452 22500
rect 1400 22457 1409 22491
rect 1409 22457 1443 22491
rect 1443 22457 1452 22491
rect 1400 22448 1452 22457
rect 27436 22380 27488 22432
rect 58256 22380 58308 22432
rect 20246 22278 20298 22330
rect 20310 22278 20362 22330
rect 20374 22278 20426 22330
rect 20438 22278 20490 22330
rect 39510 22278 39562 22330
rect 39574 22278 39626 22330
rect 39638 22278 39690 22330
rect 39702 22278 39754 22330
rect 27804 22176 27856 22228
rect 27252 22083 27304 22092
rect 27252 22049 27261 22083
rect 27261 22049 27295 22083
rect 27295 22049 27304 22083
rect 27252 22040 27304 22049
rect 27436 22083 27488 22092
rect 27436 22049 27445 22083
rect 27445 22049 27479 22083
rect 27479 22049 27488 22083
rect 27436 22040 27488 22049
rect 36268 22083 36320 22092
rect 36268 22049 36277 22083
rect 36277 22049 36311 22083
rect 36311 22049 36320 22083
rect 36268 22040 36320 22049
rect 36544 21904 36596 21956
rect 38108 21904 38160 21956
rect 38568 21904 38620 21956
rect 57336 21947 57388 21956
rect 57336 21913 57345 21947
rect 57345 21913 57379 21947
rect 57379 21913 57388 21947
rect 57336 21904 57388 21913
rect 57888 21904 57940 21956
rect 10614 21734 10666 21786
rect 10678 21734 10730 21786
rect 10742 21734 10794 21786
rect 10806 21734 10858 21786
rect 29878 21734 29930 21786
rect 29942 21734 29994 21786
rect 30006 21734 30058 21786
rect 30070 21734 30122 21786
rect 49142 21734 49194 21786
rect 49206 21734 49258 21786
rect 49270 21734 49322 21786
rect 49334 21734 49386 21786
rect 19800 21675 19852 21684
rect 19800 21641 19809 21675
rect 19809 21641 19843 21675
rect 19843 21641 19852 21675
rect 19800 21632 19852 21641
rect 19984 21632 20036 21684
rect 29460 21675 29512 21684
rect 29460 21641 29469 21675
rect 29469 21641 29503 21675
rect 29503 21641 29512 21675
rect 29460 21632 29512 21641
rect 31024 21632 31076 21684
rect 23756 21564 23808 21616
rect 20076 21496 20128 21548
rect 27252 21428 27304 21480
rect 27620 21428 27672 21480
rect 28172 21360 28224 21412
rect 29460 21428 29512 21480
rect 31392 21471 31444 21480
rect 31392 21437 31401 21471
rect 31401 21437 31435 21471
rect 31435 21437 31444 21471
rect 31392 21428 31444 21437
rect 35900 21471 35952 21480
rect 35900 21437 35909 21471
rect 35909 21437 35943 21471
rect 35943 21437 35952 21471
rect 35900 21428 35952 21437
rect 38384 21496 38436 21548
rect 29276 21292 29328 21344
rect 31300 21360 31352 21412
rect 36544 21360 36596 21412
rect 37832 21428 37884 21480
rect 36084 21335 36136 21344
rect 36084 21301 36093 21335
rect 36093 21301 36127 21335
rect 36127 21301 36136 21335
rect 36084 21292 36136 21301
rect 56784 21292 56836 21344
rect 20246 21190 20298 21242
rect 20310 21190 20362 21242
rect 20374 21190 20426 21242
rect 20438 21190 20490 21242
rect 39510 21190 39562 21242
rect 39574 21190 39626 21242
rect 39638 21190 39690 21242
rect 39702 21190 39754 21242
rect 1492 21131 1544 21140
rect 1492 21097 1501 21131
rect 1501 21097 1535 21131
rect 1535 21097 1544 21131
rect 1492 21088 1544 21097
rect 20076 21131 20128 21140
rect 20076 21097 20085 21131
rect 20085 21097 20119 21131
rect 20119 21097 20128 21131
rect 20076 21088 20128 21097
rect 28172 21088 28224 21140
rect 28540 21020 28592 21072
rect 29276 21063 29328 21072
rect 29276 21029 29285 21063
rect 29285 21029 29319 21063
rect 29319 21029 29328 21063
rect 29276 21020 29328 21029
rect 54576 21088 54628 21140
rect 1584 20995 1636 21004
rect 1584 20961 1593 20995
rect 1593 20961 1627 20995
rect 1627 20961 1636 20995
rect 1584 20952 1636 20961
rect 20076 20952 20128 21004
rect 27436 20952 27488 21004
rect 28172 20995 28224 21004
rect 28172 20961 28181 20995
rect 28181 20961 28215 20995
rect 28215 20961 28224 20995
rect 28172 20952 28224 20961
rect 27712 20927 27764 20936
rect 27712 20893 27721 20927
rect 27721 20893 27755 20927
rect 27755 20893 27764 20927
rect 27712 20884 27764 20893
rect 36084 21020 36136 21072
rect 32220 20995 32272 21004
rect 31116 20884 31168 20936
rect 32220 20961 32229 20995
rect 32229 20961 32263 20995
rect 32263 20961 32272 20995
rect 32220 20952 32272 20961
rect 35992 20995 36044 21004
rect 35992 20961 36001 20995
rect 36001 20961 36035 20995
rect 36035 20961 36044 20995
rect 35992 20952 36044 20961
rect 37832 20995 37884 21004
rect 36084 20927 36136 20936
rect 36084 20893 36093 20927
rect 36093 20893 36127 20927
rect 36127 20893 36136 20927
rect 36084 20884 36136 20893
rect 36636 20884 36688 20936
rect 37096 20884 37148 20936
rect 37832 20961 37841 20995
rect 37841 20961 37875 20995
rect 37875 20961 37884 20995
rect 37832 20952 37884 20961
rect 38016 20995 38068 21004
rect 38016 20961 38025 20995
rect 38025 20961 38059 20995
rect 38059 20961 38068 20995
rect 38016 20952 38068 20961
rect 38844 20995 38896 21004
rect 38844 20961 38853 20995
rect 38853 20961 38887 20995
rect 38887 20961 38896 20995
rect 38844 20952 38896 20961
rect 47216 20952 47268 21004
rect 47400 20884 47452 20936
rect 54392 20952 54444 21004
rect 58164 20995 58216 21004
rect 58164 20961 58173 20995
rect 58173 20961 58207 20995
rect 58207 20961 58216 20995
rect 58164 20952 58216 20961
rect 36268 20816 36320 20868
rect 57336 20816 57388 20868
rect 47216 20791 47268 20800
rect 47216 20757 47225 20791
rect 47225 20757 47259 20791
rect 47259 20757 47268 20791
rect 47216 20748 47268 20757
rect 47768 20791 47820 20800
rect 47768 20757 47777 20791
rect 47777 20757 47811 20791
rect 47811 20757 47820 20791
rect 47768 20748 47820 20757
rect 10614 20646 10666 20698
rect 10678 20646 10730 20698
rect 10742 20646 10794 20698
rect 10806 20646 10858 20698
rect 29878 20646 29930 20698
rect 29942 20646 29994 20698
rect 30006 20646 30058 20698
rect 30070 20646 30122 20698
rect 49142 20646 49194 20698
rect 49206 20646 49258 20698
rect 49270 20646 49322 20698
rect 49334 20646 49386 20698
rect 4528 20544 4580 20596
rect 38384 20587 38436 20596
rect 38384 20553 38393 20587
rect 38393 20553 38427 20587
rect 38427 20553 38436 20587
rect 38384 20544 38436 20553
rect 47400 20587 47452 20596
rect 47400 20553 47409 20587
rect 47409 20553 47443 20587
rect 47443 20553 47452 20587
rect 47400 20544 47452 20553
rect 1400 20383 1452 20392
rect 1400 20349 1409 20383
rect 1409 20349 1443 20383
rect 1443 20349 1452 20383
rect 1400 20340 1452 20349
rect 21916 20340 21968 20392
rect 22560 20340 22612 20392
rect 23112 20383 23164 20392
rect 23112 20349 23121 20383
rect 23121 20349 23155 20383
rect 23155 20349 23164 20383
rect 23112 20340 23164 20349
rect 31300 20340 31352 20392
rect 32220 20340 32272 20392
rect 32680 20340 32732 20392
rect 36544 20383 36596 20392
rect 36544 20349 36553 20383
rect 36553 20349 36587 20383
rect 36587 20349 36596 20383
rect 36544 20340 36596 20349
rect 37096 20340 37148 20392
rect 31944 20272 31996 20324
rect 2688 20247 2740 20256
rect 2688 20213 2697 20247
rect 2697 20213 2731 20247
rect 2731 20213 2740 20247
rect 2688 20204 2740 20213
rect 23296 20247 23348 20256
rect 23296 20213 23305 20247
rect 23305 20213 23339 20247
rect 23339 20213 23348 20247
rect 23296 20204 23348 20213
rect 36360 20247 36412 20256
rect 36360 20213 36369 20247
rect 36369 20213 36403 20247
rect 36403 20213 36412 20247
rect 36360 20204 36412 20213
rect 38936 20247 38988 20256
rect 38936 20213 38945 20247
rect 38945 20213 38979 20247
rect 38979 20213 38988 20247
rect 38936 20204 38988 20213
rect 20246 20102 20298 20154
rect 20310 20102 20362 20154
rect 20374 20102 20426 20154
rect 20438 20102 20490 20154
rect 39510 20102 39562 20154
rect 39574 20102 39626 20154
rect 39638 20102 39690 20154
rect 39702 20102 39754 20154
rect 1584 20000 1636 20052
rect 2504 20000 2556 20052
rect 15844 20000 15896 20052
rect 21916 20043 21968 20052
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 2688 19864 2740 19916
rect 8760 19864 8812 19916
rect 16212 19796 16264 19848
rect 21916 20009 21925 20043
rect 21925 20009 21959 20043
rect 21959 20009 21968 20043
rect 21916 20000 21968 20009
rect 23296 20000 23348 20052
rect 57796 20000 57848 20052
rect 32680 19975 32732 19984
rect 32680 19941 32689 19975
rect 32689 19941 32723 19975
rect 32723 19941 32732 19975
rect 32680 19932 32732 19941
rect 21824 19907 21876 19916
rect 21824 19873 21833 19907
rect 21833 19873 21867 19907
rect 21867 19873 21876 19907
rect 21824 19864 21876 19873
rect 31116 19907 31168 19916
rect 31116 19873 31125 19907
rect 31125 19873 31159 19907
rect 31159 19873 31168 19907
rect 31116 19864 31168 19873
rect 31392 19907 31444 19916
rect 31392 19873 31401 19907
rect 31401 19873 31435 19907
rect 31435 19873 31444 19907
rect 31392 19864 31444 19873
rect 32220 19864 32272 19916
rect 32404 19864 32456 19916
rect 35808 19864 35860 19916
rect 36544 19864 36596 19916
rect 38016 19864 38068 19916
rect 54944 19796 54996 19848
rect 3976 19703 4028 19712
rect 3976 19669 3985 19703
rect 3985 19669 4019 19703
rect 4019 19669 4028 19703
rect 3976 19660 4028 19669
rect 31484 19728 31536 19780
rect 58164 19771 58216 19780
rect 58164 19737 58173 19771
rect 58173 19737 58207 19771
rect 58207 19737 58216 19771
rect 58164 19728 58216 19737
rect 19340 19660 19392 19712
rect 35808 19703 35860 19712
rect 35808 19669 35817 19703
rect 35817 19669 35851 19703
rect 35851 19669 35860 19703
rect 35808 19660 35860 19669
rect 10614 19558 10666 19610
rect 10678 19558 10730 19610
rect 10742 19558 10794 19610
rect 10806 19558 10858 19610
rect 29878 19558 29930 19610
rect 29942 19558 29994 19610
rect 30006 19558 30058 19610
rect 30070 19558 30122 19610
rect 49142 19558 49194 19610
rect 49206 19558 49258 19610
rect 49270 19558 49322 19610
rect 49334 19558 49386 19610
rect 2320 19499 2372 19508
rect 2320 19465 2329 19499
rect 2329 19465 2363 19499
rect 2363 19465 2372 19499
rect 2320 19456 2372 19465
rect 3976 19456 4028 19508
rect 25688 19456 25740 19508
rect 7012 19388 7064 19440
rect 35808 19388 35860 19440
rect 16212 19363 16264 19372
rect 16212 19329 16221 19363
rect 16221 19329 16255 19363
rect 16255 19329 16264 19363
rect 16212 19320 16264 19329
rect 1400 19295 1452 19304
rect 1400 19261 1409 19295
rect 1409 19261 1443 19295
rect 1443 19261 1452 19295
rect 1400 19252 1452 19261
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 8668 19295 8720 19304
rect 8668 19261 8677 19295
rect 8677 19261 8711 19295
rect 8711 19261 8720 19295
rect 8668 19252 8720 19261
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 58164 19227 58216 19236
rect 58164 19193 58173 19227
rect 58173 19193 58207 19227
rect 58207 19193 58216 19227
rect 58164 19184 58216 19193
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 32220 19116 32272 19168
rect 45744 19116 45796 19168
rect 57336 19159 57388 19168
rect 57336 19125 57345 19159
rect 57345 19125 57379 19159
rect 57379 19125 57388 19159
rect 57336 19116 57388 19125
rect 20246 19014 20298 19066
rect 20310 19014 20362 19066
rect 20374 19014 20426 19066
rect 20438 19014 20490 19066
rect 39510 19014 39562 19066
rect 39574 19014 39626 19066
rect 39638 19014 39690 19066
rect 39702 19014 39754 19066
rect 1400 18955 1452 18964
rect 1400 18921 1409 18955
rect 1409 18921 1443 18955
rect 1443 18921 1452 18955
rect 1400 18912 1452 18921
rect 1584 18912 1636 18964
rect 26608 18912 26660 18964
rect 25780 18776 25832 18828
rect 26792 18776 26844 18828
rect 27068 18776 27120 18828
rect 27896 18819 27948 18828
rect 27896 18785 27905 18819
rect 27905 18785 27939 18819
rect 27939 18785 27948 18819
rect 27896 18776 27948 18785
rect 2504 18708 2556 18760
rect 4160 18708 4212 18760
rect 44456 18708 44508 18760
rect 34888 18640 34940 18692
rect 42340 18640 42392 18692
rect 57152 18640 57204 18692
rect 2044 18572 2096 18624
rect 10614 18470 10666 18522
rect 10678 18470 10730 18522
rect 10742 18470 10794 18522
rect 10806 18470 10858 18522
rect 29878 18470 29930 18522
rect 29942 18470 29994 18522
rect 30006 18470 30058 18522
rect 30070 18470 30122 18522
rect 49142 18470 49194 18522
rect 49206 18470 49258 18522
rect 49270 18470 49322 18522
rect 49334 18470 49386 18522
rect 2228 18368 2280 18420
rect 2504 18368 2556 18420
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 20246 17926 20298 17978
rect 20310 17926 20362 17978
rect 20374 17926 20426 17978
rect 20438 17926 20490 17978
rect 39510 17926 39562 17978
rect 39574 17926 39626 17978
rect 39638 17926 39690 17978
rect 39702 17926 39754 17978
rect 27068 17867 27120 17876
rect 27068 17833 27077 17867
rect 27077 17833 27111 17867
rect 27111 17833 27120 17867
rect 27068 17824 27120 17833
rect 27620 17824 27672 17876
rect 25412 17756 25464 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 2228 17688 2280 17740
rect 26608 17620 26660 17672
rect 28724 17688 28776 17740
rect 58164 17731 58216 17740
rect 58164 17697 58173 17731
rect 58173 17697 58207 17731
rect 58207 17697 58216 17731
rect 58164 17688 58216 17697
rect 36268 17620 36320 17672
rect 54392 17620 54444 17672
rect 2228 17527 2280 17536
rect 2228 17493 2237 17527
rect 2237 17493 2271 17527
rect 2271 17493 2280 17527
rect 2228 17484 2280 17493
rect 54944 17484 54996 17536
rect 10614 17382 10666 17434
rect 10678 17382 10730 17434
rect 10742 17382 10794 17434
rect 10806 17382 10858 17434
rect 29878 17382 29930 17434
rect 29942 17382 29994 17434
rect 30006 17382 30058 17434
rect 30070 17382 30122 17434
rect 49142 17382 49194 17434
rect 49206 17382 49258 17434
rect 49270 17382 49322 17434
rect 49334 17382 49386 17434
rect 25412 17323 25464 17332
rect 25412 17289 25421 17323
rect 25421 17289 25455 17323
rect 25455 17289 25464 17323
rect 25412 17280 25464 17289
rect 54392 17323 54444 17332
rect 54392 17289 54401 17323
rect 54401 17289 54435 17323
rect 54435 17289 54444 17323
rect 54392 17280 54444 17289
rect 19340 17144 19392 17196
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 25320 17119 25372 17128
rect 25320 17085 25329 17119
rect 25329 17085 25363 17119
rect 25363 17085 25372 17119
rect 25320 17076 25372 17085
rect 26608 17119 26660 17128
rect 26608 17085 26617 17119
rect 26617 17085 26651 17119
rect 26651 17085 26660 17119
rect 26608 17076 26660 17085
rect 36268 17119 36320 17128
rect 36268 17085 36277 17119
rect 36277 17085 36311 17119
rect 36311 17085 36320 17119
rect 36268 17076 36320 17085
rect 57888 17119 57940 17128
rect 57888 17085 57897 17119
rect 57897 17085 57931 17119
rect 57931 17085 57940 17119
rect 57888 17076 57940 17085
rect 36452 17008 36504 17060
rect 37648 17008 37700 17060
rect 58072 17051 58124 17060
rect 58072 17017 58081 17051
rect 58081 17017 58115 17051
rect 58115 17017 58124 17051
rect 58072 17008 58124 17017
rect 8484 16940 8536 16992
rect 20246 16838 20298 16890
rect 20310 16838 20362 16890
rect 20374 16838 20426 16890
rect 20438 16838 20490 16890
rect 39510 16838 39562 16890
rect 39574 16838 39626 16890
rect 39638 16838 39690 16890
rect 39702 16838 39754 16890
rect 10324 16779 10376 16788
rect 10324 16745 10333 16779
rect 10333 16745 10367 16779
rect 10367 16745 10376 16779
rect 10324 16736 10376 16745
rect 21364 16736 21416 16788
rect 1400 16600 1452 16652
rect 8484 16600 8536 16652
rect 21180 16600 21232 16652
rect 22744 16736 22796 16788
rect 14372 16532 14424 16584
rect 22744 16643 22796 16652
rect 22744 16609 22753 16643
rect 22753 16609 22787 16643
rect 22787 16609 22796 16643
rect 22744 16600 22796 16609
rect 25412 16600 25464 16652
rect 26792 16643 26844 16652
rect 26792 16609 26801 16643
rect 26801 16609 26835 16643
rect 26835 16609 26844 16643
rect 26792 16600 26844 16609
rect 29460 16668 29512 16720
rect 29368 16643 29420 16652
rect 29368 16609 29377 16643
rect 29377 16609 29411 16643
rect 29411 16609 29420 16643
rect 29368 16600 29420 16609
rect 37096 16643 37148 16652
rect 37096 16609 37105 16643
rect 37105 16609 37139 16643
rect 37139 16609 37148 16643
rect 37096 16600 37148 16609
rect 13544 16464 13596 16516
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 21180 16396 21232 16448
rect 25320 16464 25372 16516
rect 23296 16396 23348 16448
rect 24400 16396 24452 16448
rect 26516 16396 26568 16448
rect 26884 16396 26936 16448
rect 29276 16464 29328 16516
rect 37464 16532 37516 16584
rect 37556 16532 37608 16584
rect 57888 16668 57940 16720
rect 57980 16643 58032 16652
rect 40868 16464 40920 16516
rect 29552 16396 29604 16448
rect 38200 16439 38252 16448
rect 38200 16405 38209 16439
rect 38209 16405 38243 16439
rect 38243 16405 38252 16439
rect 38200 16396 38252 16405
rect 44548 16439 44600 16448
rect 44548 16405 44557 16439
rect 44557 16405 44591 16439
rect 44591 16405 44600 16439
rect 44548 16396 44600 16405
rect 57980 16609 57989 16643
rect 57989 16609 58023 16643
rect 58023 16609 58032 16643
rect 57980 16600 58032 16609
rect 58164 16507 58216 16516
rect 58164 16473 58173 16507
rect 58173 16473 58207 16507
rect 58207 16473 58216 16507
rect 58164 16464 58216 16473
rect 57704 16396 57756 16448
rect 10614 16294 10666 16346
rect 10678 16294 10730 16346
rect 10742 16294 10794 16346
rect 10806 16294 10858 16346
rect 29878 16294 29930 16346
rect 29942 16294 29994 16346
rect 30006 16294 30058 16346
rect 30070 16294 30122 16346
rect 49142 16294 49194 16346
rect 49206 16294 49258 16346
rect 49270 16294 49322 16346
rect 49334 16294 49386 16346
rect 1400 16235 1452 16244
rect 1400 16201 1409 16235
rect 1409 16201 1443 16235
rect 1443 16201 1452 16235
rect 1400 16192 1452 16201
rect 1584 16192 1636 16244
rect 29736 16192 29788 16244
rect 30196 16192 30248 16244
rect 37096 16192 37148 16244
rect 17868 16124 17920 16176
rect 25688 16124 25740 16176
rect 29184 16124 29236 16176
rect 21088 16099 21140 16108
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 57336 16124 57388 16176
rect 37556 16056 37608 16108
rect 38200 16056 38252 16108
rect 40868 16099 40920 16108
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 8300 15920 8352 15972
rect 18788 15988 18840 16040
rect 21364 16031 21416 16040
rect 21364 15997 21373 16031
rect 21373 15997 21407 16031
rect 21407 15997 21416 16031
rect 21364 15988 21416 15997
rect 23204 16031 23256 16040
rect 23204 15997 23213 16031
rect 23213 15997 23247 16031
rect 23247 15997 23256 16031
rect 23204 15988 23256 15997
rect 15476 15920 15528 15972
rect 22008 15920 22060 15972
rect 25504 15988 25556 16040
rect 29092 16031 29144 16040
rect 29092 15997 29101 16031
rect 29101 15997 29135 16031
rect 29135 15997 29144 16031
rect 29092 15988 29144 15997
rect 29276 16031 29328 16040
rect 29276 15997 29285 16031
rect 29285 15997 29319 16031
rect 29319 15997 29328 16031
rect 29276 15988 29328 15997
rect 29552 15988 29604 16040
rect 35992 16031 36044 16040
rect 35992 15997 36001 16031
rect 36001 15997 36035 16031
rect 36035 15997 36044 16031
rect 35992 15988 36044 15997
rect 36268 15988 36320 16040
rect 40868 16065 40877 16099
rect 40877 16065 40911 16099
rect 40911 16065 40920 16099
rect 40868 16056 40920 16065
rect 43536 16099 43588 16108
rect 43536 16065 43545 16099
rect 43545 16065 43579 16099
rect 43579 16065 43588 16099
rect 43536 16056 43588 16065
rect 25412 15852 25464 15904
rect 26792 15920 26844 15972
rect 30196 15920 30248 15972
rect 28908 15852 28960 15904
rect 29092 15852 29144 15904
rect 29736 15852 29788 15904
rect 37096 15920 37148 15972
rect 38384 15920 38436 15972
rect 41144 15988 41196 16040
rect 43628 16031 43680 16040
rect 43628 15997 43637 16031
rect 43637 15997 43671 16031
rect 43671 15997 43680 16031
rect 43628 15988 43680 15997
rect 44548 16031 44600 16040
rect 44548 15997 44557 16031
rect 44557 15997 44591 16031
rect 44591 15997 44600 16031
rect 44548 15988 44600 15997
rect 35900 15895 35952 15904
rect 35900 15861 35909 15895
rect 35909 15861 35943 15895
rect 35943 15861 35952 15895
rect 35900 15852 35952 15861
rect 39856 15852 39908 15904
rect 57980 15920 58032 15972
rect 45836 15852 45888 15904
rect 20246 15750 20298 15802
rect 20310 15750 20362 15802
rect 20374 15750 20426 15802
rect 20438 15750 20490 15802
rect 39510 15750 39562 15802
rect 39574 15750 39626 15802
rect 39638 15750 39690 15802
rect 39702 15750 39754 15802
rect 1584 15691 1636 15700
rect 1584 15657 1593 15691
rect 1593 15657 1627 15691
rect 1627 15657 1636 15691
rect 1584 15648 1636 15657
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 18880 15648 18932 15700
rect 21180 15648 21232 15700
rect 22008 15691 22060 15700
rect 22008 15657 22017 15691
rect 22017 15657 22051 15691
rect 22051 15657 22060 15691
rect 22008 15648 22060 15657
rect 29276 15648 29328 15700
rect 35992 15648 36044 15700
rect 37096 15691 37148 15700
rect 37096 15657 37105 15691
rect 37105 15657 37139 15691
rect 37139 15657 37148 15691
rect 37096 15648 37148 15657
rect 37832 15648 37884 15700
rect 17868 15555 17920 15564
rect 17868 15521 17877 15555
rect 17877 15521 17911 15555
rect 17911 15521 17920 15555
rect 17868 15512 17920 15521
rect 18788 15555 18840 15564
rect 18788 15521 18797 15555
rect 18797 15521 18831 15555
rect 18831 15521 18840 15555
rect 18788 15512 18840 15521
rect 10324 15444 10376 15496
rect 19984 15444 20036 15496
rect 21180 15444 21232 15496
rect 21364 15512 21416 15564
rect 24400 15512 24452 15564
rect 28356 15512 28408 15564
rect 35900 15580 35952 15632
rect 23664 15444 23716 15496
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 25412 15444 25464 15453
rect 25504 15444 25556 15496
rect 38108 15580 38160 15632
rect 39856 15512 39908 15564
rect 44548 15512 44600 15564
rect 33232 15487 33284 15496
rect 33232 15453 33241 15487
rect 33241 15453 33275 15487
rect 33275 15453 33284 15487
rect 33232 15444 33284 15453
rect 37280 15444 37332 15496
rect 38660 15487 38712 15496
rect 38660 15453 38669 15487
rect 38669 15453 38703 15487
rect 38703 15453 38712 15487
rect 38660 15444 38712 15453
rect 41420 15487 41472 15496
rect 41420 15453 41429 15487
rect 41429 15453 41463 15487
rect 41463 15453 41472 15487
rect 41420 15444 41472 15453
rect 18972 15351 19024 15360
rect 18972 15317 18981 15351
rect 18981 15317 19015 15351
rect 19015 15317 19024 15351
rect 18972 15308 19024 15317
rect 10614 15206 10666 15258
rect 10678 15206 10730 15258
rect 10742 15206 10794 15258
rect 10806 15206 10858 15258
rect 29878 15206 29930 15258
rect 29942 15206 29994 15258
rect 30006 15206 30058 15258
rect 30070 15206 30122 15258
rect 49142 15206 49194 15258
rect 49206 15206 49258 15258
rect 49270 15206 49322 15258
rect 49334 15206 49386 15258
rect 1400 15147 1452 15156
rect 1400 15113 1409 15147
rect 1409 15113 1443 15147
rect 1443 15113 1452 15147
rect 1400 15104 1452 15113
rect 18880 15147 18932 15156
rect 18880 15113 18889 15147
rect 18889 15113 18923 15147
rect 18923 15113 18932 15147
rect 18880 15104 18932 15113
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 18052 14943 18104 14952
rect 18052 14909 18061 14943
rect 18061 14909 18095 14943
rect 18095 14909 18104 14943
rect 18052 14900 18104 14909
rect 36820 14943 36872 14952
rect 36820 14909 36829 14943
rect 36829 14909 36863 14943
rect 36863 14909 36872 14943
rect 36820 14900 36872 14909
rect 38108 14900 38160 14952
rect 58164 14943 58216 14952
rect 58164 14909 58173 14943
rect 58173 14909 58207 14943
rect 58207 14909 58216 14943
rect 58164 14900 58216 14909
rect 35440 14832 35492 14884
rect 57980 14807 58032 14816
rect 57980 14773 57989 14807
rect 57989 14773 58023 14807
rect 58023 14773 58032 14807
rect 57980 14764 58032 14773
rect 20246 14662 20298 14714
rect 20310 14662 20362 14714
rect 20374 14662 20426 14714
rect 20438 14662 20490 14714
rect 39510 14662 39562 14714
rect 39574 14662 39626 14714
rect 39638 14662 39690 14714
rect 39702 14662 39754 14714
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 57980 14560 58032 14612
rect 23664 14535 23716 14544
rect 23664 14501 23673 14535
rect 23673 14501 23707 14535
rect 23707 14501 23716 14535
rect 23664 14492 23716 14501
rect 52460 14535 52512 14544
rect 52460 14501 52469 14535
rect 52469 14501 52503 14535
rect 52503 14501 52512 14535
rect 52460 14492 52512 14501
rect 22560 14424 22612 14476
rect 37004 14424 37056 14476
rect 54392 14492 54444 14544
rect 53104 14467 53156 14476
rect 53104 14433 53113 14467
rect 53113 14433 53147 14467
rect 53147 14433 53156 14467
rect 53104 14424 53156 14433
rect 58164 14467 58216 14476
rect 58164 14433 58173 14467
rect 58173 14433 58207 14467
rect 58207 14433 58216 14467
rect 58164 14424 58216 14433
rect 17684 14288 17736 14340
rect 18052 14288 18104 14340
rect 23204 14288 23256 14340
rect 36820 14288 36872 14340
rect 13728 14220 13780 14272
rect 23572 14263 23624 14272
rect 23572 14229 23581 14263
rect 23581 14229 23615 14263
rect 23615 14229 23624 14263
rect 23572 14220 23624 14229
rect 54392 14220 54444 14272
rect 56324 14220 56376 14272
rect 10614 14118 10666 14170
rect 10678 14118 10730 14170
rect 10742 14118 10794 14170
rect 10806 14118 10858 14170
rect 29878 14118 29930 14170
rect 29942 14118 29994 14170
rect 30006 14118 30058 14170
rect 30070 14118 30122 14170
rect 49142 14118 49194 14170
rect 49206 14118 49258 14170
rect 49270 14118 49322 14170
rect 49334 14118 49386 14170
rect 1400 13855 1452 13864
rect 1400 13821 1409 13855
rect 1409 13821 1443 13855
rect 1443 13821 1452 13855
rect 1400 13812 1452 13821
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 13728 13855 13780 13864
rect 13728 13821 13737 13855
rect 13737 13821 13771 13855
rect 13771 13821 13780 13855
rect 13728 13812 13780 13821
rect 21088 13812 21140 13864
rect 22836 13855 22888 13864
rect 22836 13821 22845 13855
rect 22845 13821 22879 13855
rect 22879 13821 22888 13855
rect 22836 13812 22888 13821
rect 23572 13812 23624 13864
rect 34704 13812 34756 13864
rect 2136 13744 2188 13796
rect 13820 13787 13872 13796
rect 13820 13753 13829 13787
rect 13829 13753 13863 13787
rect 13863 13753 13872 13787
rect 13820 13744 13872 13753
rect 19892 13744 19944 13796
rect 2412 13676 2464 13728
rect 23572 13719 23624 13728
rect 23572 13685 23581 13719
rect 23581 13685 23615 13719
rect 23615 13685 23624 13719
rect 34612 13719 34664 13728
rect 23572 13676 23624 13685
rect 34612 13685 34621 13719
rect 34621 13685 34655 13719
rect 34655 13685 34664 13719
rect 34612 13676 34664 13685
rect 55128 13676 55180 13728
rect 20246 13574 20298 13626
rect 20310 13574 20362 13626
rect 20374 13574 20426 13626
rect 20438 13574 20490 13626
rect 39510 13574 39562 13626
rect 39574 13574 39626 13626
rect 39638 13574 39690 13626
rect 39702 13574 39754 13626
rect 2412 13515 2464 13524
rect 2412 13481 2421 13515
rect 2421 13481 2455 13515
rect 2455 13481 2464 13515
rect 2412 13472 2464 13481
rect 1584 13404 1636 13456
rect 2504 13404 2556 13456
rect 1676 13132 1728 13184
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 15568 13472 15620 13524
rect 10600 13404 10652 13456
rect 10508 13379 10560 13388
rect 10508 13345 10517 13379
rect 10517 13345 10551 13379
rect 10551 13345 10560 13379
rect 10508 13336 10560 13345
rect 2412 13200 2464 13252
rect 11888 13336 11940 13388
rect 13728 13404 13780 13456
rect 11060 13268 11112 13320
rect 18972 13336 19024 13388
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 10614 13030 10666 13082
rect 10678 13030 10730 13082
rect 10742 13030 10794 13082
rect 10806 13030 10858 13082
rect 29878 13030 29930 13082
rect 29942 13030 29994 13082
rect 30006 13030 30058 13082
rect 30070 13030 30122 13082
rect 49142 13030 49194 13082
rect 49206 13030 49258 13082
rect 49270 13030 49322 13082
rect 49334 13030 49386 13082
rect 10508 12928 10560 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 57888 12792 57940 12844
rect 1860 12588 1912 12640
rect 38936 12588 38988 12640
rect 20246 12486 20298 12538
rect 20310 12486 20362 12538
rect 20374 12486 20426 12538
rect 20438 12486 20490 12538
rect 39510 12486 39562 12538
rect 39574 12486 39626 12538
rect 39638 12486 39690 12538
rect 39702 12486 39754 12538
rect 58164 12291 58216 12300
rect 58164 12257 58173 12291
rect 58173 12257 58207 12291
rect 58207 12257 58216 12291
rect 58164 12248 58216 12257
rect 2228 12180 2280 12232
rect 36176 12180 36228 12232
rect 11888 12112 11940 12164
rect 10614 11942 10666 11994
rect 10678 11942 10730 11994
rect 10742 11942 10794 11994
rect 10806 11942 10858 11994
rect 29878 11942 29930 11994
rect 29942 11942 29994 11994
rect 30006 11942 30058 11994
rect 30070 11942 30122 11994
rect 49142 11942 49194 11994
rect 49206 11942 49258 11994
rect 49270 11942 49322 11994
rect 49334 11942 49386 11994
rect 1400 11611 1452 11620
rect 1400 11577 1409 11611
rect 1409 11577 1443 11611
rect 1443 11577 1452 11611
rect 1400 11568 1452 11577
rect 2228 11611 2280 11620
rect 2228 11577 2237 11611
rect 2237 11577 2271 11611
rect 2271 11577 2280 11611
rect 2228 11568 2280 11577
rect 57888 11568 57940 11620
rect 58164 11611 58216 11620
rect 58164 11577 58173 11611
rect 58173 11577 58207 11611
rect 58207 11577 58216 11611
rect 58164 11568 58216 11577
rect 20246 11398 20298 11450
rect 20310 11398 20362 11450
rect 20374 11398 20426 11450
rect 20438 11398 20490 11450
rect 39510 11398 39562 11450
rect 39574 11398 39626 11450
rect 39638 11398 39690 11450
rect 39702 11398 39754 11450
rect 57888 11339 57940 11348
rect 57888 11305 57897 11339
rect 57897 11305 57931 11339
rect 57931 11305 57940 11339
rect 57888 11296 57940 11305
rect 58256 11228 58308 11280
rect 41420 11160 41472 11212
rect 56416 11092 56468 11144
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 28540 10956 28592 11008
rect 10614 10854 10666 10906
rect 10678 10854 10730 10906
rect 10742 10854 10794 10906
rect 10806 10854 10858 10906
rect 29878 10854 29930 10906
rect 29942 10854 29994 10906
rect 30006 10854 30058 10906
rect 30070 10854 30122 10906
rect 49142 10854 49194 10906
rect 49206 10854 49258 10906
rect 49270 10854 49322 10906
rect 49334 10854 49386 10906
rect 23296 10752 23348 10804
rect 2228 10412 2280 10464
rect 30932 10548 30984 10600
rect 25044 10480 25096 10532
rect 56416 10412 56468 10464
rect 20246 10310 20298 10362
rect 20310 10310 20362 10362
rect 20374 10310 20426 10362
rect 20438 10310 20490 10362
rect 39510 10310 39562 10362
rect 39574 10310 39626 10362
rect 39638 10310 39690 10362
rect 39702 10310 39754 10362
rect 57796 10140 57848 10192
rect 58164 10183 58216 10192
rect 58164 10149 58173 10183
rect 58173 10149 58207 10183
rect 58207 10149 58216 10183
rect 58164 10140 58216 10149
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 33324 9868 33376 9920
rect 42340 9868 42392 9920
rect 10614 9766 10666 9818
rect 10678 9766 10730 9818
rect 10742 9766 10794 9818
rect 10806 9766 10858 9818
rect 29878 9766 29930 9818
rect 29942 9766 29994 9818
rect 30006 9766 30058 9818
rect 30070 9766 30122 9818
rect 49142 9766 49194 9818
rect 49206 9766 49258 9818
rect 49270 9766 49322 9818
rect 49334 9766 49386 9818
rect 19064 9664 19116 9716
rect 49976 9664 50028 9716
rect 30932 9596 30984 9648
rect 1492 9503 1544 9512
rect 1492 9469 1501 9503
rect 1501 9469 1535 9503
rect 1535 9469 1544 9503
rect 1492 9460 1544 9469
rect 58164 9571 58216 9580
rect 58164 9537 58173 9571
rect 58173 9537 58207 9571
rect 58207 9537 58216 9571
rect 58164 9528 58216 9537
rect 35348 9503 35400 9512
rect 35348 9469 35357 9503
rect 35357 9469 35391 9503
rect 35391 9469 35400 9503
rect 35348 9460 35400 9469
rect 21824 9324 21876 9376
rect 20246 9222 20298 9274
rect 20310 9222 20362 9274
rect 20374 9222 20426 9274
rect 20438 9222 20490 9274
rect 39510 9222 39562 9274
rect 39574 9222 39626 9274
rect 39638 9222 39690 9274
rect 39702 9222 39754 9274
rect 9220 9052 9272 9104
rect 1400 8891 1452 8900
rect 1400 8857 1409 8891
rect 1409 8857 1443 8891
rect 1443 8857 1452 8891
rect 1400 8848 1452 8857
rect 10614 8678 10666 8730
rect 10678 8678 10730 8730
rect 10742 8678 10794 8730
rect 10806 8678 10858 8730
rect 29878 8678 29930 8730
rect 29942 8678 29994 8730
rect 30006 8678 30058 8730
rect 30070 8678 30122 8730
rect 49142 8678 49194 8730
rect 49206 8678 49258 8730
rect 49270 8678 49322 8730
rect 49334 8678 49386 8730
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 9588 8576 9640 8628
rect 26516 8619 26568 8628
rect 1492 8279 1544 8288
rect 1492 8245 1501 8279
rect 1501 8245 1535 8279
rect 1535 8245 1544 8279
rect 1492 8236 1544 8245
rect 2504 8236 2556 8288
rect 13728 8440 13780 8492
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 26516 8585 26525 8619
rect 26525 8585 26559 8619
rect 26559 8585 26568 8619
rect 26516 8576 26568 8585
rect 41788 8372 41840 8424
rect 25596 8304 25648 8356
rect 38660 8304 38712 8356
rect 58164 8347 58216 8356
rect 58164 8313 58173 8347
rect 58173 8313 58207 8347
rect 58207 8313 58216 8347
rect 58164 8304 58216 8313
rect 9680 8279 9732 8288
rect 9680 8245 9689 8279
rect 9689 8245 9723 8279
rect 9723 8245 9732 8279
rect 9680 8236 9732 8245
rect 20246 8134 20298 8186
rect 20310 8134 20362 8186
rect 20374 8134 20426 8186
rect 20438 8134 20490 8186
rect 39510 8134 39562 8186
rect 39574 8134 39626 8186
rect 39638 8134 39690 8186
rect 39702 8134 39754 8186
rect 25596 8032 25648 8084
rect 25780 7939 25832 7948
rect 25780 7905 25789 7939
rect 25789 7905 25823 7939
rect 25823 7905 25832 7939
rect 25780 7896 25832 7905
rect 26516 7896 26568 7948
rect 27896 7964 27948 8016
rect 20628 7828 20680 7880
rect 10614 7590 10666 7642
rect 10678 7590 10730 7642
rect 10742 7590 10794 7642
rect 10806 7590 10858 7642
rect 29878 7590 29930 7642
rect 29942 7590 29994 7642
rect 30006 7590 30058 7642
rect 30070 7590 30122 7642
rect 49142 7590 49194 7642
rect 49206 7590 49258 7642
rect 49270 7590 49322 7642
rect 49334 7590 49386 7642
rect 26516 7488 26568 7540
rect 27896 7488 27948 7540
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 58164 7327 58216 7336
rect 58164 7293 58173 7327
rect 58173 7293 58207 7327
rect 58207 7293 58216 7327
rect 58164 7284 58216 7293
rect 57888 7216 57940 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 57980 7191 58032 7200
rect 57980 7157 57989 7191
rect 57989 7157 58023 7191
rect 58023 7157 58032 7191
rect 57980 7148 58032 7157
rect 20246 7046 20298 7098
rect 20310 7046 20362 7098
rect 20374 7046 20426 7098
rect 20438 7046 20490 7098
rect 39510 7046 39562 7098
rect 39574 7046 39626 7098
rect 39638 7046 39690 7098
rect 39702 7046 39754 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 1584 6944 1636 6996
rect 2504 6876 2556 6928
rect 57888 6919 57940 6928
rect 57888 6885 57897 6919
rect 57897 6885 57931 6919
rect 57931 6885 57940 6919
rect 57888 6876 57940 6885
rect 1676 6740 1728 6792
rect 57980 6808 58032 6860
rect 58072 6851 58124 6860
rect 58072 6817 58081 6851
rect 58081 6817 58115 6851
rect 58115 6817 58124 6851
rect 58072 6808 58124 6817
rect 57520 6672 57572 6724
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 54024 6647 54076 6656
rect 54024 6613 54033 6647
rect 54033 6613 54067 6647
rect 54067 6613 54076 6647
rect 54024 6604 54076 6613
rect 10614 6502 10666 6554
rect 10678 6502 10730 6554
rect 10742 6502 10794 6554
rect 10806 6502 10858 6554
rect 29878 6502 29930 6554
rect 29942 6502 29994 6554
rect 30006 6502 30058 6554
rect 30070 6502 30122 6554
rect 49142 6502 49194 6554
rect 49206 6502 49258 6554
rect 49270 6502 49322 6554
rect 49334 6502 49386 6554
rect 1584 6239 1636 6248
rect 1584 6205 1593 6239
rect 1593 6205 1627 6239
rect 1627 6205 1636 6239
rect 1584 6196 1636 6205
rect 1400 6171 1452 6180
rect 1400 6137 1409 6171
rect 1409 6137 1443 6171
rect 1443 6137 1452 6171
rect 1400 6128 1452 6137
rect 57704 6103 57756 6112
rect 57704 6069 57713 6103
rect 57713 6069 57747 6103
rect 57747 6069 57756 6103
rect 57704 6060 57756 6069
rect 20246 5958 20298 6010
rect 20310 5958 20362 6010
rect 20374 5958 20426 6010
rect 20438 5958 20490 6010
rect 39510 5958 39562 6010
rect 39574 5958 39626 6010
rect 39638 5958 39690 6010
rect 39702 5958 39754 6010
rect 1768 5788 1820 5840
rect 33968 5788 34020 5840
rect 56876 5720 56928 5772
rect 57704 5720 57756 5772
rect 58164 5627 58216 5636
rect 58164 5593 58173 5627
rect 58173 5593 58207 5627
rect 58207 5593 58216 5627
rect 58164 5584 58216 5593
rect 40408 5516 40460 5568
rect 53472 5516 53524 5568
rect 57060 5559 57112 5568
rect 57060 5525 57069 5559
rect 57069 5525 57103 5559
rect 57103 5525 57112 5559
rect 57060 5516 57112 5525
rect 10614 5414 10666 5466
rect 10678 5414 10730 5466
rect 10742 5414 10794 5466
rect 10806 5414 10858 5466
rect 29878 5414 29930 5466
rect 29942 5414 29994 5466
rect 30006 5414 30058 5466
rect 30070 5414 30122 5466
rect 49142 5414 49194 5466
rect 49206 5414 49258 5466
rect 49270 5414 49322 5466
rect 49334 5414 49386 5466
rect 16856 5312 16908 5364
rect 33968 5355 34020 5364
rect 1584 5244 1636 5296
rect 18144 5244 18196 5296
rect 33968 5321 33977 5355
rect 33977 5321 34011 5355
rect 34011 5321 34020 5355
rect 33968 5312 34020 5321
rect 36084 5312 36136 5364
rect 34796 5219 34848 5228
rect 34796 5185 34805 5219
rect 34805 5185 34839 5219
rect 34839 5185 34848 5219
rect 34796 5176 34848 5185
rect 21916 5108 21968 5160
rect 25780 5108 25832 5160
rect 41328 5176 41380 5228
rect 41512 5176 41564 5228
rect 56416 5219 56468 5228
rect 56416 5185 56425 5219
rect 56425 5185 56459 5219
rect 56459 5185 56468 5219
rect 56416 5176 56468 5185
rect 57796 5108 57848 5160
rect 56692 5040 56744 5092
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 33968 4972 34020 5024
rect 35624 4972 35676 5024
rect 40500 4972 40552 5024
rect 57612 4972 57664 5024
rect 20246 4870 20298 4922
rect 20310 4870 20362 4922
rect 20374 4870 20426 4922
rect 20438 4870 20490 4922
rect 39510 4870 39562 4922
rect 39574 4870 39626 4922
rect 39638 4870 39690 4922
rect 39702 4870 39754 4922
rect 2412 4811 2464 4820
rect 2412 4777 2421 4811
rect 2421 4777 2455 4811
rect 2455 4777 2464 4811
rect 2412 4768 2464 4777
rect 26240 4768 26292 4820
rect 35624 4768 35676 4820
rect 56876 4768 56928 4820
rect 1400 4700 1452 4752
rect 37648 4743 37700 4752
rect 37648 4709 37657 4743
rect 37657 4709 37691 4743
rect 37691 4709 37700 4743
rect 37648 4700 37700 4709
rect 41236 4700 41288 4752
rect 58072 4743 58124 4752
rect 58072 4709 58081 4743
rect 58081 4709 58115 4743
rect 58115 4709 58124 4743
rect 58072 4700 58124 4709
rect 27436 4675 27488 4684
rect 27436 4641 27445 4675
rect 27445 4641 27479 4675
rect 27479 4641 27488 4675
rect 27436 4632 27488 4641
rect 40500 4632 40552 4684
rect 57612 4632 57664 4684
rect 28724 4564 28776 4616
rect 38476 4564 38528 4616
rect 41144 4564 41196 4616
rect 41420 4564 41472 4616
rect 10232 4496 10284 4548
rect 27712 4496 27764 4548
rect 39120 4496 39172 4548
rect 39856 4496 39908 4548
rect 41052 4496 41104 4548
rect 41328 4496 41380 4548
rect 16028 4428 16080 4480
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 17776 4428 17828 4480
rect 20536 4428 20588 4480
rect 27252 4428 27304 4480
rect 28816 4428 28868 4480
rect 36360 4428 36412 4480
rect 36820 4428 36872 4480
rect 39304 4428 39356 4480
rect 41144 4471 41196 4480
rect 41144 4437 41153 4471
rect 41153 4437 41187 4471
rect 41187 4437 41196 4471
rect 41144 4428 41196 4437
rect 42432 4428 42484 4480
rect 44088 4496 44140 4548
rect 52368 4496 52420 4548
rect 57888 4539 57940 4548
rect 57888 4505 57897 4539
rect 57897 4505 57931 4539
rect 57931 4505 57940 4539
rect 57888 4496 57940 4505
rect 44640 4428 44692 4480
rect 57244 4471 57296 4480
rect 57244 4437 57253 4471
rect 57253 4437 57287 4471
rect 57287 4437 57296 4471
rect 57244 4428 57296 4437
rect 10614 4326 10666 4378
rect 10678 4326 10730 4378
rect 10742 4326 10794 4378
rect 10806 4326 10858 4378
rect 29878 4326 29930 4378
rect 29942 4326 29994 4378
rect 30006 4326 30058 4378
rect 30070 4326 30122 4378
rect 49142 4326 49194 4378
rect 49206 4326 49258 4378
rect 49270 4326 49322 4378
rect 49334 4326 49386 4378
rect 4252 4224 4304 4276
rect 10324 4267 10376 4276
rect 10324 4233 10333 4267
rect 10333 4233 10367 4267
rect 10367 4233 10376 4267
rect 10324 4224 10376 4233
rect 19432 4224 19484 4276
rect 21548 4224 21600 4276
rect 21824 4224 21876 4276
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 25688 4156 25740 4208
rect 25872 4224 25924 4276
rect 28908 4267 28960 4276
rect 28908 4233 28917 4267
rect 28917 4233 28951 4267
rect 28951 4233 28960 4267
rect 28908 4224 28960 4233
rect 29460 4267 29512 4276
rect 29460 4233 29469 4267
rect 29469 4233 29503 4267
rect 29503 4233 29512 4267
rect 29460 4224 29512 4233
rect 37004 4267 37056 4276
rect 37004 4233 37013 4267
rect 37013 4233 37047 4267
rect 37047 4233 37056 4267
rect 37004 4224 37056 4233
rect 43628 4224 43680 4276
rect 43996 4224 44048 4276
rect 57244 4224 57296 4276
rect 58256 4224 58308 4276
rect 26976 4156 27028 4208
rect 28816 4156 28868 4208
rect 57888 4156 57940 4208
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 1952 4020 2004 4072
rect 15200 4063 15252 4072
rect 15200 4029 15209 4063
rect 15209 4029 15243 4063
rect 15243 4029 15252 4063
rect 15200 4020 15252 4029
rect 17592 4020 17644 4072
rect 1308 3952 1360 4004
rect 16672 3952 16724 4004
rect 25780 4088 25832 4140
rect 27252 4088 27304 4140
rect 25044 4063 25096 4072
rect 25044 4029 25053 4063
rect 25053 4029 25087 4063
rect 25087 4029 25096 4063
rect 25044 4020 25096 4029
rect 25688 4063 25740 4072
rect 25688 4029 25697 4063
rect 25697 4029 25731 4063
rect 25731 4029 25740 4063
rect 25688 4020 25740 4029
rect 25872 4063 25924 4072
rect 25872 4029 25881 4063
rect 25881 4029 25915 4063
rect 25915 4029 25924 4063
rect 25872 4020 25924 4029
rect 34612 4020 34664 4072
rect 36820 4063 36872 4072
rect 36820 4029 36829 4063
rect 36829 4029 36863 4063
rect 36863 4029 36872 4063
rect 36820 4020 36872 4029
rect 36084 3952 36136 4004
rect 37464 4020 37516 4072
rect 39396 4020 39448 4072
rect 39856 4020 39908 4072
rect 41052 4020 41104 4072
rect 41420 4020 41472 4072
rect 42432 4063 42484 4072
rect 37372 3952 37424 4004
rect 42432 4029 42441 4063
rect 42441 4029 42475 4063
rect 42475 4029 42484 4063
rect 42432 4020 42484 4029
rect 43812 4020 43864 4072
rect 44088 4063 44140 4072
rect 44088 4029 44097 4063
rect 44097 4029 44131 4063
rect 44131 4029 44140 4063
rect 44088 4020 44140 4029
rect 44272 4088 44324 4140
rect 48412 4088 48464 4140
rect 55128 4131 55180 4140
rect 55128 4097 55137 4131
rect 55137 4097 55171 4131
rect 55171 4097 55180 4131
rect 55128 4088 55180 4097
rect 57980 4088 58032 4140
rect 47124 4020 47176 4072
rect 57796 4020 57848 4072
rect 57888 4020 57940 4072
rect 3148 3927 3200 3936
rect 3148 3893 3157 3927
rect 3157 3893 3191 3927
rect 3191 3893 3200 3927
rect 3148 3884 3200 3893
rect 17408 3884 17460 3936
rect 18696 3927 18748 3936
rect 18696 3893 18705 3927
rect 18705 3893 18739 3927
rect 18739 3893 18748 3927
rect 18696 3884 18748 3893
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 21180 3884 21232 3893
rect 25136 3927 25188 3936
rect 25136 3893 25145 3927
rect 25145 3893 25179 3927
rect 25179 3893 25188 3927
rect 25136 3884 25188 3893
rect 25964 3884 26016 3936
rect 27620 3927 27672 3936
rect 27620 3893 27629 3927
rect 27629 3893 27663 3927
rect 27663 3893 27672 3927
rect 27620 3884 27672 3893
rect 28080 3884 28132 3936
rect 34980 3884 35032 3936
rect 38200 3884 38252 3936
rect 38660 3884 38712 3936
rect 39396 3884 39448 3936
rect 40132 3927 40184 3936
rect 40132 3893 40141 3927
rect 40141 3893 40175 3927
rect 40175 3893 40184 3927
rect 40132 3884 40184 3893
rect 41604 3884 41656 3936
rect 45468 3952 45520 4004
rect 45560 3952 45612 4004
rect 51080 3952 51132 4004
rect 43444 3927 43496 3936
rect 43444 3893 43453 3927
rect 43453 3893 43487 3927
rect 43487 3893 43496 3927
rect 43444 3884 43496 3893
rect 44548 3927 44600 3936
rect 44548 3893 44557 3927
rect 44557 3893 44591 3927
rect 44591 3893 44600 3927
rect 44548 3884 44600 3893
rect 44640 3884 44692 3936
rect 46296 3927 46348 3936
rect 46296 3893 46305 3927
rect 46305 3893 46339 3927
rect 46339 3893 46348 3927
rect 46296 3884 46348 3893
rect 47308 3884 47360 3936
rect 47584 3927 47636 3936
rect 47584 3893 47593 3927
rect 47593 3893 47627 3927
rect 47627 3893 47636 3927
rect 47584 3884 47636 3893
rect 55588 3884 55640 3936
rect 57520 3927 57572 3936
rect 57520 3893 57529 3927
rect 57529 3893 57563 3927
rect 57563 3893 57572 3927
rect 57520 3884 57572 3893
rect 20246 3782 20298 3834
rect 20310 3782 20362 3834
rect 20374 3782 20426 3834
rect 20438 3782 20490 3834
rect 39510 3782 39562 3834
rect 39574 3782 39626 3834
rect 39638 3782 39690 3834
rect 39702 3782 39754 3834
rect 11520 3723 11572 3732
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 14372 3723 14424 3732
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 15476 3680 15528 3732
rect 22560 3723 22612 3732
rect 22560 3689 22569 3723
rect 22569 3689 22603 3723
rect 22603 3689 22612 3723
rect 22560 3680 22612 3689
rect 25780 3723 25832 3732
rect 25780 3689 25789 3723
rect 25789 3689 25823 3723
rect 25823 3689 25832 3723
rect 25780 3680 25832 3689
rect 30472 3723 30524 3732
rect 30472 3689 30481 3723
rect 30481 3689 30515 3723
rect 30515 3689 30524 3723
rect 30472 3680 30524 3689
rect 31208 3680 31260 3732
rect 32404 3723 32456 3732
rect 32404 3689 32413 3723
rect 32413 3689 32447 3723
rect 32447 3689 32456 3723
rect 32404 3680 32456 3689
rect 34796 3680 34848 3732
rect 38752 3680 38804 3732
rect 41420 3680 41472 3732
rect 42432 3680 42484 3732
rect 43628 3680 43680 3732
rect 2044 3612 2096 3664
rect 4252 3612 4304 3664
rect 11060 3612 11112 3664
rect 9220 3544 9272 3596
rect 15384 3544 15436 3596
rect 16488 3612 16540 3664
rect 57980 3655 58032 3664
rect 57980 3621 57989 3655
rect 57989 3621 58023 3655
rect 58023 3621 58032 3655
rect 57980 3612 58032 3621
rect 16764 3587 16816 3596
rect 16764 3553 16773 3587
rect 16773 3553 16807 3587
rect 16807 3553 16816 3587
rect 16764 3544 16816 3553
rect 17408 3587 17460 3596
rect 17408 3553 17417 3587
rect 17417 3553 17451 3587
rect 17451 3553 17460 3587
rect 17408 3544 17460 3553
rect 18420 3587 18472 3596
rect 18420 3553 18429 3587
rect 18429 3553 18463 3587
rect 18463 3553 18472 3587
rect 18420 3544 18472 3553
rect 18696 3544 18748 3596
rect 21180 3544 21232 3596
rect 22652 3544 22704 3596
rect 26148 3544 26200 3596
rect 27804 3544 27856 3596
rect 28080 3544 28132 3596
rect 28724 3587 28776 3596
rect 28724 3553 28733 3587
rect 28733 3553 28767 3587
rect 28767 3553 28776 3587
rect 28724 3544 28776 3553
rect 480 3408 532 3460
rect 21916 3476 21968 3528
rect 22192 3476 22244 3528
rect 27620 3476 27672 3528
rect 30196 3544 30248 3596
rect 32220 3587 32272 3596
rect 32220 3553 32229 3587
rect 32229 3553 32263 3587
rect 32263 3553 32272 3587
rect 32220 3544 32272 3553
rect 34060 3587 34112 3596
rect 34060 3553 34069 3587
rect 34069 3553 34103 3587
rect 34103 3553 34112 3587
rect 34060 3544 34112 3553
rect 34980 3544 35032 3596
rect 36636 3544 36688 3596
rect 37372 3544 37424 3596
rect 38200 3544 38252 3596
rect 38660 3587 38712 3596
rect 38660 3553 38669 3587
rect 38669 3553 38703 3587
rect 38703 3553 38712 3587
rect 38660 3544 38712 3553
rect 40132 3544 40184 3596
rect 41144 3587 41196 3596
rect 41144 3553 41153 3587
rect 41153 3553 41187 3587
rect 41187 3553 41196 3587
rect 41144 3544 41196 3553
rect 41604 3544 41656 3596
rect 43444 3544 43496 3596
rect 43996 3587 44048 3596
rect 43996 3553 44005 3587
rect 44005 3553 44039 3587
rect 44039 3553 44048 3587
rect 43996 3544 44048 3553
rect 18144 3408 18196 3460
rect 19432 3408 19484 3460
rect 26332 3408 26384 3460
rect 27160 3451 27212 3460
rect 27160 3417 27169 3451
rect 27169 3417 27203 3451
rect 27203 3417 27212 3451
rect 27160 3408 27212 3417
rect 43720 3476 43772 3528
rect 36360 3451 36412 3460
rect 36360 3417 36369 3451
rect 36369 3417 36403 3451
rect 36403 3417 36412 3451
rect 36360 3408 36412 3417
rect 39396 3408 39448 3460
rect 41880 3451 41932 3460
rect 41880 3417 41889 3451
rect 41889 3417 41923 3451
rect 41923 3417 41932 3451
rect 41880 3408 41932 3417
rect 43996 3408 44048 3460
rect 47860 3476 47912 3528
rect 57060 3544 57112 3596
rect 57244 3587 57296 3596
rect 57244 3553 57253 3587
rect 57253 3553 57287 3587
rect 57287 3553 57296 3587
rect 57244 3544 57296 3553
rect 58072 3476 58124 3528
rect 54208 3408 54260 3460
rect 57428 3451 57480 3460
rect 57428 3417 57437 3451
rect 57437 3417 57471 3451
rect 57471 3417 57480 3451
rect 57428 3408 57480 3417
rect 58900 3408 58952 3460
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 2596 3340 2648 3392
rect 3240 3340 3292 3392
rect 6460 3340 6512 3392
rect 10508 3340 10560 3392
rect 13268 3383 13320 3392
rect 13268 3349 13277 3383
rect 13277 3349 13311 3383
rect 13311 3349 13320 3383
rect 13268 3340 13320 3349
rect 14372 3340 14424 3392
rect 17500 3383 17552 3392
rect 17500 3349 17509 3383
rect 17509 3349 17543 3383
rect 17543 3349 17552 3383
rect 17500 3340 17552 3349
rect 18604 3383 18656 3392
rect 18604 3349 18613 3383
rect 18613 3349 18647 3383
rect 18647 3349 18656 3383
rect 18604 3340 18656 3349
rect 19616 3383 19668 3392
rect 19616 3349 19625 3383
rect 19625 3349 19659 3383
rect 19659 3349 19668 3383
rect 19616 3340 19668 3349
rect 20536 3340 20588 3392
rect 20720 3340 20772 3392
rect 22008 3383 22060 3392
rect 22008 3349 22017 3383
rect 22017 3349 22051 3383
rect 22051 3349 22060 3383
rect 22008 3340 22060 3349
rect 24308 3383 24360 3392
rect 24308 3349 24317 3383
rect 24317 3349 24351 3383
rect 24351 3349 24360 3383
rect 24308 3340 24360 3349
rect 28632 3383 28684 3392
rect 28632 3349 28641 3383
rect 28641 3349 28675 3383
rect 28675 3349 28684 3383
rect 28632 3340 28684 3349
rect 29736 3340 29788 3392
rect 34612 3340 34664 3392
rect 36452 3340 36504 3392
rect 38292 3340 38344 3392
rect 40592 3340 40644 3392
rect 41788 3340 41840 3392
rect 42800 3340 42852 3392
rect 43168 3383 43220 3392
rect 43168 3349 43177 3383
rect 43177 3349 43211 3383
rect 43211 3349 43220 3383
rect 43168 3340 43220 3349
rect 44088 3340 44140 3392
rect 45836 3383 45888 3392
rect 45836 3349 45845 3383
rect 45845 3349 45879 3383
rect 45879 3349 45888 3383
rect 45836 3340 45888 3349
rect 46020 3340 46072 3392
rect 47032 3340 47084 3392
rect 49608 3383 49660 3392
rect 49608 3349 49617 3383
rect 49617 3349 49651 3383
rect 49651 3349 49660 3383
rect 49608 3340 49660 3349
rect 50068 3383 50120 3392
rect 50068 3349 50077 3383
rect 50077 3349 50111 3383
rect 50111 3349 50120 3383
rect 50068 3340 50120 3349
rect 52368 3340 52420 3392
rect 52552 3383 52604 3392
rect 52552 3349 52561 3383
rect 52561 3349 52595 3383
rect 52595 3349 52604 3383
rect 52552 3340 52604 3349
rect 53196 3383 53248 3392
rect 53196 3349 53205 3383
rect 53205 3349 53239 3383
rect 53239 3349 53248 3383
rect 53196 3340 53248 3349
rect 53380 3340 53432 3392
rect 55680 3340 55732 3392
rect 56324 3383 56376 3392
rect 56324 3349 56333 3383
rect 56333 3349 56367 3383
rect 56367 3349 56376 3383
rect 56324 3340 56376 3349
rect 10614 3238 10666 3290
rect 10678 3238 10730 3290
rect 10742 3238 10794 3290
rect 10806 3238 10858 3290
rect 29878 3238 29930 3290
rect 29942 3238 29994 3290
rect 30006 3238 30058 3290
rect 30070 3238 30122 3290
rect 49142 3238 49194 3290
rect 49206 3238 49258 3290
rect 49270 3238 49322 3290
rect 49334 3238 49386 3290
rect 7012 3179 7064 3188
rect 7012 3145 7021 3179
rect 7021 3145 7055 3179
rect 7055 3145 7064 3179
rect 7012 3136 7064 3145
rect 8668 3136 8720 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 14188 3136 14240 3188
rect 16764 3136 16816 3188
rect 17040 3179 17092 3188
rect 17040 3145 17049 3179
rect 17049 3145 17083 3179
rect 17083 3145 17092 3179
rect 17040 3136 17092 3145
rect 19800 3179 19852 3188
rect 19800 3145 19809 3179
rect 19809 3145 19843 3179
rect 19843 3145 19852 3179
rect 19800 3136 19852 3145
rect 27804 3179 27856 3188
rect 27804 3145 27813 3179
rect 27813 3145 27847 3179
rect 27847 3145 27856 3179
rect 27804 3136 27856 3145
rect 29368 3136 29420 3188
rect 1400 2975 1452 2984
rect 1400 2941 1409 2975
rect 1409 2941 1443 2975
rect 1443 2941 1452 2975
rect 1400 2932 1452 2941
rect 2412 2932 2464 2984
rect 3148 2932 3200 2984
rect 35072 3068 35124 3120
rect 36544 3068 36596 3120
rect 37832 3068 37884 3120
rect 38384 3111 38436 3120
rect 38384 3077 38393 3111
rect 38393 3077 38427 3111
rect 38427 3077 38436 3111
rect 38384 3068 38436 3077
rect 16212 3000 16264 3052
rect 6460 2932 6512 2984
rect 8760 2932 8812 2984
rect 9680 2932 9732 2984
rect 11520 2932 11572 2984
rect 13084 2975 13136 2984
rect 13084 2941 13093 2975
rect 13093 2941 13127 2975
rect 13127 2941 13136 2975
rect 13084 2932 13136 2941
rect 13268 2932 13320 2984
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 15476 2932 15528 2984
rect 16856 2932 16908 2984
rect 17500 2932 17552 2984
rect 19432 3000 19484 3052
rect 27620 3000 27672 3052
rect 29644 3000 29696 3052
rect 35348 3000 35400 3052
rect 36176 3043 36228 3052
rect 36176 3009 36185 3043
rect 36185 3009 36219 3043
rect 36219 3009 36228 3043
rect 36176 3000 36228 3009
rect 41604 3068 41656 3120
rect 42340 3111 42392 3120
rect 40040 3000 40092 3052
rect 41052 3043 41104 3052
rect 41052 3009 41061 3043
rect 41061 3009 41095 3043
rect 41095 3009 41104 3043
rect 41052 3000 41104 3009
rect 41236 3043 41288 3052
rect 41236 3009 41245 3043
rect 41245 3009 41279 3043
rect 41279 3009 41288 3043
rect 41236 3000 41288 3009
rect 19340 2932 19392 2984
rect 19616 2975 19668 2984
rect 19616 2941 19625 2975
rect 19625 2941 19659 2975
rect 19659 2941 19668 2975
rect 19616 2932 19668 2941
rect 20720 2975 20772 2984
rect 20720 2941 20729 2975
rect 20729 2941 20763 2975
rect 20763 2941 20772 2975
rect 20720 2932 20772 2941
rect 22100 2932 22152 2984
rect 2320 2907 2372 2916
rect 2320 2873 2329 2907
rect 2329 2873 2363 2907
rect 2363 2873 2372 2907
rect 2320 2864 2372 2873
rect 2780 2907 2832 2916
rect 2780 2873 2789 2907
rect 2789 2873 2823 2907
rect 2823 2873 2832 2907
rect 2780 2864 2832 2873
rect 4160 2907 4212 2916
rect 4160 2873 4169 2907
rect 4169 2873 4203 2907
rect 4203 2873 4212 2907
rect 4160 2864 4212 2873
rect 4620 2864 4672 2916
rect 5724 2907 5776 2916
rect 5724 2873 5733 2907
rect 5733 2873 5767 2907
rect 5767 2873 5776 2907
rect 5724 2864 5776 2873
rect 12164 2864 12216 2916
rect 12900 2907 12952 2916
rect 12900 2873 12909 2907
rect 12909 2873 12943 2907
rect 12943 2873 12952 2907
rect 12900 2864 12952 2873
rect 14280 2907 14332 2916
rect 14280 2873 14289 2907
rect 14289 2873 14323 2907
rect 14323 2873 14332 2907
rect 14280 2864 14332 2873
rect 14464 2907 14516 2916
rect 14464 2873 14473 2907
rect 14473 2873 14507 2907
rect 14507 2873 14516 2907
rect 14464 2864 14516 2873
rect 16120 2907 16172 2916
rect 16120 2873 16129 2907
rect 16129 2873 16163 2907
rect 16163 2873 16172 2907
rect 16120 2864 16172 2873
rect 24308 2932 24360 2984
rect 25136 2975 25188 2984
rect 25136 2941 25145 2975
rect 25145 2941 25179 2975
rect 25179 2941 25188 2975
rect 25136 2932 25188 2941
rect 25964 2975 26016 2984
rect 25964 2941 25973 2975
rect 25973 2941 26007 2975
rect 26007 2941 26016 2975
rect 25964 2932 26016 2941
rect 26240 2932 26292 2984
rect 26976 2932 27028 2984
rect 28816 2932 28868 2984
rect 28908 2932 28960 2984
rect 29736 2932 29788 2984
rect 31208 2932 31260 2984
rect 31944 2975 31996 2984
rect 31944 2941 31953 2975
rect 31953 2941 31987 2975
rect 31987 2941 31996 2975
rect 31944 2932 31996 2941
rect 33600 2975 33652 2984
rect 33600 2941 33609 2975
rect 33609 2941 33643 2975
rect 33643 2941 33652 2975
rect 33600 2932 33652 2941
rect 34612 2975 34664 2984
rect 34612 2941 34621 2975
rect 34621 2941 34655 2975
rect 34655 2941 34664 2975
rect 34612 2932 34664 2941
rect 36452 2975 36504 2984
rect 36452 2941 36461 2975
rect 36461 2941 36495 2975
rect 36495 2941 36504 2975
rect 36452 2932 36504 2941
rect 37648 2932 37700 2984
rect 38292 2975 38344 2984
rect 38292 2941 38301 2975
rect 38301 2941 38335 2975
rect 38335 2941 38344 2975
rect 38292 2932 38344 2941
rect 39488 2932 39540 2984
rect 7380 2796 7432 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 11980 2796 12032 2848
rect 19064 2839 19116 2848
rect 19064 2805 19073 2839
rect 19073 2805 19107 2839
rect 19107 2805 19116 2839
rect 19064 2796 19116 2805
rect 24860 2864 24912 2916
rect 25320 2907 25372 2916
rect 25320 2873 25329 2907
rect 25329 2873 25363 2907
rect 25363 2873 25372 2907
rect 25320 2864 25372 2873
rect 25780 2907 25832 2916
rect 25780 2873 25789 2907
rect 25789 2873 25823 2907
rect 25823 2873 25832 2907
rect 25780 2864 25832 2873
rect 30380 2864 30432 2916
rect 31760 2907 31812 2916
rect 31760 2873 31769 2907
rect 31769 2873 31803 2907
rect 31803 2873 31812 2907
rect 31760 2864 31812 2873
rect 34704 2864 34756 2916
rect 36268 2864 36320 2916
rect 40132 2864 40184 2916
rect 22100 2796 22152 2848
rect 22560 2839 22612 2848
rect 22560 2805 22569 2839
rect 22569 2805 22603 2839
rect 22603 2805 22612 2839
rect 22560 2796 22612 2805
rect 25872 2796 25924 2848
rect 26792 2839 26844 2848
rect 26792 2805 26801 2839
rect 26801 2805 26835 2839
rect 26835 2805 26844 2839
rect 26792 2796 26844 2805
rect 33784 2839 33836 2848
rect 33784 2805 33793 2839
rect 33793 2805 33827 2839
rect 33827 2805 33836 2839
rect 33784 2796 33836 2805
rect 39948 2796 40000 2848
rect 40592 2932 40644 2984
rect 41512 3000 41564 3052
rect 42340 3077 42349 3111
rect 42349 3077 42383 3111
rect 42383 3077 42392 3111
rect 42340 3068 42392 3077
rect 43628 3111 43680 3120
rect 43628 3077 43637 3111
rect 43637 3077 43671 3111
rect 43671 3077 43680 3111
rect 43628 3068 43680 3077
rect 45468 3111 45520 3120
rect 45468 3077 45477 3111
rect 45477 3077 45511 3111
rect 45511 3077 45520 3111
rect 45468 3068 45520 3077
rect 47124 3136 47176 3188
rect 53104 3179 53156 3188
rect 49700 3111 49752 3120
rect 49700 3077 49709 3111
rect 49709 3077 49743 3111
rect 49743 3077 49752 3111
rect 49700 3068 49752 3077
rect 50804 3068 50856 3120
rect 53104 3145 53113 3179
rect 53113 3145 53147 3179
rect 53147 3145 53156 3179
rect 53104 3136 53156 3145
rect 44088 3043 44140 3052
rect 44088 3009 44097 3043
rect 44097 3009 44131 3043
rect 44131 3009 44140 3043
rect 44088 3000 44140 3009
rect 55588 3068 55640 3120
rect 56416 3136 56468 3188
rect 57152 3136 57204 3188
rect 45100 2932 45152 2984
rect 45836 2932 45888 2984
rect 46940 2932 46992 2984
rect 47032 2932 47084 2984
rect 47584 2932 47636 2984
rect 41236 2864 41288 2916
rect 42064 2864 42116 2916
rect 42800 2864 42852 2916
rect 44180 2907 44232 2916
rect 44180 2873 44189 2907
rect 44189 2873 44223 2907
rect 44223 2873 44232 2907
rect 44180 2864 44232 2873
rect 44640 2864 44692 2916
rect 44916 2907 44968 2916
rect 44916 2873 44925 2907
rect 44925 2873 44959 2907
rect 44959 2873 44968 2907
rect 44916 2864 44968 2873
rect 46480 2907 46532 2916
rect 46480 2873 46489 2907
rect 46489 2873 46523 2907
rect 46523 2873 46532 2907
rect 46480 2864 46532 2873
rect 43996 2796 44048 2848
rect 44272 2796 44324 2848
rect 44364 2796 44416 2848
rect 48320 2864 48372 2916
rect 49700 2932 49752 2984
rect 50068 2932 50120 2984
rect 52552 2932 52604 2984
rect 52920 2975 52972 2984
rect 52920 2941 52929 2975
rect 52929 2941 52963 2975
rect 52963 2941 52972 2975
rect 52920 2932 52972 2941
rect 53196 2932 53248 2984
rect 54024 2975 54076 2984
rect 54024 2941 54033 2975
rect 54033 2941 54067 2975
rect 54067 2941 54076 2975
rect 54024 2932 54076 2941
rect 54208 2975 54260 2984
rect 54208 2941 54217 2975
rect 54217 2941 54251 2975
rect 54251 2941 54260 2975
rect 54208 2932 54260 2941
rect 54944 2975 54996 2984
rect 54944 2941 54953 2975
rect 54953 2941 54987 2975
rect 54987 2941 54996 2975
rect 54944 2932 54996 2941
rect 56324 2932 56376 2984
rect 57520 2975 57572 2984
rect 57520 2941 57529 2975
rect 57529 2941 57563 2975
rect 57563 2941 57572 2975
rect 57520 2932 57572 2941
rect 50160 2864 50212 2916
rect 50620 2907 50672 2916
rect 50620 2873 50629 2907
rect 50629 2873 50663 2907
rect 50663 2873 50672 2907
rect 50620 2864 50672 2873
rect 51540 2907 51592 2916
rect 51540 2873 51549 2907
rect 51549 2873 51583 2907
rect 51583 2873 51592 2907
rect 51540 2864 51592 2873
rect 54760 2907 54812 2916
rect 54760 2873 54769 2907
rect 54769 2873 54803 2907
rect 54803 2873 54812 2907
rect 54760 2864 54812 2873
rect 56508 2907 56560 2916
rect 56508 2873 56517 2907
rect 56517 2873 56551 2907
rect 56551 2873 56560 2907
rect 56508 2864 56560 2873
rect 52276 2839 52328 2848
rect 52276 2805 52285 2839
rect 52285 2805 52319 2839
rect 52319 2805 52328 2839
rect 52276 2796 52328 2805
rect 54116 2839 54168 2848
rect 54116 2805 54125 2839
rect 54125 2805 54159 2839
rect 54159 2805 54168 2839
rect 54116 2796 54168 2805
rect 56600 2839 56652 2848
rect 56600 2805 56609 2839
rect 56609 2805 56643 2839
rect 56643 2805 56652 2839
rect 56600 2796 56652 2805
rect 20246 2694 20298 2746
rect 20310 2694 20362 2746
rect 20374 2694 20426 2746
rect 20438 2694 20490 2746
rect 39510 2694 39562 2746
rect 39574 2694 39626 2746
rect 39638 2694 39690 2746
rect 39702 2694 39754 2746
rect 8760 2592 8812 2644
rect 1676 2567 1728 2576
rect 1676 2533 1685 2567
rect 1685 2533 1719 2567
rect 1719 2533 1728 2567
rect 1676 2524 1728 2533
rect 8300 2567 8352 2576
rect 8300 2533 8309 2567
rect 8309 2533 8343 2567
rect 8343 2533 8352 2567
rect 8300 2524 8352 2533
rect 10324 2524 10376 2576
rect 940 2456 992 2508
rect 3240 2456 3292 2508
rect 5540 2456 5592 2508
rect 7380 2456 7432 2508
rect 12440 2592 12492 2644
rect 14372 2592 14424 2644
rect 14464 2592 14516 2644
rect 15292 2635 15344 2644
rect 15292 2601 15301 2635
rect 15301 2601 15335 2635
rect 15335 2601 15344 2635
rect 15292 2592 15344 2601
rect 13820 2567 13872 2576
rect 10508 2456 10560 2508
rect 13820 2533 13829 2567
rect 13829 2533 13863 2567
rect 13863 2533 13872 2567
rect 13820 2524 13872 2533
rect 16028 2524 16080 2576
rect 16212 2524 16264 2576
rect 11980 2456 12032 2508
rect 14188 2456 14240 2508
rect 17500 2524 17552 2576
rect 18144 2567 18196 2576
rect 18144 2533 18153 2567
rect 18153 2533 18187 2567
rect 18187 2533 18196 2567
rect 18144 2524 18196 2533
rect 19892 2524 19944 2576
rect 20628 2524 20680 2576
rect 22008 2592 22060 2644
rect 23480 2592 23532 2644
rect 29368 2635 29420 2644
rect 21916 2524 21968 2576
rect 29368 2601 29377 2635
rect 29377 2601 29411 2635
rect 29411 2601 29420 2635
rect 29368 2592 29420 2601
rect 33140 2592 33192 2644
rect 35072 2635 35124 2644
rect 35072 2601 35081 2635
rect 35081 2601 35115 2635
rect 35115 2601 35124 2635
rect 35072 2592 35124 2601
rect 37372 2635 37424 2644
rect 37372 2601 37381 2635
rect 37381 2601 37415 2635
rect 37415 2601 37424 2635
rect 37372 2592 37424 2601
rect 40132 2592 40184 2644
rect 41604 2592 41656 2644
rect 43076 2592 43128 2644
rect 43168 2635 43220 2644
rect 43168 2601 43177 2635
rect 43177 2601 43211 2635
rect 43211 2601 43220 2635
rect 43168 2592 43220 2601
rect 43352 2592 43404 2644
rect 44364 2592 44416 2644
rect 44916 2592 44968 2644
rect 46940 2635 46992 2644
rect 46940 2601 46949 2635
rect 46949 2601 46983 2635
rect 46983 2601 46992 2635
rect 46940 2592 46992 2601
rect 49608 2592 49660 2644
rect 50804 2592 50856 2644
rect 51080 2592 51132 2644
rect 27436 2524 27488 2576
rect 28540 2524 28592 2576
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 13728 2388 13780 2440
rect 20536 2456 20588 2508
rect 22560 2456 22612 2508
rect 6000 2320 6052 2372
rect 7840 2320 7892 2372
rect 15660 2320 15712 2372
rect 17776 2320 17828 2372
rect 22192 2388 22244 2440
rect 18880 2363 18932 2372
rect 18880 2329 18889 2363
rect 18889 2329 18923 2363
rect 18923 2329 18932 2363
rect 18880 2320 18932 2329
rect 20260 2363 20312 2372
rect 20260 2329 20269 2363
rect 20269 2329 20303 2363
rect 20303 2329 20312 2363
rect 20260 2320 20312 2329
rect 21640 2320 21692 2372
rect 23940 2363 23992 2372
rect 23940 2329 23949 2363
rect 23949 2329 23983 2363
rect 23983 2329 23992 2363
rect 23940 2320 23992 2329
rect 25872 2456 25924 2508
rect 26332 2499 26384 2508
rect 26332 2465 26341 2499
rect 26341 2465 26375 2499
rect 26375 2465 26384 2499
rect 26332 2456 26384 2465
rect 29000 2456 29052 2508
rect 31484 2567 31536 2576
rect 31484 2533 31493 2567
rect 31493 2533 31527 2567
rect 31527 2533 31536 2567
rect 31484 2524 31536 2533
rect 29460 2456 29512 2508
rect 29736 2456 29788 2508
rect 26056 2431 26108 2440
rect 26056 2397 26065 2431
rect 26065 2397 26099 2431
rect 26099 2397 26108 2431
rect 26056 2388 26108 2397
rect 26148 2388 26200 2440
rect 28264 2320 28316 2372
rect 31300 2363 31352 2372
rect 31300 2329 31309 2363
rect 31309 2329 31343 2363
rect 31343 2329 31352 2363
rect 31300 2320 31352 2329
rect 3792 2252 3844 2304
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 12348 2252 12400 2304
rect 13728 2252 13780 2304
rect 13820 2252 13872 2304
rect 17684 2295 17736 2304
rect 17684 2261 17693 2295
rect 17693 2261 17727 2295
rect 17727 2261 17736 2295
rect 17684 2252 17736 2261
rect 21364 2295 21416 2304
rect 21364 2261 21373 2295
rect 21373 2261 21407 2295
rect 21407 2261 21416 2295
rect 21364 2252 21416 2261
rect 33232 2456 33284 2508
rect 36084 2456 36136 2508
rect 36268 2499 36320 2508
rect 36268 2465 36277 2499
rect 36277 2465 36311 2499
rect 36311 2465 36320 2499
rect 36268 2456 36320 2465
rect 36544 2499 36596 2508
rect 36544 2465 36553 2499
rect 36553 2465 36587 2499
rect 36587 2465 36596 2499
rect 36544 2456 36596 2465
rect 37832 2499 37884 2508
rect 37832 2465 37841 2499
rect 37841 2465 37875 2499
rect 37875 2465 37884 2499
rect 39120 2499 39172 2508
rect 37832 2456 37884 2465
rect 39120 2465 39129 2499
rect 39129 2465 39163 2499
rect 39163 2465 39172 2499
rect 39120 2456 39172 2465
rect 39304 2456 39356 2508
rect 39764 2456 39816 2508
rect 40408 2499 40460 2508
rect 40408 2465 40417 2499
rect 40417 2465 40451 2499
rect 40451 2465 40460 2499
rect 41604 2499 41656 2508
rect 40408 2456 40460 2465
rect 41604 2465 41613 2499
rect 41613 2465 41647 2499
rect 41647 2465 41656 2499
rect 41604 2456 41656 2465
rect 41788 2499 41840 2508
rect 41788 2465 41797 2499
rect 41797 2465 41831 2499
rect 41831 2465 41840 2499
rect 41788 2456 41840 2465
rect 39856 2388 39908 2440
rect 41236 2388 41288 2440
rect 35440 2320 35492 2372
rect 36452 2320 36504 2372
rect 42064 2388 42116 2440
rect 44548 2456 44600 2508
rect 44916 2499 44968 2508
rect 44916 2465 44925 2499
rect 44925 2465 44959 2499
rect 44959 2465 44968 2499
rect 44916 2456 44968 2465
rect 45560 2456 45612 2508
rect 45744 2499 45796 2508
rect 45744 2465 45753 2499
rect 45753 2465 45787 2499
rect 45787 2465 45796 2499
rect 45744 2456 45796 2465
rect 46020 2456 46072 2508
rect 47308 2499 47360 2508
rect 47308 2465 47317 2499
rect 47317 2465 47351 2499
rect 47351 2465 47360 2499
rect 47308 2456 47360 2465
rect 43812 2388 43864 2440
rect 44180 2388 44232 2440
rect 47400 2431 47452 2440
rect 47400 2397 47409 2431
rect 47409 2397 47443 2431
rect 47443 2397 47452 2431
rect 47400 2388 47452 2397
rect 48412 2456 48464 2508
rect 49516 2456 49568 2508
rect 52276 2524 52328 2576
rect 54116 2524 54168 2576
rect 55588 2524 55640 2576
rect 50528 2499 50580 2508
rect 50528 2465 50537 2499
rect 50537 2465 50571 2499
rect 50571 2465 50580 2499
rect 50528 2456 50580 2465
rect 52368 2456 52420 2508
rect 53380 2456 53432 2508
rect 55680 2456 55732 2508
rect 57704 2499 57756 2508
rect 57704 2465 57713 2499
rect 57713 2465 57747 2499
rect 57747 2465 57756 2499
rect 57704 2456 57756 2465
rect 58072 2499 58124 2508
rect 58072 2465 58081 2499
rect 58081 2465 58115 2499
rect 58115 2465 58124 2499
rect 58072 2456 58124 2465
rect 59360 2456 59412 2508
rect 35348 2252 35400 2304
rect 37280 2252 37332 2304
rect 42524 2252 42576 2304
rect 42708 2295 42760 2304
rect 42708 2261 42717 2295
rect 42717 2261 42751 2295
rect 42751 2261 42760 2295
rect 42708 2252 42760 2261
rect 46296 2252 46348 2304
rect 50804 2388 50856 2440
rect 48504 2295 48556 2304
rect 48504 2261 48513 2295
rect 48513 2261 48547 2295
rect 48547 2261 48556 2295
rect 48504 2252 48556 2261
rect 49516 2252 49568 2304
rect 50620 2252 50672 2304
rect 53472 2295 53524 2304
rect 53472 2261 53481 2295
rect 53481 2261 53515 2295
rect 53515 2261 53524 2295
rect 53472 2252 53524 2261
rect 54300 2320 54352 2372
rect 56140 2320 56192 2372
rect 55864 2252 55916 2304
rect 57244 2252 57296 2304
rect 10614 2150 10666 2202
rect 10678 2150 10730 2202
rect 10742 2150 10794 2202
rect 10806 2150 10858 2202
rect 29878 2150 29930 2202
rect 29942 2150 29994 2202
rect 30006 2150 30058 2202
rect 30070 2150 30122 2202
rect 49142 2150 49194 2202
rect 49206 2150 49258 2202
rect 49270 2150 49322 2202
rect 49334 2150 49386 2202
rect 13084 2048 13136 2100
rect 37372 2048 37424 2100
rect 40316 2048 40368 2100
rect 48504 2048 48556 2100
rect 24308 1980 24360 2032
rect 42708 1980 42760 2032
rect 47400 1980 47452 2032
rect 56692 1980 56744 2032
rect 1860 1912 1912 1964
rect 17684 1912 17736 1964
rect 18604 1912 18656 1964
rect 41512 1912 41564 1964
rect 42524 1912 42576 1964
rect 48412 1912 48464 1964
rect 55864 1912 55916 1964
rect 14924 1844 14976 1896
rect 21364 1844 21416 1896
rect 22008 1844 22060 1896
rect 53472 1844 53524 1896
rect 12348 1776 12400 1828
rect 20076 1776 20128 1828
rect 26056 1776 26108 1828
rect 52368 1776 52420 1828
rect 5724 1708 5776 1760
rect 47308 1708 47360 1760
rect 56508 1708 56560 1760
rect 3792 1640 3844 1692
rect 28356 1640 28408 1692
rect 33784 1640 33836 1692
rect 50528 1640 50580 1692
rect 7564 1572 7616 1624
rect 39764 1572 39816 1624
rect 13728 1504 13780 1556
rect 44916 1504 44968 1556
<< metal2 >>
rect 938 29200 994 30000
rect 1398 29200 1454 30000
rect 2318 29200 2374 30000
rect 2778 29200 2834 30000
rect 3238 29200 3294 30000
rect 4158 29200 4214 30000
rect 4618 29200 4674 30000
rect 5538 29200 5594 30000
rect 5998 29200 6054 30000
rect 6458 29200 6514 30000
rect 7378 29200 7434 30000
rect 7838 29200 7894 30000
rect 8758 29200 8814 30000
rect 9218 29200 9274 30000
rect 9678 29200 9734 30000
rect 10598 29200 10654 30000
rect 11058 29200 11114 30000
rect 11978 29200 12034 30000
rect 12438 29200 12494 30000
rect 12898 29200 12954 30000
rect 13818 29200 13874 30000
rect 14278 29200 14334 30000
rect 14738 29200 14794 30000
rect 15658 29200 15714 30000
rect 16118 29200 16174 30000
rect 17038 29200 17094 30000
rect 17498 29200 17554 30000
rect 17958 29200 18014 30000
rect 18878 29200 18934 30000
rect 19338 29200 19394 30000
rect 20258 29200 20314 30000
rect 20718 29200 20774 30000
rect 21178 29200 21234 30000
rect 22098 29200 22154 30000
rect 22558 29200 22614 30000
rect 23478 29200 23534 30000
rect 23938 29200 23994 30000
rect 24398 29200 24454 30000
rect 25318 29200 25374 30000
rect 25778 29200 25834 30000
rect 26698 29200 26754 30000
rect 27158 29200 27214 30000
rect 27618 29200 27674 30000
rect 28538 29200 28594 30000
rect 28998 29200 29054 30000
rect 29918 29200 29974 30000
rect 30378 29200 30434 30000
rect 30838 29200 30894 30000
rect 31758 29200 31814 30000
rect 32218 29200 32274 30000
rect 33138 29200 33194 30000
rect 33598 29200 33654 30000
rect 34058 29200 34114 30000
rect 34978 29200 35034 30000
rect 35438 29200 35494 30000
rect 36358 29200 36414 30000
rect 36818 29200 36874 30000
rect 37278 29200 37334 30000
rect 38198 29200 38254 30000
rect 38658 29200 38714 30000
rect 39578 29200 39634 30000
rect 40038 29200 40094 30000
rect 40498 29200 40554 30000
rect 41418 29200 41474 30000
rect 41878 29200 41934 30000
rect 42798 29200 42854 30000
rect 43258 29200 43314 30000
rect 43718 29200 43774 30000
rect 44638 29200 44694 30000
rect 45098 29200 45154 30000
rect 45558 29200 45614 30000
rect 46478 29200 46534 30000
rect 46938 29200 46994 30000
rect 47858 29200 47914 30000
rect 48318 29200 48374 30000
rect 48778 29200 48834 30000
rect 49698 29200 49754 30000
rect 50158 29200 50214 30000
rect 51078 29200 51134 30000
rect 51538 29200 51594 30000
rect 51998 29200 52054 30000
rect 52918 29200 52974 30000
rect 53378 29200 53434 30000
rect 54298 29200 54354 30000
rect 54758 29200 54814 30000
rect 55218 29200 55274 30000
rect 56138 29200 56194 30000
rect 56598 29200 56654 30000
rect 57518 29200 57574 30000
rect 57978 29200 58034 30000
rect 58438 29200 58494 30000
rect 59358 29200 59414 30000
rect 952 27538 980 29200
rect 940 27532 992 27538
rect 940 27474 992 27480
rect 1412 27062 1440 29200
rect 2228 27532 2280 27538
rect 2228 27474 2280 27480
rect 1582 27432 1638 27441
rect 1582 27367 1638 27376
rect 1490 27296 1546 27305
rect 1490 27231 1546 27240
rect 1400 27056 1452 27062
rect 1400 26998 1452 27004
rect 1504 26926 1532 27231
rect 1492 26920 1544 26926
rect 1492 26862 1544 26868
rect 1398 25936 1454 25945
rect 1398 25871 1400 25880
rect 1452 25871 1454 25880
rect 1400 25842 1452 25848
rect 1398 25256 1454 25265
rect 1398 25191 1400 25200
rect 1452 25191 1454 25200
rect 1400 25162 1452 25168
rect 1504 24954 1532 26862
rect 1596 26518 1624 27367
rect 1768 27328 1820 27334
rect 1768 27270 1820 27276
rect 1676 26852 1728 26858
rect 1676 26794 1728 26800
rect 1584 26512 1636 26518
rect 1584 26454 1636 26460
rect 1596 24954 1624 26454
rect 1492 24948 1544 24954
rect 1492 24890 1544 24896
rect 1584 24948 1636 24954
rect 1584 24890 1636 24896
rect 1490 23896 1546 23905
rect 1490 23831 1492 23840
rect 1544 23831 1546 23840
rect 1492 23802 1544 23808
rect 1398 23216 1454 23225
rect 1398 23151 1400 23160
rect 1452 23151 1454 23160
rect 1400 23122 1452 23128
rect 1688 22982 1716 26794
rect 1676 22976 1728 22982
rect 1676 22918 1728 22924
rect 1398 22536 1454 22545
rect 1398 22471 1400 22480
rect 1452 22471 1454 22480
rect 1400 22442 1452 22448
rect 1490 21176 1546 21185
rect 1490 21111 1492 21120
rect 1544 21111 1546 21120
rect 1492 21082 1544 21088
rect 1584 21004 1636 21010
rect 1584 20946 1636 20952
rect 1398 20496 1454 20505
rect 1398 20431 1454 20440
rect 1412 20398 1440 20431
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1596 20058 1624 20946
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1400 19304 1452 19310
rect 1400 19246 1452 19252
rect 1412 19145 1440 19246
rect 1584 19168 1636 19174
rect 1398 19136 1454 19145
rect 1584 19110 1636 19116
rect 1398 19071 1454 19080
rect 1412 18970 1440 19071
rect 1596 18970 1624 19110
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1398 18456 1454 18465
rect 1398 18391 1454 18400
rect 1412 18222 1440 18391
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1398 17776 1454 17785
rect 1398 17711 1400 17720
rect 1452 17711 1454 17720
rect 1400 17682 1452 17688
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 16425 1440 16594
rect 1584 16448 1636 16454
rect 1398 16416 1454 16425
rect 1584 16390 1636 16396
rect 1398 16351 1454 16360
rect 1412 16250 1440 16351
rect 1596 16250 1624 16390
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1584 15700 1636 15706
rect 1412 15570 1440 15671
rect 1584 15642 1636 15648
rect 1596 15609 1624 15642
rect 1582 15600 1638 15609
rect 1400 15564 1452 15570
rect 1582 15535 1638 15544
rect 1400 15506 1452 15512
rect 1412 15162 1440 15506
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 14385 1440 14418
rect 1398 14376 1454 14385
rect 1398 14311 1454 14320
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1412 13705 1440 13806
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1584 13456 1636 13462
rect 1584 13398 1636 13404
rect 1398 13016 1454 13025
rect 1398 12951 1454 12960
rect 1412 12850 1440 12951
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1398 11656 1454 11665
rect 1398 11591 1400 11600
rect 1452 11591 1454 11600
rect 1400 11562 1452 11568
rect 1492 11008 1544 11014
rect 1490 10976 1492 10985
rect 1544 10976 1546 10985
rect 1490 10911 1546 10920
rect 1492 9920 1544 9926
rect 1492 9862 1544 9868
rect 1504 9625 1532 9862
rect 1490 9616 1546 9625
rect 1490 9551 1546 9560
rect 1504 9518 1532 9551
rect 1492 9512 1544 9518
rect 1492 9454 1544 9460
rect 1398 8936 1454 8945
rect 1398 8871 1400 8880
rect 1452 8871 1454 8880
rect 1400 8842 1452 8848
rect 1492 8288 1544 8294
rect 1490 8256 1492 8265
rect 1544 8256 1546 8265
rect 1490 8191 1546 8200
rect 1596 8106 1624 13398
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1504 8078 1624 8106
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1412 6905 1440 7278
rect 1504 7002 1532 8078
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 7002 1624 7142
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1398 6896 1454 6905
rect 1688 6882 1716 13126
rect 1398 6831 1454 6840
rect 1596 6854 1716 6882
rect 1596 6254 1624 6854
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1584 6248 1636 6254
rect 1398 6216 1454 6225
rect 1584 6190 1636 6196
rect 1398 6151 1400 6160
rect 1452 6151 1454 6160
rect 1400 6122 1452 6128
rect 1584 5296 1636 5302
rect 1584 5238 1636 5244
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4865 1440 4966
rect 1398 4856 1454 4865
rect 1398 4791 1454 4800
rect 1412 4758 1440 4791
rect 1400 4752 1452 4758
rect 1400 4694 1452 4700
rect 1398 4176 1454 4185
rect 1398 4111 1400 4120
rect 1452 4111 1454 4120
rect 1400 4082 1452 4088
rect 1596 4078 1624 5238
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1308 4004 1360 4010
rect 1308 3946 1360 3952
rect 480 3460 532 3466
rect 480 3402 532 3408
rect 492 800 520 3402
rect 940 2508 992 2514
rect 940 2450 992 2456
rect 952 800 980 2450
rect 1320 1986 1348 3946
rect 1398 3496 1454 3505
rect 1398 3431 1454 3440
rect 1412 2990 1440 3431
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1320 1958 1440 1986
rect 1412 800 1440 1958
rect 1504 1465 1532 3334
rect 1688 2582 1716 6734
rect 1780 5846 1808 27270
rect 2240 26518 2268 27474
rect 2228 26512 2280 26518
rect 2228 26454 2280 26460
rect 2332 26450 2360 29200
rect 2594 28656 2650 28665
rect 2594 28591 2650 28600
rect 2608 26586 2636 28591
rect 2792 27606 2820 29200
rect 2870 27976 2926 27985
rect 2870 27911 2926 27920
rect 2780 27600 2832 27606
rect 2780 27542 2832 27548
rect 2884 26926 2912 27911
rect 3252 27674 3280 29200
rect 3240 27668 3292 27674
rect 3240 27610 3292 27616
rect 3240 27532 3292 27538
rect 3240 27474 3292 27480
rect 3884 27532 3936 27538
rect 3884 27474 3936 27480
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 2596 26580 2648 26586
rect 2596 26522 2648 26528
rect 2320 26444 2372 26450
rect 2320 26386 2372 26392
rect 2332 26042 2360 26386
rect 3252 26042 3280 27474
rect 3896 27062 3924 27474
rect 3884 27056 3936 27062
rect 3884 26998 3936 27004
rect 3332 26852 3384 26858
rect 3332 26794 3384 26800
rect 3344 26489 3372 26794
rect 4172 26518 4200 29200
rect 4436 27328 4488 27334
rect 4436 27270 4488 27276
rect 4252 27056 4304 27062
rect 4252 26998 4304 27004
rect 4160 26512 4212 26518
rect 3330 26480 3386 26489
rect 4160 26454 4212 26460
rect 3330 26415 3386 26424
rect 2320 26036 2372 26042
rect 2320 25978 2372 25984
rect 3240 26036 3292 26042
rect 3240 25978 3292 25984
rect 2504 25832 2556 25838
rect 2504 25774 2556 25780
rect 2136 23520 2188 23526
rect 2136 23462 2188 23468
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 1860 12640 1912 12646
rect 1860 12582 1912 12588
rect 1768 5840 1820 5846
rect 1768 5782 1820 5788
rect 1676 2576 1728 2582
rect 1676 2518 1728 2524
rect 1872 1970 1900 12582
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1964 4078 1992 6598
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 2056 3670 2084 18566
rect 2148 13802 2176 23462
rect 2516 20058 2544 25774
rect 3344 25498 3372 26415
rect 3516 26036 3568 26042
rect 3516 25978 3568 25984
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3528 24138 3556 25978
rect 3516 24132 3568 24138
rect 3516 24074 3568 24080
rect 4160 23180 4212 23186
rect 4160 23122 4212 23128
rect 4172 22778 4200 23122
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2504 20052 2556 20058
rect 2504 19994 2556 20000
rect 2700 19922 2728 20198
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2332 19514 2360 19858
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3988 19514 4016 19654
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 3976 19508 4028 19514
rect 3976 19450 4028 19456
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 18426 2268 19246
rect 4172 18766 4200 22714
rect 2504 18760 2556 18766
rect 2504 18702 2556 18708
rect 4160 18760 4212 18766
rect 4160 18702 4212 18708
rect 2516 18426 2544 18702
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2504 18420 2556 18426
rect 2504 18362 2556 18368
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 17542 2268 17682
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 2240 12238 2268 17478
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2424 13530 2452 13670
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2516 13462 2544 18362
rect 2504 13456 2556 13462
rect 2504 13398 2556 13404
rect 2516 13326 2544 13398
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2240 10470 2268 11562
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2424 4826 2452 13194
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2516 6934 2544 8230
rect 2504 6928 2556 6934
rect 2504 6870 2556 6876
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2044 3664 2096 3670
rect 2044 3606 2096 3612
rect 2424 2990 2452 4762
rect 4264 4282 4292 26998
rect 4448 26518 4476 27270
rect 4632 26926 4660 29200
rect 5552 27606 5580 29200
rect 5724 28008 5776 28014
rect 5724 27950 5776 27956
rect 5736 27606 5764 27950
rect 5540 27600 5592 27606
rect 5540 27542 5592 27548
rect 5724 27600 5776 27606
rect 5724 27542 5776 27548
rect 5172 27532 5224 27538
rect 5172 27474 5224 27480
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4632 26586 4660 26862
rect 4908 26858 4936 27406
rect 4896 26852 4948 26858
rect 4896 26794 4948 26800
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4436 26512 4488 26518
rect 4436 26454 4488 26460
rect 4528 26512 4580 26518
rect 4528 26454 4580 26460
rect 4436 26308 4488 26314
rect 4436 26250 4488 26256
rect 4448 26042 4476 26250
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4540 20602 4568 26454
rect 4908 25838 4936 26794
rect 5184 25974 5212 27474
rect 6012 27062 6040 29200
rect 6000 27056 6052 27062
rect 6000 26998 6052 27004
rect 6472 26994 6500 29200
rect 6920 27396 6972 27402
rect 6920 27338 6972 27344
rect 6932 27062 6960 27338
rect 6920 27056 6972 27062
rect 6920 26998 6972 27004
rect 5724 26988 5776 26994
rect 5724 26930 5776 26936
rect 6460 26988 6512 26994
rect 6460 26930 6512 26936
rect 5736 26586 5764 26930
rect 7392 26926 7420 29200
rect 7852 27606 7880 29200
rect 8024 27940 8076 27946
rect 8024 27882 8076 27888
rect 8036 27674 8064 27882
rect 8024 27668 8076 27674
rect 8024 27610 8076 27616
rect 8116 27668 8168 27674
rect 8116 27610 8168 27616
rect 7840 27600 7892 27606
rect 7840 27542 7892 27548
rect 8128 26994 8156 27610
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7392 26586 7420 26862
rect 7932 26852 7984 26858
rect 7932 26794 7984 26800
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 5172 25968 5224 25974
rect 5172 25910 5224 25916
rect 4896 25832 4948 25838
rect 4896 25774 4948 25780
rect 4908 23118 4936 25774
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2412 2984 2464 2990
rect 2412 2926 2464 2932
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 1860 1964 1912 1970
rect 1860 1906 1912 1912
rect 1490 1456 1546 1465
rect 1490 1391 1546 1400
rect 2332 800 2360 2858
rect 2608 2145 2636 3334
rect 3160 2990 3188 3878
rect 4264 3670 4292 4218
rect 4252 3664 4304 3670
rect 4252 3606 4304 3612
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 2780 2916 2832 2922
rect 2780 2858 2832 2864
rect 2594 2136 2650 2145
rect 2594 2071 2650 2080
rect 2792 800 2820 2858
rect 3252 2514 3280 3334
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 3240 2508 3292 2514
rect 3240 2450 3292 2456
rect 3252 800 3280 2450
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3804 1698 3832 2246
rect 3792 1692 3844 1698
rect 3792 1634 3844 1640
rect 4172 800 4200 2858
rect 4632 800 4660 2858
rect 5184 2417 5212 25910
rect 5736 25770 5764 26522
rect 7944 26518 7972 26794
rect 8024 26784 8076 26790
rect 8024 26726 8076 26732
rect 7932 26512 7984 26518
rect 7932 26454 7984 26460
rect 6368 26240 6420 26246
rect 6368 26182 6420 26188
rect 6380 25906 6408 26182
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 5724 25764 5776 25770
rect 5724 25706 5776 25712
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 2990 6500 3334
rect 7024 3194 7052 19382
rect 8036 17134 8064 26726
rect 8128 26586 8156 26930
rect 8772 26926 8800 29200
rect 8852 26988 8904 26994
rect 8852 26930 8904 26936
rect 8760 26920 8812 26926
rect 8760 26862 8812 26868
rect 8772 26586 8800 26862
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8864 25974 8892 26930
rect 9232 26518 9260 29200
rect 9404 27872 9456 27878
rect 9404 27814 9456 27820
rect 9416 26926 9444 27814
rect 9692 27606 9720 29200
rect 10612 27606 10640 29200
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 10600 27600 10652 27606
rect 10600 27542 10652 27548
rect 10416 27532 10468 27538
rect 10416 27474 10468 27480
rect 9864 27328 9916 27334
rect 9864 27270 9916 27276
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9220 26512 9272 26518
rect 9220 26454 9272 26460
rect 8852 25968 8904 25974
rect 8852 25910 8904 25916
rect 9416 25498 9444 26862
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 26518 9720 26726
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9680 26512 9732 26518
rect 9680 26454 9732 26460
rect 9784 25838 9812 26522
rect 9772 25832 9824 25838
rect 9772 25774 9824 25780
rect 9876 25702 9904 27270
rect 10324 26920 10376 26926
rect 10324 26862 10376 26868
rect 10336 26586 10364 26862
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10232 26444 10284 26450
rect 10232 26386 10284 26392
rect 10244 25974 10272 26386
rect 10232 25968 10284 25974
rect 10232 25910 10284 25916
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9404 25492 9456 25498
rect 9404 25434 9456 25440
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 8772 19310 8800 19858
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16658 8524 16934
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8496 16046 8524 16594
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8300 15972 8352 15978
rect 8300 15914 8352 15920
rect 7012 3188 7064 3194
rect 7012 3130 7064 3136
rect 6460 2984 6512 2990
rect 5722 2952 5778 2961
rect 6460 2926 6512 2932
rect 5722 2887 5724 2896
rect 5776 2887 5778 2896
rect 5724 2858 5776 2864
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5170 2408 5226 2417
rect 5170 2343 5226 2352
rect 5552 800 5580 2450
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5736 1766 5764 2246
rect 5724 1760 5776 1766
rect 5724 1702 5776 1708
rect 6012 800 6040 2314
rect 6472 800 6500 2926
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7392 2514 7420 2790
rect 8312 2582 8340 15914
rect 8680 3194 8708 19246
rect 9220 9104 9272 9110
rect 9220 9046 9272 9052
rect 9232 8634 9260 9046
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9600 8430 9628 8570
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9220 3596 9272 3602
rect 9220 3538 9272 3544
rect 8668 3188 8720 3194
rect 8668 3130 8720 3136
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8772 2650 8800 2926
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7392 800 7420 2450
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7576 1630 7604 2246
rect 7564 1624 7616 1630
rect 7564 1566 7616 1572
rect 7852 800 7880 2314
rect 8772 800 8800 2586
rect 9232 800 9260 3538
rect 9692 3194 9720 8230
rect 10244 4554 10272 25910
rect 10428 24486 10456 27474
rect 10588 27228 10884 27248
rect 10644 27226 10668 27228
rect 10724 27226 10748 27228
rect 10804 27226 10828 27228
rect 10666 27174 10668 27226
rect 10730 27174 10742 27226
rect 10804 27174 10806 27226
rect 10644 27172 10668 27174
rect 10724 27172 10748 27174
rect 10804 27172 10828 27174
rect 10588 27152 10884 27172
rect 11072 27146 11100 29200
rect 11992 27606 12020 29200
rect 12452 27606 12480 29200
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 12440 27600 12492 27606
rect 12440 27542 12492 27548
rect 11072 27118 11192 27146
rect 11058 27024 11114 27033
rect 11058 26959 11114 26968
rect 11072 26790 11100 26959
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 11164 26450 11192 27118
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 11256 26518 11284 26930
rect 11992 26926 12020 27542
rect 12912 26926 12940 29200
rect 13832 27674 13860 29200
rect 13820 27668 13872 27674
rect 13820 27610 13872 27616
rect 13544 27532 13596 27538
rect 13544 27474 13596 27480
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 11244 26512 11296 26518
rect 11244 26454 11296 26460
rect 11152 26444 11204 26450
rect 11152 26386 11204 26392
rect 10588 26140 10884 26160
rect 10644 26138 10668 26140
rect 10724 26138 10748 26140
rect 10804 26138 10828 26140
rect 10666 26086 10668 26138
rect 10730 26086 10742 26138
rect 10804 26086 10806 26138
rect 10644 26084 10668 26086
rect 10724 26084 10748 26086
rect 10804 26084 10828 26086
rect 10588 26064 10884 26084
rect 11256 25974 11284 26454
rect 11520 26240 11572 26246
rect 11520 26182 11572 26188
rect 11244 25968 11296 25974
rect 11244 25910 11296 25916
rect 10588 25052 10884 25072
rect 10644 25050 10668 25052
rect 10724 25050 10748 25052
rect 10804 25050 10828 25052
rect 10666 24998 10668 25050
rect 10730 24998 10742 25050
rect 10804 24998 10806 25050
rect 10644 24996 10668 24998
rect 10724 24996 10748 24998
rect 10804 24996 10828 24998
rect 10588 24976 10884 24996
rect 10336 24458 10456 24486
rect 10336 16794 10364 24458
rect 10588 23964 10884 23984
rect 10644 23962 10668 23964
rect 10724 23962 10748 23964
rect 10804 23962 10828 23964
rect 10666 23910 10668 23962
rect 10730 23910 10742 23962
rect 10804 23910 10806 23962
rect 10644 23908 10668 23910
rect 10724 23908 10748 23910
rect 10804 23908 10828 23910
rect 10588 23888 10884 23908
rect 10588 22876 10884 22896
rect 10644 22874 10668 22876
rect 10724 22874 10748 22876
rect 10804 22874 10828 22876
rect 10666 22822 10668 22874
rect 10730 22822 10742 22874
rect 10804 22822 10806 22874
rect 10644 22820 10668 22822
rect 10724 22820 10748 22822
rect 10804 22820 10828 22822
rect 10588 22800 10884 22820
rect 10588 21788 10884 21808
rect 10644 21786 10668 21788
rect 10724 21786 10748 21788
rect 10804 21786 10828 21788
rect 10666 21734 10668 21786
rect 10730 21734 10742 21786
rect 10804 21734 10806 21786
rect 10644 21732 10668 21734
rect 10724 21732 10748 21734
rect 10804 21732 10828 21734
rect 10588 21712 10884 21732
rect 10588 20700 10884 20720
rect 10644 20698 10668 20700
rect 10724 20698 10748 20700
rect 10804 20698 10828 20700
rect 10666 20646 10668 20698
rect 10730 20646 10742 20698
rect 10804 20646 10806 20698
rect 10644 20644 10668 20646
rect 10724 20644 10748 20646
rect 10804 20644 10828 20646
rect 10588 20624 10884 20644
rect 10588 19612 10884 19632
rect 10644 19610 10668 19612
rect 10724 19610 10748 19612
rect 10804 19610 10828 19612
rect 10666 19558 10668 19610
rect 10730 19558 10742 19610
rect 10804 19558 10806 19610
rect 10644 19556 10668 19558
rect 10724 19556 10748 19558
rect 10804 19556 10828 19558
rect 10588 19536 10884 19556
rect 10588 18524 10884 18544
rect 10644 18522 10668 18524
rect 10724 18522 10748 18524
rect 10804 18522 10828 18524
rect 10666 18470 10668 18522
rect 10730 18470 10742 18522
rect 10804 18470 10806 18522
rect 10644 18468 10668 18470
rect 10724 18468 10748 18470
rect 10804 18468 10828 18470
rect 10588 18448 10884 18468
rect 10588 17436 10884 17456
rect 10644 17434 10668 17436
rect 10724 17434 10748 17436
rect 10804 17434 10828 17436
rect 10666 17382 10668 17434
rect 10730 17382 10742 17434
rect 10804 17382 10806 17434
rect 10644 17380 10668 17382
rect 10724 17380 10748 17382
rect 10804 17380 10828 17382
rect 10588 17360 10884 17380
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10588 16348 10884 16368
rect 10644 16346 10668 16348
rect 10724 16346 10748 16348
rect 10804 16346 10828 16348
rect 10666 16294 10668 16346
rect 10730 16294 10742 16346
rect 10804 16294 10806 16346
rect 10644 16292 10668 16294
rect 10724 16292 10748 16294
rect 10804 16292 10828 16294
rect 10588 16272 10884 16292
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 10336 4282 10364 15438
rect 10588 15260 10884 15280
rect 10644 15258 10668 15260
rect 10724 15258 10748 15260
rect 10804 15258 10828 15260
rect 10666 15206 10668 15258
rect 10730 15206 10742 15258
rect 10804 15206 10806 15258
rect 10644 15204 10668 15206
rect 10724 15204 10748 15206
rect 10804 15204 10828 15206
rect 10588 15184 10884 15204
rect 10588 14172 10884 14192
rect 10644 14170 10668 14172
rect 10724 14170 10748 14172
rect 10804 14170 10828 14172
rect 10666 14118 10668 14170
rect 10730 14118 10742 14170
rect 10804 14118 10806 14170
rect 10644 14116 10668 14118
rect 10724 14116 10748 14118
rect 10804 14116 10828 14118
rect 10588 14096 10884 14116
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10612 13462 10640 13806
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10520 12986 10548 13330
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10588 13084 10884 13104
rect 10644 13082 10668 13084
rect 10724 13082 10748 13084
rect 10804 13082 10828 13084
rect 10666 13030 10668 13082
rect 10730 13030 10742 13082
rect 10804 13030 10806 13082
rect 10644 13028 10668 13030
rect 10724 13028 10748 13030
rect 10804 13028 10828 13030
rect 10588 13008 10884 13028
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10588 11996 10884 12016
rect 10644 11994 10668 11996
rect 10724 11994 10748 11996
rect 10804 11994 10828 11996
rect 10666 11942 10668 11994
rect 10730 11942 10742 11994
rect 10804 11942 10806 11994
rect 10644 11940 10668 11942
rect 10724 11940 10748 11942
rect 10804 11940 10828 11942
rect 10588 11920 10884 11940
rect 10588 10908 10884 10928
rect 10644 10906 10668 10908
rect 10724 10906 10748 10908
rect 10804 10906 10828 10908
rect 10666 10854 10668 10906
rect 10730 10854 10742 10906
rect 10804 10854 10806 10906
rect 10644 10852 10668 10854
rect 10724 10852 10748 10854
rect 10804 10852 10828 10854
rect 10588 10832 10884 10852
rect 10588 9820 10884 9840
rect 10644 9818 10668 9820
rect 10724 9818 10748 9820
rect 10804 9818 10828 9820
rect 10666 9766 10668 9818
rect 10730 9766 10742 9818
rect 10804 9766 10806 9818
rect 10644 9764 10668 9766
rect 10724 9764 10748 9766
rect 10804 9764 10828 9766
rect 10588 9744 10884 9764
rect 10588 8732 10884 8752
rect 10644 8730 10668 8732
rect 10724 8730 10748 8732
rect 10804 8730 10828 8732
rect 10666 8678 10668 8730
rect 10730 8678 10742 8730
rect 10804 8678 10806 8730
rect 10644 8676 10668 8678
rect 10724 8676 10748 8678
rect 10804 8676 10828 8678
rect 10588 8656 10884 8676
rect 10588 7644 10884 7664
rect 10644 7642 10668 7644
rect 10724 7642 10748 7644
rect 10804 7642 10828 7644
rect 10666 7590 10668 7642
rect 10730 7590 10742 7642
rect 10804 7590 10806 7642
rect 10644 7588 10668 7590
rect 10724 7588 10748 7590
rect 10804 7588 10828 7590
rect 10588 7568 10884 7588
rect 10588 6556 10884 6576
rect 10644 6554 10668 6556
rect 10724 6554 10748 6556
rect 10804 6554 10828 6556
rect 10666 6502 10668 6554
rect 10730 6502 10742 6554
rect 10804 6502 10806 6554
rect 10644 6500 10668 6502
rect 10724 6500 10748 6502
rect 10804 6500 10828 6502
rect 10588 6480 10884 6500
rect 10588 5468 10884 5488
rect 10644 5466 10668 5468
rect 10724 5466 10748 5468
rect 10804 5466 10828 5468
rect 10666 5414 10668 5466
rect 10730 5414 10742 5466
rect 10804 5414 10806 5466
rect 10644 5412 10668 5414
rect 10724 5412 10748 5414
rect 10804 5412 10828 5414
rect 10588 5392 10884 5412
rect 10588 4380 10884 4400
rect 10644 4378 10668 4380
rect 10724 4378 10748 4380
rect 10804 4378 10828 4380
rect 10666 4326 10668 4378
rect 10730 4326 10742 4378
rect 10804 4326 10806 4378
rect 10644 4324 10668 4326
rect 10724 4324 10748 4326
rect 10804 4324 10828 4326
rect 10588 4304 10884 4324
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9680 2984 9732 2990
rect 9680 2926 9732 2932
rect 9692 800 9720 2926
rect 10336 2582 10364 4218
rect 11072 3670 11100 13262
rect 11532 3738 11560 26182
rect 12268 25430 12296 26726
rect 12912 26353 12940 26726
rect 12898 26344 12954 26353
rect 12898 26279 12954 26288
rect 12912 25974 12940 26279
rect 13556 26246 13584 27474
rect 14292 26926 14320 29200
rect 14752 27606 14780 29200
rect 14740 27600 14792 27606
rect 14740 27542 14792 27548
rect 15016 27532 15068 27538
rect 15016 27474 15068 27480
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14464 26784 14516 26790
rect 14464 26726 14516 26732
rect 14476 26518 14504 26726
rect 14464 26512 14516 26518
rect 14464 26454 14516 26460
rect 14188 26308 14240 26314
rect 14188 26250 14240 26256
rect 13544 26240 13596 26246
rect 14200 26217 14228 26250
rect 15028 26246 15056 27474
rect 15672 26926 15700 29200
rect 16132 27606 16160 29200
rect 17052 28150 17080 29200
rect 17040 28144 17092 28150
rect 17040 28086 17092 28092
rect 16488 28076 16540 28082
rect 16488 28018 16540 28024
rect 16500 27606 16528 28018
rect 17408 28008 17460 28014
rect 17408 27950 17460 27956
rect 16120 27600 16172 27606
rect 16120 27542 16172 27548
rect 16488 27600 16540 27606
rect 16488 27542 16540 27548
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15660 26920 15712 26926
rect 15660 26862 15712 26868
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15016 26240 15068 26246
rect 13544 26182 13596 26188
rect 14186 26208 14242 26217
rect 12900 25968 12952 25974
rect 12900 25910 12952 25916
rect 12256 25424 12308 25430
rect 12256 25366 12308 25372
rect 13556 16522 13584 26182
rect 15016 26182 15068 26188
rect 14186 26143 14242 26152
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 13544 16516 13596 16522
rect 13544 16458 13596 16464
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13870 13768 14214
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13740 13462 13768 13806
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 13190 11928 13330
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12170 11928 13126
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10324 2576 10376 2582
rect 10324 2518 10376 2524
rect 10520 2514 10548 3334
rect 10588 3292 10884 3312
rect 10644 3290 10668 3292
rect 10724 3290 10748 3292
rect 10804 3290 10828 3292
rect 10666 3238 10668 3290
rect 10730 3238 10742 3290
rect 10804 3238 10806 3290
rect 10644 3236 10668 3238
rect 10724 3236 10748 3238
rect 10804 3236 10828 3238
rect 10588 3216 10884 3236
rect 11532 2990 11560 3674
rect 13268 3392 13320 3398
rect 13268 3334 13320 3340
rect 13280 2990 13308 3334
rect 13740 3194 13768 8434
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 10520 1986 10548 2450
rect 10588 2204 10884 2224
rect 10644 2202 10668 2204
rect 10724 2202 10748 2204
rect 10804 2202 10828 2204
rect 10666 2150 10668 2202
rect 10730 2150 10742 2202
rect 10804 2150 10806 2202
rect 10644 2148 10668 2150
rect 10724 2148 10748 2150
rect 10804 2148 10828 2150
rect 10588 2128 10884 2148
rect 10520 1958 10640 1986
rect 10612 800 10640 1958
rect 10980 1442 11008 2790
rect 11992 2514 12020 2790
rect 12176 2689 12204 2858
rect 12162 2680 12218 2689
rect 12162 2615 12218 2624
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 10980 1414 11100 1442
rect 11072 800 11100 1414
rect 11992 800 12020 2450
rect 12348 2304 12400 2310
rect 12348 2246 12400 2252
rect 12360 1834 12388 2246
rect 12348 1828 12400 1834
rect 12348 1770 12400 1776
rect 12452 800 12480 2586
rect 12912 800 12940 2858
rect 13096 2106 13124 2926
rect 13740 2446 13768 3130
rect 13832 2582 13860 13738
rect 14384 3738 14412 16526
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 14200 2514 14228 3130
rect 14280 2916 14332 2922
rect 14280 2858 14332 2864
rect 14188 2508 14240 2514
rect 14188 2450 14240 2456
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13820 2304 13872 2310
rect 13820 2246 13872 2252
rect 13084 2100 13136 2106
rect 13084 2042 13136 2048
rect 13740 1562 13768 2246
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13832 800 13860 2246
rect 14292 800 14320 2858
rect 14384 2650 14412 3334
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14476 2650 14504 2858
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 15028 2590 15056 26182
rect 15476 15972 15528 15978
rect 15476 15914 15528 15920
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 14936 2562 15056 2590
rect 14936 1902 14964 2562
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 15212 800 15240 4014
rect 15488 3738 15516 15914
rect 15580 13530 15608 26726
rect 15672 26586 15700 26862
rect 15660 26580 15712 26586
rect 15660 26522 15712 26528
rect 15856 20058 15884 27474
rect 17420 27470 17448 27950
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17512 27418 17540 29200
rect 17972 27606 18000 29200
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 18616 27538 18644 28086
rect 17684 27532 17736 27538
rect 17684 27474 17736 27480
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 18604 27532 18656 27538
rect 18604 27474 18656 27480
rect 16948 27056 17000 27062
rect 16948 26998 17000 27004
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 16764 26920 16816 26926
rect 16764 26862 16816 26868
rect 16408 25974 16436 26862
rect 16776 26450 16804 26862
rect 16960 26450 16988 26998
rect 17052 26586 17080 27406
rect 17512 27390 17632 27418
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17500 27328 17552 27334
rect 17500 27270 17552 27276
rect 17144 26586 17172 27270
rect 17512 26858 17540 27270
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16948 26444 17000 26450
rect 16948 26386 17000 26392
rect 16396 25968 16448 25974
rect 16396 25910 16448 25916
rect 16776 25498 16804 26386
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 16960 25906 16988 26182
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 17604 25838 17632 27390
rect 17696 27062 17724 27474
rect 17684 27056 17736 27062
rect 17684 26998 17736 27004
rect 17684 26852 17736 26858
rect 17684 26794 17736 26800
rect 17696 25974 17724 26794
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17788 26450 17816 26522
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 17880 26382 17908 27474
rect 17960 27056 18012 27062
rect 17960 26998 18012 27004
rect 17868 26376 17920 26382
rect 17868 26318 17920 26324
rect 17684 25968 17736 25974
rect 17684 25910 17736 25916
rect 17592 25832 17644 25838
rect 17592 25774 17644 25780
rect 17604 25498 17632 25774
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 17592 25492 17644 25498
rect 17592 25434 17644 25440
rect 16776 25362 16804 25434
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16224 19378 16252 19790
rect 16212 19372 16264 19378
rect 16212 19314 16264 19320
rect 17696 14346 17724 25910
rect 17880 16182 17908 26318
rect 17972 25430 18000 26998
rect 18052 26852 18104 26858
rect 18052 26794 18104 26800
rect 18064 26246 18092 26794
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 18616 25974 18644 27474
rect 18892 26450 18920 29200
rect 18972 28144 19024 28150
rect 18972 28086 19024 28092
rect 18984 26586 19012 28086
rect 19352 27606 19380 29200
rect 20272 27962 20300 29200
rect 20088 27934 20300 27962
rect 20628 28008 20680 28014
rect 20628 27950 20680 27956
rect 19340 27600 19392 27606
rect 19340 27542 19392 27548
rect 19800 27532 19852 27538
rect 19800 27474 19852 27480
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 18972 26580 19024 26586
rect 18972 26522 19024 26528
rect 18880 26444 18932 26450
rect 18880 26386 18932 26392
rect 18984 25974 19012 26522
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 17960 25424 18012 25430
rect 17960 25366 18012 25372
rect 19076 20622 19104 26794
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 19524 26240 19576 26246
rect 19524 26182 19576 26188
rect 19536 25974 19564 26182
rect 19524 25968 19576 25974
rect 19524 25910 19576 25916
rect 19628 25906 19656 26726
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 18984 20594 19104 20622
rect 19628 20622 19656 25842
rect 19812 21690 19840 27474
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19892 26308 19944 26314
rect 19892 26250 19944 26256
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19904 20622 19932 26250
rect 19996 21690 20024 27066
rect 20088 26518 20116 27934
rect 20220 27772 20516 27792
rect 20276 27770 20300 27772
rect 20356 27770 20380 27772
rect 20436 27770 20460 27772
rect 20298 27718 20300 27770
rect 20362 27718 20374 27770
rect 20436 27718 20438 27770
rect 20276 27716 20300 27718
rect 20356 27716 20380 27718
rect 20436 27716 20460 27718
rect 20220 27696 20516 27716
rect 20640 27606 20668 27950
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 20260 27532 20312 27538
rect 20260 27474 20312 27480
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20536 27532 20588 27538
rect 20536 27474 20588 27480
rect 20272 26858 20300 27474
rect 20456 26926 20484 27474
rect 20548 27130 20576 27474
rect 20732 27470 20760 29200
rect 20720 27464 20772 27470
rect 20720 27406 20772 27412
rect 20536 27124 20588 27130
rect 20536 27066 20588 27072
rect 20444 26920 20496 26926
rect 21088 26920 21140 26926
rect 20994 26888 21050 26897
rect 20496 26868 20576 26874
rect 20444 26862 20576 26868
rect 20260 26852 20312 26858
rect 20456 26846 20576 26862
rect 20260 26794 20312 26800
rect 20220 26684 20516 26704
rect 20276 26682 20300 26684
rect 20356 26682 20380 26684
rect 20436 26682 20460 26684
rect 20298 26630 20300 26682
rect 20362 26630 20374 26682
rect 20436 26630 20438 26682
rect 20276 26628 20300 26630
rect 20356 26628 20380 26630
rect 20436 26628 20460 26630
rect 20220 26608 20516 26628
rect 20076 26512 20128 26518
rect 20076 26454 20128 26460
rect 20548 25838 20576 26846
rect 21088 26862 21140 26868
rect 20994 26823 21050 26832
rect 21008 26790 21036 26823
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20996 26784 21048 26790
rect 20996 26726 21048 26732
rect 20732 26586 20760 26726
rect 20720 26580 20772 26586
rect 20720 26522 20772 26528
rect 21100 26353 21128 26862
rect 21192 26518 21220 29200
rect 22112 27538 22140 29200
rect 22100 27532 22152 27538
rect 22100 27474 22152 27480
rect 22572 27062 22600 29200
rect 22284 27056 22336 27062
rect 22284 26998 22336 27004
rect 22560 27056 22612 27062
rect 22560 26998 22612 27004
rect 21180 26512 21232 26518
rect 21180 26454 21232 26460
rect 22296 26450 22324 26998
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 23492 26908 23520 29200
rect 23952 27606 23980 29200
rect 24308 28076 24360 28082
rect 24308 28018 24360 28024
rect 23940 27600 23992 27606
rect 23940 27542 23992 27548
rect 23756 27532 23808 27538
rect 23756 27474 23808 27480
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 23572 26920 23624 26926
rect 23492 26880 23572 26908
rect 22744 26852 22796 26858
rect 22744 26794 22796 26800
rect 22284 26444 22336 26450
rect 22284 26386 22336 26392
rect 21086 26344 21142 26353
rect 21086 26279 21142 26288
rect 21100 25838 21128 26279
rect 20536 25832 20588 25838
rect 20536 25774 20588 25780
rect 21088 25832 21140 25838
rect 21088 25774 21140 25780
rect 20220 25596 20516 25616
rect 20276 25594 20300 25596
rect 20356 25594 20380 25596
rect 20436 25594 20460 25596
rect 20298 25542 20300 25594
rect 20362 25542 20374 25594
rect 20436 25542 20438 25594
rect 20276 25540 20300 25542
rect 20356 25540 20380 25542
rect 20436 25540 20460 25542
rect 20220 25520 20516 25540
rect 20220 24508 20516 24528
rect 20276 24506 20300 24508
rect 20356 24506 20380 24508
rect 20436 24506 20460 24508
rect 20298 24454 20300 24506
rect 20362 24454 20374 24506
rect 20436 24454 20438 24506
rect 20276 24452 20300 24454
rect 20356 24452 20380 24454
rect 20436 24452 20460 24454
rect 20220 24432 20516 24452
rect 20220 23420 20516 23440
rect 20276 23418 20300 23420
rect 20356 23418 20380 23420
rect 20436 23418 20460 23420
rect 20298 23366 20300 23418
rect 20362 23366 20374 23418
rect 20436 23366 20438 23418
rect 20276 23364 20300 23366
rect 20356 23364 20380 23366
rect 20436 23364 20460 23366
rect 20220 23344 20516 23364
rect 20220 22332 20516 22352
rect 20276 22330 20300 22332
rect 20356 22330 20380 22332
rect 20436 22330 20460 22332
rect 20298 22278 20300 22330
rect 20362 22278 20374 22330
rect 20436 22278 20438 22330
rect 20276 22276 20300 22278
rect 20356 22276 20380 22278
rect 20436 22276 20460 22278
rect 20220 22256 20516 22276
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20088 21146 20116 21490
rect 20220 21244 20516 21264
rect 20276 21242 20300 21244
rect 20356 21242 20380 21244
rect 20436 21242 20460 21244
rect 20298 21190 20300 21242
rect 20362 21190 20374 21242
rect 20436 21190 20438 21242
rect 20276 21188 20300 21190
rect 20356 21188 20380 21190
rect 20436 21188 20460 21190
rect 20220 21168 20516 21188
rect 20076 21140 20128 21146
rect 20076 21082 20128 21088
rect 20076 21004 20128 21010
rect 20076 20946 20128 20952
rect 19628 20594 19840 20622
rect 19904 20594 20024 20622
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17880 15570 17908 16118
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18800 15570 18828 15982
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 17880 14958 17908 15506
rect 18892 15162 18920 15642
rect 18984 15366 19012 20594
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 17202 19380 19654
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 19352 15470 19380 17138
rect 19352 15442 19472 15470
rect 18972 15360 19024 15366
rect 18972 15302 19024 15308
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14346 18092 14894
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16028 4480 16080 4486
rect 16028 4422 16080 4428
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15396 2990 15424 3538
rect 15488 2990 15516 3674
rect 16040 3097 16068 4422
rect 16500 3670 16528 4422
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16488 3664 16540 3670
rect 16488 3606 16540 3612
rect 16026 3088 16082 3097
rect 16026 3023 16082 3032
rect 16212 3052 16264 3058
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15290 2680 15346 2689
rect 15290 2615 15292 2624
rect 15344 2615 15346 2624
rect 15292 2586 15344 2592
rect 16040 2582 16068 3023
rect 16212 2994 16264 3000
rect 16120 2916 16172 2922
rect 16120 2858 16172 2864
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 15660 2372 15712 2378
rect 15660 2314 15712 2320
rect 15672 800 15700 2314
rect 16132 800 16160 2858
rect 16224 2582 16252 2994
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16684 2514 16712 3946
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16776 3194 16804 3538
rect 16764 3188 16816 3194
rect 16764 3130 16816 3136
rect 16868 2990 16896 5306
rect 18156 5302 18184 14962
rect 18984 13394 19012 15302
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 18144 5296 18196 5302
rect 18144 5238 18196 5244
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17420 3602 17448 3878
rect 17408 3596 17460 3602
rect 17408 3538 17460 3544
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 16856 2984 16908 2990
rect 16856 2926 16908 2932
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 17052 800 17080 3130
rect 17512 2990 17540 3334
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17512 2582 17540 2926
rect 17500 2576 17552 2582
rect 17500 2518 17552 2524
rect 17604 2428 17632 4014
rect 17512 2400 17632 2428
rect 17512 800 17540 2400
rect 17788 2378 17816 4422
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18708 3602 18736 3878
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18156 2582 18184 3402
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17696 1970 17724 2246
rect 17684 1964 17736 1970
rect 17684 1906 17736 1912
rect 18432 800 18460 3538
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 1970 18644 3334
rect 19076 2854 19104 9658
rect 19444 4282 19472 15442
rect 19432 4276 19484 4282
rect 19432 4218 19484 4224
rect 19444 3466 19472 4218
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 19444 3058 19472 3402
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 19628 2990 19656 3334
rect 19812 3194 19840 20594
rect 19996 15502 20024 20594
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19892 13796 19944 13802
rect 19892 13738 19944 13744
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19616 2984 19668 2990
rect 19616 2926 19668 2932
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 18880 2372 18932 2378
rect 18880 2314 18932 2320
rect 18604 1964 18656 1970
rect 18604 1906 18656 1912
rect 18892 800 18920 2314
rect 19352 800 19380 2926
rect 19904 2582 19932 13738
rect 19892 2576 19944 2582
rect 19892 2518 19944 2524
rect 20088 1834 20116 20946
rect 20220 20156 20516 20176
rect 20276 20154 20300 20156
rect 20356 20154 20380 20156
rect 20436 20154 20460 20156
rect 20298 20102 20300 20154
rect 20362 20102 20374 20154
rect 20436 20102 20438 20154
rect 20276 20100 20300 20102
rect 20356 20100 20380 20102
rect 20436 20100 20460 20102
rect 20220 20080 20516 20100
rect 20220 19068 20516 19088
rect 20276 19066 20300 19068
rect 20356 19066 20380 19068
rect 20436 19066 20460 19068
rect 20298 19014 20300 19066
rect 20362 19014 20374 19066
rect 20436 19014 20438 19066
rect 20276 19012 20300 19014
rect 20356 19012 20380 19014
rect 20436 19012 20460 19014
rect 20220 18992 20516 19012
rect 20220 17980 20516 18000
rect 20276 17978 20300 17980
rect 20356 17978 20380 17980
rect 20436 17978 20460 17980
rect 20298 17926 20300 17978
rect 20362 17926 20374 17978
rect 20436 17926 20438 17978
rect 20276 17924 20300 17926
rect 20356 17924 20380 17926
rect 20436 17924 20460 17926
rect 20220 17904 20516 17924
rect 20220 16892 20516 16912
rect 20276 16890 20300 16892
rect 20356 16890 20380 16892
rect 20436 16890 20460 16892
rect 20298 16838 20300 16890
rect 20362 16838 20374 16890
rect 20436 16838 20438 16890
rect 20276 16836 20300 16838
rect 20356 16836 20380 16838
rect 20436 16836 20460 16838
rect 20220 16816 20516 16836
rect 21100 16114 21128 25774
rect 22756 23866 22784 26794
rect 22848 26246 22876 26862
rect 23204 26852 23256 26858
rect 23204 26794 23256 26800
rect 23216 26246 23244 26794
rect 23492 26586 23520 26880
rect 23572 26862 23624 26868
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 23204 26240 23256 26246
rect 23204 26182 23256 26188
rect 22744 23860 22796 23866
rect 22744 23802 22796 23808
rect 22560 23656 22612 23662
rect 22560 23598 22612 23604
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 21192 22574 21220 23122
rect 21548 23044 21600 23050
rect 21548 22986 21600 22992
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 21364 16788 21416 16794
rect 21364 16730 21416 16736
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21192 16454 21220 16594
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 20220 15804 20516 15824
rect 20276 15802 20300 15804
rect 20356 15802 20380 15804
rect 20436 15802 20460 15804
rect 20298 15750 20300 15802
rect 20362 15750 20374 15802
rect 20436 15750 20438 15802
rect 20276 15748 20300 15750
rect 20356 15748 20380 15750
rect 20436 15748 20460 15750
rect 20220 15728 20516 15748
rect 20220 14716 20516 14736
rect 20276 14714 20300 14716
rect 20356 14714 20380 14716
rect 20436 14714 20460 14716
rect 20298 14662 20300 14714
rect 20362 14662 20374 14714
rect 20436 14662 20438 14714
rect 20276 14660 20300 14662
rect 20356 14660 20380 14662
rect 20436 14660 20460 14662
rect 20220 14640 20516 14660
rect 21100 13870 21128 16050
rect 21376 16046 21404 16730
rect 21364 16040 21416 16046
rect 21364 15982 21416 15988
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21192 15502 21220 15642
rect 21376 15570 21404 15982
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 20220 13628 20516 13648
rect 20276 13626 20300 13628
rect 20356 13626 20380 13628
rect 20436 13626 20460 13628
rect 20298 13574 20300 13626
rect 20362 13574 20374 13626
rect 20436 13574 20438 13626
rect 20276 13572 20300 13574
rect 20356 13572 20380 13574
rect 20436 13572 20460 13574
rect 20220 13552 20516 13572
rect 20220 12540 20516 12560
rect 20276 12538 20300 12540
rect 20356 12538 20380 12540
rect 20436 12538 20460 12540
rect 20298 12486 20300 12538
rect 20362 12486 20374 12538
rect 20436 12486 20438 12538
rect 20276 12484 20300 12486
rect 20356 12484 20380 12486
rect 20436 12484 20460 12486
rect 20220 12464 20516 12484
rect 20220 11452 20516 11472
rect 20276 11450 20300 11452
rect 20356 11450 20380 11452
rect 20436 11450 20460 11452
rect 20298 11398 20300 11450
rect 20362 11398 20374 11450
rect 20436 11398 20438 11450
rect 20276 11396 20300 11398
rect 20356 11396 20380 11398
rect 20436 11396 20460 11398
rect 20220 11376 20516 11396
rect 20220 10364 20516 10384
rect 20276 10362 20300 10364
rect 20356 10362 20380 10364
rect 20436 10362 20460 10364
rect 20298 10310 20300 10362
rect 20362 10310 20374 10362
rect 20436 10310 20438 10362
rect 20276 10308 20300 10310
rect 20356 10308 20380 10310
rect 20436 10308 20460 10310
rect 20220 10288 20516 10308
rect 20220 9276 20516 9296
rect 20276 9274 20300 9276
rect 20356 9274 20380 9276
rect 20436 9274 20460 9276
rect 20298 9222 20300 9274
rect 20362 9222 20374 9274
rect 20436 9222 20438 9274
rect 20276 9220 20300 9222
rect 20356 9220 20380 9222
rect 20436 9220 20460 9222
rect 20220 9200 20516 9220
rect 20220 8188 20516 8208
rect 20276 8186 20300 8188
rect 20356 8186 20380 8188
rect 20436 8186 20460 8188
rect 20298 8134 20300 8186
rect 20362 8134 20374 8186
rect 20436 8134 20438 8186
rect 20276 8132 20300 8134
rect 20356 8132 20380 8134
rect 20436 8132 20460 8134
rect 20220 8112 20516 8132
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20220 7100 20516 7120
rect 20276 7098 20300 7100
rect 20356 7098 20380 7100
rect 20436 7098 20460 7100
rect 20298 7046 20300 7098
rect 20362 7046 20374 7098
rect 20436 7046 20438 7098
rect 20276 7044 20300 7046
rect 20356 7044 20380 7046
rect 20436 7044 20460 7046
rect 20220 7024 20516 7044
rect 20220 6012 20516 6032
rect 20276 6010 20300 6012
rect 20356 6010 20380 6012
rect 20436 6010 20460 6012
rect 20298 5958 20300 6010
rect 20362 5958 20374 6010
rect 20436 5958 20438 6010
rect 20276 5956 20300 5958
rect 20356 5956 20380 5958
rect 20436 5956 20460 5958
rect 20220 5936 20516 5956
rect 20220 4924 20516 4944
rect 20276 4922 20300 4924
rect 20356 4922 20380 4924
rect 20436 4922 20460 4924
rect 20298 4870 20300 4922
rect 20362 4870 20374 4922
rect 20436 4870 20438 4922
rect 20276 4868 20300 4870
rect 20356 4868 20380 4870
rect 20436 4868 20460 4870
rect 20220 4848 20516 4868
rect 20536 4480 20588 4486
rect 20536 4422 20588 4428
rect 20220 3836 20516 3856
rect 20276 3834 20300 3836
rect 20356 3834 20380 3836
rect 20436 3834 20460 3836
rect 20298 3782 20300 3834
rect 20362 3782 20374 3834
rect 20436 3782 20438 3834
rect 20276 3780 20300 3782
rect 20356 3780 20380 3782
rect 20436 3780 20460 3782
rect 20220 3760 20516 3780
rect 20548 3398 20576 4422
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20220 2748 20516 2768
rect 20276 2746 20300 2748
rect 20356 2746 20380 2748
rect 20436 2746 20460 2748
rect 20298 2694 20300 2746
rect 20362 2694 20374 2746
rect 20436 2694 20438 2746
rect 20276 2692 20300 2694
rect 20356 2692 20380 2694
rect 20436 2692 20460 2694
rect 20220 2672 20516 2692
rect 20548 2514 20576 3334
rect 20640 2582 20668 7822
rect 21560 4282 21588 22986
rect 22572 20398 22600 23598
rect 22756 22574 22784 23598
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 21928 20058 21956 20334
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 21824 19916 21876 19922
rect 21824 19858 21876 19864
rect 21836 9382 21864 19858
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22756 16658 22784 16730
rect 22744 16652 22796 16658
rect 22744 16594 22796 16600
rect 22008 15972 22060 15978
rect 22008 15914 22060 15920
rect 22020 15706 22048 15914
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21916 5160 21968 5166
rect 21916 5102 21968 5108
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21824 4276 21876 4282
rect 21824 4218 21876 4224
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21192 3602 21220 3878
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 20732 2990 20760 3334
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20628 2576 20680 2582
rect 20628 2518 20680 2524
rect 20536 2508 20588 2514
rect 20536 2450 20588 2456
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20076 1828 20128 1834
rect 20076 1770 20128 1776
rect 20272 800 20300 2314
rect 20732 800 20760 2926
rect 21836 2564 21864 4218
rect 21928 3534 21956 5102
rect 22572 3738 22600 14418
rect 22848 13870 22876 26182
rect 23216 26042 23244 26182
rect 23204 26036 23256 26042
rect 23204 25978 23256 25984
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 23124 23322 23152 24210
rect 23112 23316 23164 23322
rect 23112 23258 23164 23264
rect 23124 23186 23152 23258
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 23124 20398 23152 23122
rect 23112 20392 23164 20398
rect 23112 20334 23164 20340
rect 23216 19530 23244 25978
rect 23584 24750 23612 26726
rect 23768 25838 23796 27474
rect 24136 27130 24164 27474
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 24320 26994 24348 28018
rect 24412 27588 24440 29200
rect 24492 27600 24544 27606
rect 24412 27560 24492 27588
rect 24492 27542 24544 27548
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 25332 26926 25360 29200
rect 25792 27334 25820 29200
rect 25872 27668 25924 27674
rect 25872 27610 25924 27616
rect 25780 27328 25832 27334
rect 25780 27270 25832 27276
rect 25884 27130 25912 27610
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 26332 26920 26384 26926
rect 26332 26862 26384 26868
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24504 26217 24532 26250
rect 24490 26208 24546 26217
rect 24490 26143 24546 26152
rect 23756 25832 23808 25838
rect 23756 25774 23808 25780
rect 23664 25696 23716 25702
rect 23664 25638 23716 25644
rect 23676 25226 23704 25638
rect 23664 25220 23716 25226
rect 23664 25162 23716 25168
rect 23572 24744 23624 24750
rect 23572 24686 23624 24692
rect 23480 24608 23532 24614
rect 23480 24550 23532 24556
rect 23492 24206 23520 24550
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23492 23730 23520 24142
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23768 21622 23796 25774
rect 25976 22574 26004 26726
rect 26344 26518 26372 26862
rect 26608 26852 26660 26858
rect 26608 26794 26660 26800
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26344 25838 26372 26454
rect 26332 25832 26384 25838
rect 26332 25774 26384 25780
rect 26240 23588 26292 23594
rect 26240 23530 26292 23536
rect 25964 22568 26016 22574
rect 25964 22510 26016 22516
rect 23756 21616 23808 21622
rect 23756 21558 23808 21564
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23308 20058 23336 20198
rect 23296 20052 23348 20058
rect 23296 19994 23348 20000
rect 23216 19502 23336 19530
rect 23308 16454 23336 19502
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25412 17808 25464 17814
rect 25412 17750 25464 17756
rect 25424 17338 25452 17750
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25320 17128 25372 17134
rect 25320 17070 25372 17076
rect 25332 16522 25360 17070
rect 25424 16658 25452 17274
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25320 16516 25372 16522
rect 25320 16458 25372 16464
rect 23296 16448 23348 16454
rect 23296 16390 23348 16396
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 23216 14346 23244 15982
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 23308 10810 23336 16390
rect 24412 15570 24440 16390
rect 25700 16182 25728 19450
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25688 16176 25740 16182
rect 25688 16118 25740 16124
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 24400 15564 24452 15570
rect 24400 15506 24452 15512
rect 25424 15502 25452 15846
rect 25516 15502 25544 15982
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 23676 14550 23704 15438
rect 23664 14544 23716 14550
rect 23664 14486 23716 14492
rect 23572 14272 23624 14278
rect 23572 14214 23624 14220
rect 23584 13870 23612 14214
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23584 13734 23612 13806
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 25044 10532 25096 10538
rect 25044 10474 25096 10480
rect 25056 4078 25084 10474
rect 25596 8356 25648 8362
rect 25596 8298 25648 8304
rect 25608 8090 25636 8298
rect 25596 8084 25648 8090
rect 25596 8026 25648 8032
rect 25700 4298 25728 16118
rect 25792 7954 25820 18770
rect 25780 7948 25832 7954
rect 25780 7890 25832 7896
rect 25792 5166 25820 7890
rect 25780 5160 25832 5166
rect 25780 5102 25832 5108
rect 26252 4826 26280 23530
rect 26620 18970 26648 26794
rect 26712 26450 26740 29200
rect 26976 27532 27028 27538
rect 26804 27492 26976 27520
rect 26700 26444 26752 26450
rect 26700 26386 26752 26392
rect 26804 25838 26832 27492
rect 26976 27474 27028 27480
rect 27172 27062 27200 29200
rect 27252 27464 27304 27470
rect 27252 27406 27304 27412
rect 27160 27056 27212 27062
rect 27160 26998 27212 27004
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 26896 26246 26924 26862
rect 27264 26858 27292 27406
rect 27252 26852 27304 26858
rect 27252 26794 27304 26800
rect 27632 26518 27660 29200
rect 28552 27606 28580 29200
rect 28540 27600 28592 27606
rect 28540 27542 28592 27548
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28080 26920 28132 26926
rect 28080 26862 28132 26868
rect 27986 26616 28042 26625
rect 28092 26586 28120 26862
rect 28172 26852 28224 26858
rect 28172 26794 28224 26800
rect 28356 26852 28408 26858
rect 28356 26794 28408 26800
rect 27986 26551 27988 26560
rect 28040 26551 28042 26560
rect 28080 26580 28132 26586
rect 27988 26522 28040 26528
rect 28080 26522 28132 26528
rect 27620 26512 27672 26518
rect 27620 26454 27672 26460
rect 27804 26444 27856 26450
rect 27804 26386 27856 26392
rect 26884 26240 26936 26246
rect 26884 26182 26936 26188
rect 26792 25832 26844 25838
rect 26792 25774 26844 25780
rect 26608 18964 26660 18970
rect 26608 18906 26660 18912
rect 26804 18834 26832 25774
rect 26792 18828 26844 18834
rect 26792 18770 26844 18776
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26620 17134 26648 17614
rect 26608 17128 26660 17134
rect 26608 17070 26660 17076
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26516 16448 26568 16454
rect 26516 16390 26568 16396
rect 26528 8634 26556 16390
rect 26804 15978 26832 16594
rect 26896 16454 26924 26182
rect 27436 24268 27488 24274
rect 27436 24210 27488 24216
rect 27448 23526 27476 24210
rect 27436 23520 27488 23526
rect 27436 23462 27488 23468
rect 27448 23254 27476 23462
rect 27436 23248 27488 23254
rect 27436 23190 27488 23196
rect 27620 23248 27672 23254
rect 27620 23190 27672 23196
rect 27436 22432 27488 22438
rect 27436 22374 27488 22380
rect 27448 22098 27476 22374
rect 27252 22092 27304 22098
rect 27252 22034 27304 22040
rect 27436 22092 27488 22098
rect 27436 22034 27488 22040
rect 27264 21486 27292 22034
rect 27252 21480 27304 21486
rect 27252 21422 27304 21428
rect 27448 21010 27476 22034
rect 27632 21486 27660 23190
rect 27816 22234 27844 26386
rect 28184 26353 28212 26794
rect 28170 26344 28226 26353
rect 28170 26279 28226 26288
rect 28368 24138 28396 26794
rect 28448 24268 28500 24274
rect 28448 24210 28500 24216
rect 28356 24132 28408 24138
rect 28356 24074 28408 24080
rect 28460 23730 28488 24210
rect 28448 23724 28500 23730
rect 28448 23666 28500 23672
rect 28540 23656 28592 23662
rect 28540 23598 28592 23604
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 27804 22228 27856 22234
rect 27804 22170 27856 22176
rect 27620 21480 27672 21486
rect 27620 21422 27672 21428
rect 27436 21004 27488 21010
rect 27436 20946 27488 20952
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 27080 17882 27108 18770
rect 27632 17882 27660 21422
rect 28172 21412 28224 21418
rect 28172 21354 28224 21360
rect 28184 21146 28212 21354
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28184 21010 28212 21082
rect 28172 21004 28224 21010
rect 28172 20946 28224 20952
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27068 17876 27120 17882
rect 27068 17818 27120 17824
rect 27620 17876 27672 17882
rect 27620 17818 27672 17824
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26528 7954 26556 8570
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26528 7546 26556 7890
rect 26516 7540 26568 7546
rect 26516 7482 26568 7488
rect 26240 4820 26292 4826
rect 26240 4762 26292 4768
rect 25700 4282 25912 4298
rect 25700 4276 25924 4282
rect 25700 4270 25872 4276
rect 25700 4214 25728 4270
rect 25872 4218 25924 4224
rect 25688 4208 25740 4214
rect 25688 4150 25740 4156
rect 25700 4078 25728 4150
rect 25780 4140 25832 4146
rect 25780 4082 25832 4088
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 25688 4072 25740 4078
rect 25688 4014 25740 4020
rect 25136 3936 25188 3942
rect 25136 3878 25188 3884
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22652 3596 22704 3602
rect 22652 3538 22704 3544
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22008 3392 22060 3398
rect 22008 3334 22060 3340
rect 22020 2650 22048 3334
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22112 2854 22140 2926
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22008 2644 22060 2650
rect 22008 2586 22060 2592
rect 21916 2576 21968 2582
rect 21836 2536 21916 2564
rect 21916 2518 21968 2524
rect 21640 2372 21692 2378
rect 21640 2314 21692 2320
rect 21364 2304 21416 2310
rect 21364 2246 21416 2252
rect 21376 1902 21404 2246
rect 21364 1896 21416 1902
rect 21364 1838 21416 1844
rect 21652 800 21680 2314
rect 22020 1902 22048 2586
rect 22008 1896 22060 1902
rect 22008 1838 22060 1844
rect 22112 800 22140 2790
rect 22204 2446 22232 3470
rect 22560 2848 22612 2854
rect 22560 2790 22612 2796
rect 22572 2514 22600 2790
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 22192 2440 22244 2446
rect 22664 2394 22692 3538
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24320 2990 24348 3334
rect 25148 2990 25176 3878
rect 25792 3738 25820 4082
rect 25872 4072 25924 4078
rect 25872 4014 25924 4020
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 24308 2984 24360 2990
rect 24308 2926 24360 2932
rect 25136 2984 25188 2990
rect 25136 2926 25188 2932
rect 23480 2644 23532 2650
rect 23480 2586 23532 2592
rect 22192 2382 22244 2388
rect 22572 2366 22692 2394
rect 22572 800 22600 2366
rect 23492 800 23520 2586
rect 23940 2372 23992 2378
rect 23940 2314 23992 2320
rect 23952 800 23980 2314
rect 24320 2038 24348 2926
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 25320 2916 25372 2922
rect 25320 2858 25372 2864
rect 25780 2916 25832 2922
rect 25780 2858 25832 2864
rect 24308 2032 24360 2038
rect 24308 1974 24360 1980
rect 24872 800 24900 2858
rect 25332 800 25360 2858
rect 25792 800 25820 2858
rect 25884 2854 25912 4014
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25976 2990 26004 3878
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 25964 2984 26016 2990
rect 25964 2926 26016 2932
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 25884 2514 25912 2790
rect 25872 2508 25924 2514
rect 25872 2450 25924 2456
rect 26160 2446 26188 3538
rect 26252 2990 26280 4762
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27252 4480 27304 4486
rect 27252 4422 27304 4428
rect 26976 4208 27028 4214
rect 26976 4150 27028 4156
rect 26332 3460 26384 3466
rect 26332 3402 26384 3408
rect 26240 2984 26292 2990
rect 26240 2926 26292 2932
rect 26344 2514 26372 3402
rect 26988 2990 27016 4150
rect 27264 4146 27292 4422
rect 27252 4140 27304 4146
rect 27252 4082 27304 4088
rect 27160 3460 27212 3466
rect 27160 3402 27212 3408
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 26792 2848 26844 2854
rect 26712 2808 26792 2836
rect 26332 2508 26384 2514
rect 26332 2450 26384 2456
rect 26056 2440 26108 2446
rect 26056 2382 26108 2388
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26068 1834 26096 2382
rect 26056 1828 26108 1834
rect 26056 1770 26108 1776
rect 26712 800 26740 2808
rect 26792 2790 26844 2796
rect 27172 800 27200 3402
rect 27448 2582 27476 4626
rect 27724 4554 27752 20878
rect 27896 18828 27948 18834
rect 27896 18770 27948 18776
rect 27908 8022 27936 18770
rect 27896 8016 27948 8022
rect 27896 7958 27948 7964
rect 27908 7546 27936 7958
rect 27896 7540 27948 7546
rect 27896 7482 27948 7488
rect 27712 4548 27764 4554
rect 27712 4490 27764 4496
rect 27620 3936 27672 3942
rect 27620 3878 27672 3884
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 27632 3534 27660 3878
rect 28092 3602 28120 3878
rect 27804 3596 27856 3602
rect 27804 3538 27856 3544
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 27620 3528 27672 3534
rect 27620 3470 27672 3476
rect 27632 3058 27660 3470
rect 27816 3194 27844 3538
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 27620 3052 27672 3058
rect 27620 2994 27672 3000
rect 27436 2576 27488 2582
rect 27436 2518 27488 2524
rect 28092 800 28120 3538
rect 28276 2378 28304 23462
rect 28552 23322 28580 23598
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28552 21078 28580 23258
rect 28540 21072 28592 21078
rect 28540 21014 28592 21020
rect 28736 17746 28764 27270
rect 29012 27062 29040 29200
rect 29736 28008 29788 28014
rect 29736 27950 29788 27956
rect 29748 27606 29776 27950
rect 29932 27674 29960 29200
rect 30196 27940 30248 27946
rect 30196 27882 30248 27888
rect 29920 27668 29972 27674
rect 29920 27610 29972 27616
rect 29736 27600 29788 27606
rect 29736 27542 29788 27548
rect 29368 27532 29420 27538
rect 29368 27474 29420 27480
rect 29184 27328 29236 27334
rect 29184 27270 29236 27276
rect 29000 27056 29052 27062
rect 29000 26998 29052 27004
rect 28908 24608 28960 24614
rect 28908 24550 28960 24556
rect 28920 24274 28948 24550
rect 28908 24268 28960 24274
rect 28908 24210 28960 24216
rect 28724 17740 28776 17746
rect 28724 17682 28776 17688
rect 29196 16182 29224 27270
rect 29276 21344 29328 21350
rect 29276 21286 29328 21292
rect 29288 21078 29316 21286
rect 29276 21072 29328 21078
rect 29276 21014 29328 21020
rect 29380 20622 29408 27474
rect 29852 27228 30148 27248
rect 29908 27226 29932 27228
rect 29988 27226 30012 27228
rect 30068 27226 30092 27228
rect 29930 27174 29932 27226
rect 29994 27174 30006 27226
rect 30068 27174 30070 27226
rect 29908 27172 29932 27174
rect 29988 27172 30012 27174
rect 30068 27172 30092 27174
rect 29852 27152 30148 27172
rect 30208 27130 30236 27882
rect 30288 27396 30340 27402
rect 30288 27338 30340 27344
rect 30300 27130 30328 27338
rect 30196 27124 30248 27130
rect 30196 27066 30248 27072
rect 30288 27124 30340 27130
rect 30288 27066 30340 27072
rect 29552 27056 29604 27062
rect 29552 26998 29604 27004
rect 29460 26988 29512 26994
rect 29460 26930 29512 26936
rect 29472 25838 29500 26930
rect 29564 26489 29592 26998
rect 29550 26480 29606 26489
rect 30392 26450 30420 29200
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 30484 26994 30512 27270
rect 30852 27062 30880 29200
rect 31484 27668 31536 27674
rect 31484 27610 31536 27616
rect 31496 27470 31524 27610
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31208 27328 31260 27334
rect 31208 27270 31260 27276
rect 30840 27056 30892 27062
rect 30840 26998 30892 27004
rect 30472 26988 30524 26994
rect 30472 26930 30524 26936
rect 29550 26415 29606 26424
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 29852 26140 30148 26160
rect 29908 26138 29932 26140
rect 29988 26138 30012 26140
rect 30068 26138 30092 26140
rect 29930 26086 29932 26138
rect 29994 26086 30006 26138
rect 30068 26086 30070 26138
rect 29908 26084 29932 26086
rect 29988 26084 30012 26086
rect 30068 26084 30092 26086
rect 29852 26064 30148 26084
rect 29460 25832 29512 25838
rect 29460 25774 29512 25780
rect 29472 21690 29500 25774
rect 29852 25052 30148 25072
rect 29908 25050 29932 25052
rect 29988 25050 30012 25052
rect 30068 25050 30092 25052
rect 29930 24998 29932 25050
rect 29994 24998 30006 25050
rect 30068 24998 30070 25050
rect 29908 24996 29932 24998
rect 29988 24996 30012 24998
rect 30068 24996 30092 24998
rect 29852 24976 30148 24996
rect 29644 24880 29696 24886
rect 29644 24822 29696 24828
rect 29460 21684 29512 21690
rect 29460 21626 29512 21632
rect 29472 21486 29500 21626
rect 29460 21480 29512 21486
rect 29460 21422 29512 21428
rect 29288 20594 29408 20622
rect 29472 20622 29500 21422
rect 29472 20594 29592 20622
rect 29288 16522 29316 20594
rect 29460 16720 29512 16726
rect 29460 16662 29512 16668
rect 29368 16652 29420 16658
rect 29368 16594 29420 16600
rect 29276 16516 29328 16522
rect 29276 16458 29328 16464
rect 29380 16266 29408 16594
rect 29288 16238 29408 16266
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29288 16046 29316 16238
rect 29092 16040 29144 16046
rect 29092 15982 29144 15988
rect 29276 16040 29328 16046
rect 29276 15982 29328 15988
rect 29104 15910 29132 15982
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 29092 15904 29144 15910
rect 29092 15846 29144 15852
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 28264 2372 28316 2378
rect 28264 2314 28316 2320
rect 28368 1698 28396 15506
rect 28540 11008 28592 11014
rect 28540 10950 28592 10956
rect 28552 2582 28580 10950
rect 28724 4616 28776 4622
rect 28724 4558 28776 4564
rect 28736 3602 28764 4558
rect 28816 4480 28868 4486
rect 28816 4422 28868 4428
rect 28828 4214 28856 4422
rect 28920 4282 28948 15846
rect 29288 15706 29316 15982
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 29472 4282 29500 16662
rect 29564 16454 29592 20594
rect 29552 16448 29604 16454
rect 29552 16390 29604 16396
rect 29564 16046 29592 16390
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 28908 4276 28960 4282
rect 28908 4218 28960 4224
rect 29460 4276 29512 4282
rect 29460 4218 29512 4224
rect 28816 4208 28868 4214
rect 28816 4150 28868 4156
rect 28724 3596 28776 3602
rect 28724 3538 28776 3544
rect 28632 3392 28684 3398
rect 28632 3334 28684 3340
rect 28540 2576 28592 2582
rect 28540 2518 28592 2524
rect 28644 1714 28672 3334
rect 28828 2990 28856 4150
rect 28920 2990 28948 4218
rect 29368 3188 29420 3194
rect 29368 3130 29420 3136
rect 28816 2984 28868 2990
rect 28816 2926 28868 2932
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 29380 2650 29408 3130
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 29472 2514 29500 4218
rect 29656 3058 29684 24822
rect 29852 23964 30148 23984
rect 29908 23962 29932 23964
rect 29988 23962 30012 23964
rect 30068 23962 30092 23964
rect 29930 23910 29932 23962
rect 29994 23910 30006 23962
rect 30068 23910 30070 23962
rect 29908 23908 29932 23910
rect 29988 23908 30012 23910
rect 30068 23908 30092 23910
rect 29852 23888 30148 23908
rect 29852 22876 30148 22896
rect 29908 22874 29932 22876
rect 29988 22874 30012 22876
rect 30068 22874 30092 22876
rect 29930 22822 29932 22874
rect 29994 22822 30006 22874
rect 30068 22822 30070 22874
rect 29908 22820 29932 22822
rect 29988 22820 30012 22822
rect 30068 22820 30092 22822
rect 29852 22800 30148 22820
rect 29852 21788 30148 21808
rect 29908 21786 29932 21788
rect 29988 21786 30012 21788
rect 30068 21786 30092 21788
rect 29930 21734 29932 21786
rect 29994 21734 30006 21786
rect 30068 21734 30070 21786
rect 29908 21732 29932 21734
rect 29988 21732 30012 21734
rect 30068 21732 30092 21734
rect 29852 21712 30148 21732
rect 29852 20700 30148 20720
rect 29908 20698 29932 20700
rect 29988 20698 30012 20700
rect 30068 20698 30092 20700
rect 29930 20646 29932 20698
rect 29994 20646 30006 20698
rect 30068 20646 30070 20698
rect 29908 20644 29932 20646
rect 29988 20644 30012 20646
rect 30068 20644 30092 20646
rect 29852 20624 30148 20644
rect 29852 19612 30148 19632
rect 29908 19610 29932 19612
rect 29988 19610 30012 19612
rect 30068 19610 30092 19612
rect 29930 19558 29932 19610
rect 29994 19558 30006 19610
rect 30068 19558 30070 19610
rect 29908 19556 29932 19558
rect 29988 19556 30012 19558
rect 30068 19556 30092 19558
rect 29852 19536 30148 19556
rect 29852 18524 30148 18544
rect 29908 18522 29932 18524
rect 29988 18522 30012 18524
rect 30068 18522 30092 18524
rect 29930 18470 29932 18522
rect 29994 18470 30006 18522
rect 30068 18470 30070 18522
rect 29908 18468 29932 18470
rect 29988 18468 30012 18470
rect 30068 18468 30092 18470
rect 29852 18448 30148 18468
rect 29852 17436 30148 17456
rect 29908 17434 29932 17436
rect 29988 17434 30012 17436
rect 30068 17434 30092 17436
rect 29930 17382 29932 17434
rect 29994 17382 30006 17434
rect 30068 17382 30070 17434
rect 29908 17380 29932 17382
rect 29988 17380 30012 17382
rect 30068 17380 30092 17382
rect 29852 17360 30148 17380
rect 29852 16348 30148 16368
rect 29908 16346 29932 16348
rect 29988 16346 30012 16348
rect 30068 16346 30092 16348
rect 29930 16294 29932 16346
rect 29994 16294 30006 16346
rect 30068 16294 30070 16346
rect 29908 16292 29932 16294
rect 29988 16292 30012 16294
rect 30068 16292 30092 16294
rect 29852 16272 30148 16292
rect 29736 16244 29788 16250
rect 29736 16186 29788 16192
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 29748 15910 29776 16186
rect 30208 15978 30236 16186
rect 30196 15972 30248 15978
rect 30196 15914 30248 15920
rect 29736 15904 29788 15910
rect 29736 15846 29788 15852
rect 29852 15260 30148 15280
rect 29908 15258 29932 15260
rect 29988 15258 30012 15260
rect 30068 15258 30092 15260
rect 29930 15206 29932 15258
rect 29994 15206 30006 15258
rect 30068 15206 30070 15258
rect 29908 15204 29932 15206
rect 29988 15204 30012 15206
rect 30068 15204 30092 15206
rect 29852 15184 30148 15204
rect 29852 14172 30148 14192
rect 29908 14170 29932 14172
rect 29988 14170 30012 14172
rect 30068 14170 30092 14172
rect 29930 14118 29932 14170
rect 29994 14118 30006 14170
rect 30068 14118 30070 14170
rect 29908 14116 29932 14118
rect 29988 14116 30012 14118
rect 30068 14116 30092 14118
rect 29852 14096 30148 14116
rect 29852 13084 30148 13104
rect 29908 13082 29932 13084
rect 29988 13082 30012 13084
rect 30068 13082 30092 13084
rect 29930 13030 29932 13082
rect 29994 13030 30006 13082
rect 30068 13030 30070 13082
rect 29908 13028 29932 13030
rect 29988 13028 30012 13030
rect 30068 13028 30092 13030
rect 29852 13008 30148 13028
rect 29852 11996 30148 12016
rect 29908 11994 29932 11996
rect 29988 11994 30012 11996
rect 30068 11994 30092 11996
rect 29930 11942 29932 11994
rect 29994 11942 30006 11994
rect 30068 11942 30070 11994
rect 29908 11940 29932 11942
rect 29988 11940 30012 11942
rect 30068 11940 30092 11942
rect 29852 11920 30148 11940
rect 29852 10908 30148 10928
rect 29908 10906 29932 10908
rect 29988 10906 30012 10908
rect 30068 10906 30092 10908
rect 29930 10854 29932 10906
rect 29994 10854 30006 10906
rect 30068 10854 30070 10906
rect 29908 10852 29932 10854
rect 29988 10852 30012 10854
rect 30068 10852 30092 10854
rect 29852 10832 30148 10852
rect 29852 9820 30148 9840
rect 29908 9818 29932 9820
rect 29988 9818 30012 9820
rect 30068 9818 30092 9820
rect 29930 9766 29932 9818
rect 29994 9766 30006 9818
rect 30068 9766 30070 9818
rect 29908 9764 29932 9766
rect 29988 9764 30012 9766
rect 30068 9764 30092 9766
rect 29852 9744 30148 9764
rect 29852 8732 30148 8752
rect 29908 8730 29932 8732
rect 29988 8730 30012 8732
rect 30068 8730 30092 8732
rect 29930 8678 29932 8730
rect 29994 8678 30006 8730
rect 30068 8678 30070 8730
rect 29908 8676 29932 8678
rect 29988 8676 30012 8678
rect 30068 8676 30092 8678
rect 29852 8656 30148 8676
rect 29852 7644 30148 7664
rect 29908 7642 29932 7644
rect 29988 7642 30012 7644
rect 30068 7642 30092 7644
rect 29930 7590 29932 7642
rect 29994 7590 30006 7642
rect 30068 7590 30070 7642
rect 29908 7588 29932 7590
rect 29988 7588 30012 7590
rect 30068 7588 30092 7590
rect 29852 7568 30148 7588
rect 29852 6556 30148 6576
rect 29908 6554 29932 6556
rect 29988 6554 30012 6556
rect 30068 6554 30092 6556
rect 29930 6502 29932 6554
rect 29994 6502 30006 6554
rect 30068 6502 30070 6554
rect 29908 6500 29932 6502
rect 29988 6500 30012 6502
rect 30068 6500 30092 6502
rect 29852 6480 30148 6500
rect 29852 5468 30148 5488
rect 29908 5466 29932 5468
rect 29988 5466 30012 5468
rect 30068 5466 30092 5468
rect 29930 5414 29932 5466
rect 29994 5414 30006 5466
rect 30068 5414 30070 5466
rect 29908 5412 29932 5414
rect 29988 5412 30012 5414
rect 30068 5412 30092 5414
rect 29852 5392 30148 5412
rect 29852 4380 30148 4400
rect 29908 4378 29932 4380
rect 29988 4378 30012 4380
rect 30068 4378 30092 4380
rect 29930 4326 29932 4378
rect 29994 4326 30006 4378
rect 30068 4326 30070 4378
rect 29908 4324 29932 4326
rect 29988 4324 30012 4326
rect 30068 4324 30092 4326
rect 29852 4304 30148 4324
rect 30484 3738 30512 26930
rect 31024 26852 31076 26858
rect 31024 26794 31076 26800
rect 30932 26784 30984 26790
rect 30932 26726 30984 26732
rect 30944 25770 30972 26726
rect 30932 25764 30984 25770
rect 30932 25706 30984 25712
rect 31036 21690 31064 26794
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 31116 20936 31168 20942
rect 31116 20878 31168 20884
rect 31128 19922 31156 20878
rect 31116 19916 31168 19922
rect 31116 19858 31168 19864
rect 30932 10600 30984 10606
rect 30932 10542 30984 10548
rect 30944 9654 30972 10542
rect 30932 9648 30984 9654
rect 30932 9590 30984 9596
rect 31220 3738 31248 27270
rect 31772 26926 31800 29200
rect 32232 27606 32260 29200
rect 32220 27600 32272 27606
rect 32220 27542 32272 27548
rect 31760 26920 31812 26926
rect 31760 26862 31812 26868
rect 31772 26586 31800 26862
rect 32588 26852 32640 26858
rect 32588 26794 32640 26800
rect 31760 26580 31812 26586
rect 31760 26522 31812 26528
rect 32600 26246 32628 26794
rect 33152 26518 33180 29200
rect 33612 27538 33640 29200
rect 33968 28008 34020 28014
rect 33968 27950 34020 27956
rect 33980 27606 34008 27950
rect 33968 27600 34020 27606
rect 33968 27542 34020 27548
rect 33600 27532 33652 27538
rect 33600 27474 33652 27480
rect 33508 27464 33560 27470
rect 33508 27406 33560 27412
rect 33416 26988 33468 26994
rect 33416 26930 33468 26936
rect 33324 26784 33376 26790
rect 33324 26726 33376 26732
rect 33336 26518 33364 26726
rect 33140 26512 33192 26518
rect 33140 26454 33192 26460
rect 33324 26512 33376 26518
rect 33324 26454 33376 26460
rect 32588 26240 32640 26246
rect 32588 26182 32640 26188
rect 32312 25968 32364 25974
rect 32312 25910 32364 25916
rect 32324 24750 32352 25910
rect 32600 25498 32628 26182
rect 33324 25832 33376 25838
rect 33428 25820 33456 26930
rect 33520 26790 33548 27406
rect 33876 26920 33928 26926
rect 33876 26862 33928 26868
rect 33508 26784 33560 26790
rect 33508 26726 33560 26732
rect 33376 25792 33456 25820
rect 33324 25774 33376 25780
rect 32588 25492 32640 25498
rect 32588 25434 32640 25440
rect 32312 24744 32364 24750
rect 32312 24686 32364 24692
rect 31392 21480 31444 21486
rect 31392 21422 31444 21428
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 31312 20398 31340 21354
rect 31300 20392 31352 20398
rect 31300 20334 31352 20340
rect 31404 19922 31432 21422
rect 32220 21004 32272 21010
rect 32220 20946 32272 20952
rect 32232 20398 32260 20946
rect 32220 20392 32272 20398
rect 32220 20334 32272 20340
rect 32680 20392 32732 20398
rect 32680 20334 32732 20340
rect 31944 20324 31996 20330
rect 31944 20266 31996 20272
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 31484 19780 31536 19786
rect 31484 19722 31536 19728
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 31208 3732 31260 3738
rect 31208 3674 31260 3680
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 29736 3392 29788 3398
rect 29736 3334 29788 3340
rect 29644 3052 29696 3058
rect 29644 2994 29696 3000
rect 29748 2990 29776 3334
rect 29852 3292 30148 3312
rect 29908 3290 29932 3292
rect 29988 3290 30012 3292
rect 30068 3290 30092 3292
rect 29930 3238 29932 3290
rect 29994 3238 30006 3290
rect 30068 3238 30070 3290
rect 29908 3236 29932 3238
rect 29988 3236 30012 3238
rect 30068 3236 30092 3238
rect 29852 3216 30148 3236
rect 29736 2984 29788 2990
rect 29736 2926 29788 2932
rect 29748 2514 29776 2926
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 29460 2508 29512 2514
rect 29460 2450 29512 2456
rect 29736 2508 29788 2514
rect 29736 2450 29788 2456
rect 28356 1692 28408 1698
rect 28356 1634 28408 1640
rect 28552 1686 28672 1714
rect 28552 800 28580 1686
rect 29012 800 29040 2450
rect 29852 2204 30148 2224
rect 29908 2202 29932 2204
rect 29988 2202 30012 2204
rect 30068 2202 30092 2204
rect 29930 2150 29932 2202
rect 29994 2150 30006 2202
rect 30068 2150 30070 2202
rect 29908 2148 29932 2150
rect 29988 2148 30012 2150
rect 30068 2148 30092 2150
rect 29852 2128 30148 2148
rect 30208 2020 30236 3538
rect 31220 2990 31248 3674
rect 31208 2984 31260 2990
rect 31208 2926 31260 2932
rect 30380 2916 30432 2922
rect 30380 2858 30432 2864
rect 29932 1992 30236 2020
rect 29932 800 29960 1992
rect 30392 800 30420 2858
rect 31496 2582 31524 19722
rect 31956 2990 31984 20266
rect 32692 19990 32720 20334
rect 32680 19984 32732 19990
rect 32680 19926 32732 19932
rect 32220 19916 32272 19922
rect 32220 19858 32272 19864
rect 32404 19916 32456 19922
rect 32404 19858 32456 19864
rect 32232 19174 32260 19858
rect 32220 19168 32272 19174
rect 32220 19110 32272 19116
rect 32416 3738 32444 19858
rect 33232 15496 33284 15502
rect 33232 15438 33284 15444
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 31760 2916 31812 2922
rect 31760 2858 31812 2864
rect 31484 2576 31536 2582
rect 31484 2518 31536 2524
rect 31300 2372 31352 2378
rect 31300 2314 31352 2320
rect 31312 800 31340 2314
rect 31772 800 31800 2858
rect 32232 800 32260 3538
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 33152 800 33180 2586
rect 33244 2514 33272 15438
rect 33336 9926 33364 25774
rect 33520 25770 33548 26726
rect 33888 26042 33916 26862
rect 34072 26450 34100 29200
rect 34336 28076 34388 28082
rect 34336 28018 34388 28024
rect 34152 27600 34204 27606
rect 34152 27542 34204 27548
rect 34164 26586 34192 27542
rect 34152 26580 34204 26586
rect 34152 26522 34204 26528
rect 34348 26450 34376 28018
rect 34612 27940 34664 27946
rect 34612 27882 34664 27888
rect 34428 27532 34480 27538
rect 34428 27474 34480 27480
rect 34060 26444 34112 26450
rect 34060 26386 34112 26392
rect 34336 26444 34388 26450
rect 34336 26386 34388 26392
rect 34072 26042 34100 26386
rect 33876 26036 33928 26042
rect 33876 25978 33928 25984
rect 34060 26036 34112 26042
rect 34060 25978 34112 25984
rect 33508 25764 33560 25770
rect 33508 25706 33560 25712
rect 33520 25294 33548 25706
rect 33888 25498 33916 25978
rect 33876 25492 33928 25498
rect 33876 25434 33928 25440
rect 33508 25288 33560 25294
rect 33508 25230 33560 25236
rect 34348 24954 34376 26386
rect 34440 26042 34468 27474
rect 34520 26784 34572 26790
rect 34520 26726 34572 26732
rect 34532 26489 34560 26726
rect 34518 26480 34574 26489
rect 34518 26415 34574 26424
rect 34428 26036 34480 26042
rect 34428 25978 34480 25984
rect 34336 24948 34388 24954
rect 34336 24890 34388 24896
rect 34624 22778 34652 27882
rect 34888 27328 34940 27334
rect 34888 27270 34940 27276
rect 34704 26920 34756 26926
rect 34704 26862 34756 26868
rect 34716 26246 34744 26862
rect 34704 26240 34756 26246
rect 34704 26182 34756 26188
rect 34612 22772 34664 22778
rect 34612 22714 34664 22720
rect 34716 13870 34744 26182
rect 34900 18698 34928 27270
rect 34992 25838 35020 29200
rect 35452 27606 35480 29200
rect 35440 27600 35492 27606
rect 35440 27542 35492 27548
rect 35808 26920 35860 26926
rect 35808 26862 35860 26868
rect 35714 26616 35770 26625
rect 35820 26586 35848 26862
rect 36268 26852 36320 26858
rect 36268 26794 36320 26800
rect 36176 26784 36228 26790
rect 36176 26726 36228 26732
rect 35714 26551 35770 26560
rect 35808 26580 35860 26586
rect 35728 26450 35756 26551
rect 35808 26522 35860 26528
rect 35716 26444 35768 26450
rect 35716 26386 35768 26392
rect 34980 25832 35032 25838
rect 34980 25774 35032 25780
rect 35728 25498 35756 26386
rect 35716 25492 35768 25498
rect 35716 25434 35768 25440
rect 36188 25226 36216 26726
rect 36280 26586 36308 26794
rect 36268 26580 36320 26586
rect 36268 26522 36320 26528
rect 36372 26450 36400 29200
rect 36636 27532 36688 27538
rect 36636 27474 36688 27480
rect 36360 26444 36412 26450
rect 36360 26386 36412 26392
rect 36372 26042 36400 26386
rect 36360 26036 36412 26042
rect 36360 25978 36412 25984
rect 36176 25220 36228 25226
rect 36176 25162 36228 25168
rect 36452 25152 36504 25158
rect 36452 25094 36504 25100
rect 35900 23588 35952 23594
rect 35900 23530 35952 23536
rect 35912 21486 35940 23530
rect 35992 22568 36044 22574
rect 35992 22510 36044 22516
rect 35900 21480 35952 21486
rect 35900 21422 35952 21428
rect 36004 21010 36032 22510
rect 36268 22092 36320 22098
rect 36268 22034 36320 22040
rect 36084 21344 36136 21350
rect 36084 21286 36136 21292
rect 36096 21078 36124 21286
rect 36084 21072 36136 21078
rect 36084 21014 36136 21020
rect 35992 21004 36044 21010
rect 35992 20946 36044 20952
rect 36084 20936 36136 20942
rect 36084 20878 36136 20884
rect 35808 19916 35860 19922
rect 35808 19858 35860 19864
rect 35820 19718 35848 19858
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35820 19446 35848 19654
rect 35808 19440 35860 19446
rect 35808 19382 35860 19388
rect 34888 18692 34940 18698
rect 34888 18634 34940 18640
rect 35992 16040 36044 16046
rect 35992 15982 36044 15988
rect 35900 15904 35952 15910
rect 35900 15846 35952 15852
rect 35912 15638 35940 15846
rect 36004 15706 36032 15982
rect 35992 15700 36044 15706
rect 35992 15642 36044 15648
rect 35900 15632 35952 15638
rect 35900 15574 35952 15580
rect 35440 14884 35492 14890
rect 35440 14826 35492 14832
rect 34704 13864 34756 13870
rect 34704 13806 34756 13812
rect 34612 13728 34664 13734
rect 34612 13670 34664 13676
rect 33324 9920 33376 9926
rect 33324 9862 33376 9868
rect 33968 5840 34020 5846
rect 33968 5782 34020 5788
rect 33980 5370 34008 5782
rect 33968 5364 34020 5370
rect 33968 5306 34020 5312
rect 33980 5030 34008 5306
rect 33968 5024 34020 5030
rect 33968 4966 34020 4972
rect 34624 4078 34652 13670
rect 35348 9512 35400 9518
rect 35348 9454 35400 9460
rect 34796 5228 34848 5234
rect 34796 5170 34848 5176
rect 34612 4072 34664 4078
rect 34612 4014 34664 4020
rect 34060 3596 34112 3602
rect 34060 3538 34112 3544
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33232 2508 33284 2514
rect 33232 2450 33284 2456
rect 33612 800 33640 2926
rect 33784 2848 33836 2854
rect 33784 2790 33836 2796
rect 33796 1698 33824 2790
rect 33784 1692 33836 1698
rect 33784 1634 33836 1640
rect 34072 800 34100 3538
rect 34624 3482 34652 4014
rect 34808 3738 34836 5170
rect 34980 3936 35032 3942
rect 34980 3878 35032 3884
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 34992 3602 35020 3878
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 34624 3454 34744 3482
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34624 2990 34652 3334
rect 34612 2984 34664 2990
rect 34612 2926 34664 2932
rect 34716 2922 34744 3454
rect 34704 2916 34756 2922
rect 34704 2858 34756 2864
rect 34992 800 35020 3538
rect 35072 3120 35124 3126
rect 35072 3062 35124 3068
rect 35084 2650 35112 3062
rect 35360 3058 35388 9454
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 35072 2644 35124 2650
rect 35072 2586 35124 2592
rect 35452 2496 35480 14826
rect 36096 5370 36124 20878
rect 36280 20874 36308 22034
rect 36268 20868 36320 20874
rect 36268 20810 36320 20816
rect 36360 20256 36412 20262
rect 36360 20198 36412 20204
rect 36268 17672 36320 17678
rect 36268 17614 36320 17620
rect 36280 17134 36308 17614
rect 36268 17128 36320 17134
rect 36268 17070 36320 17076
rect 36280 16046 36308 17070
rect 36268 16040 36320 16046
rect 36268 15982 36320 15988
rect 36176 12232 36228 12238
rect 36176 12174 36228 12180
rect 36084 5364 36136 5370
rect 36084 5306 36136 5312
rect 35624 5024 35676 5030
rect 35624 4966 35676 4972
rect 35636 4826 35664 4966
rect 35624 4820 35676 4826
rect 35624 4762 35676 4768
rect 36084 4004 36136 4010
rect 36084 3946 36136 3952
rect 36096 2514 36124 3946
rect 36188 3058 36216 12174
rect 36372 4486 36400 20198
rect 36464 17066 36492 25094
rect 36648 24970 36676 27474
rect 36832 27402 36860 29200
rect 37292 27606 37320 29200
rect 37464 28144 37516 28150
rect 37464 28086 37516 28092
rect 37280 27600 37332 27606
rect 37280 27542 37332 27548
rect 36820 27396 36872 27402
rect 36820 27338 36872 27344
rect 36728 26920 36780 26926
rect 36728 26862 36780 26868
rect 36740 25158 36768 26862
rect 37476 26450 37504 28086
rect 37832 27668 37884 27674
rect 37832 27610 37884 27616
rect 37556 27600 37608 27606
rect 37556 27542 37608 27548
rect 37280 26444 37332 26450
rect 37280 26386 37332 26392
rect 37464 26444 37516 26450
rect 37464 26386 37516 26392
rect 36820 25832 36872 25838
rect 36820 25774 36872 25780
rect 36728 25152 36780 25158
rect 36728 25094 36780 25100
rect 36648 24942 36768 24970
rect 36740 24614 36768 24942
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 36740 23526 36768 24550
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36544 22568 36596 22574
rect 36544 22510 36596 22516
rect 36556 21962 36584 22510
rect 36544 21956 36596 21962
rect 36544 21898 36596 21904
rect 36556 21418 36584 21898
rect 36544 21412 36596 21418
rect 36544 21354 36596 21360
rect 36556 20398 36584 21354
rect 36636 20936 36688 20942
rect 36636 20878 36688 20884
rect 36544 20392 36596 20398
rect 36544 20334 36596 20340
rect 36556 19922 36584 20334
rect 36544 19916 36596 19922
rect 36544 19858 36596 19864
rect 36452 17060 36504 17066
rect 36452 17002 36504 17008
rect 36360 4480 36412 4486
rect 36360 4422 36412 4428
rect 36648 3602 36676 20878
rect 36832 14958 36860 25774
rect 37292 24614 37320 26386
rect 37476 25498 37504 26386
rect 37568 25838 37596 27542
rect 37648 26308 37700 26314
rect 37648 26250 37700 26256
rect 37660 25906 37688 26250
rect 37844 26042 37872 27610
rect 38016 27600 38068 27606
rect 38016 27542 38068 27548
rect 37832 26036 37884 26042
rect 37832 25978 37884 25984
rect 37648 25900 37700 25906
rect 37648 25842 37700 25848
rect 37556 25832 37608 25838
rect 37556 25774 37608 25780
rect 37740 25832 37792 25838
rect 37740 25774 37792 25780
rect 37464 25492 37516 25498
rect 37516 25452 37596 25480
rect 37464 25434 37516 25440
rect 37464 25220 37516 25226
rect 37464 25162 37516 25168
rect 37280 24608 37332 24614
rect 37280 24550 37332 24556
rect 37096 20936 37148 20942
rect 37096 20878 37148 20884
rect 37108 20398 37136 20878
rect 37096 20392 37148 20398
rect 37096 20334 37148 20340
rect 37096 16652 37148 16658
rect 37096 16594 37148 16600
rect 37108 16250 37136 16594
rect 37096 16244 37148 16250
rect 37096 16186 37148 16192
rect 37096 15972 37148 15978
rect 37096 15914 37148 15920
rect 37108 15706 37136 15914
rect 37096 15700 37148 15706
rect 37096 15642 37148 15648
rect 37292 15502 37320 24550
rect 37476 16590 37504 25162
rect 37568 24410 37596 25452
rect 37752 25362 37780 25774
rect 38028 25770 38056 27542
rect 38212 26450 38240 29200
rect 38476 27328 38528 27334
rect 38476 27270 38528 27276
rect 38200 26444 38252 26450
rect 38200 26386 38252 26392
rect 38488 26042 38516 27270
rect 38672 26926 38700 29200
rect 39592 27962 39620 29200
rect 39592 27934 39896 27962
rect 39484 27772 39780 27792
rect 39540 27770 39564 27772
rect 39620 27770 39644 27772
rect 39700 27770 39724 27772
rect 39562 27718 39564 27770
rect 39626 27718 39638 27770
rect 39700 27718 39702 27770
rect 39540 27716 39564 27718
rect 39620 27716 39644 27718
rect 39700 27716 39724 27718
rect 39484 27696 39780 27716
rect 39304 27532 39356 27538
rect 39304 27474 39356 27480
rect 39026 27432 39082 27441
rect 39026 27367 39028 27376
rect 39080 27367 39082 27376
rect 39028 27338 39080 27344
rect 39120 27328 39172 27334
rect 39120 27270 39172 27276
rect 38660 26920 38712 26926
rect 38660 26862 38712 26868
rect 38752 26512 38804 26518
rect 38752 26454 38804 26460
rect 38568 26444 38620 26450
rect 38568 26386 38620 26392
rect 38580 26042 38608 26386
rect 38660 26376 38712 26382
rect 38660 26318 38712 26324
rect 38476 26036 38528 26042
rect 38476 25978 38528 25984
rect 38568 26036 38620 26042
rect 38568 25978 38620 25984
rect 38016 25764 38068 25770
rect 38016 25706 38068 25712
rect 37740 25356 37792 25362
rect 37740 25298 37792 25304
rect 37556 24404 37608 24410
rect 37556 24346 37608 24352
rect 37752 24274 37780 25298
rect 37924 25288 37976 25294
rect 37924 25230 37976 25236
rect 37740 24268 37792 24274
rect 37740 24210 37792 24216
rect 37752 23798 37780 24210
rect 37740 23792 37792 23798
rect 37740 23734 37792 23740
rect 37832 21480 37884 21486
rect 37832 21422 37884 21428
rect 37844 21010 37872 21422
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 37936 20622 37964 25230
rect 38028 24886 38056 25706
rect 38488 24886 38516 25978
rect 38672 25838 38700 26318
rect 38660 25832 38712 25838
rect 38660 25774 38712 25780
rect 38568 25764 38620 25770
rect 38568 25706 38620 25712
rect 38580 25362 38608 25706
rect 38764 25498 38792 26454
rect 38844 26240 38896 26246
rect 38844 26182 38896 26188
rect 38752 25492 38804 25498
rect 38752 25434 38804 25440
rect 38568 25356 38620 25362
rect 38568 25298 38620 25304
rect 38016 24880 38068 24886
rect 38016 24822 38068 24828
rect 38476 24880 38528 24886
rect 38476 24822 38528 24828
rect 38476 24200 38528 24206
rect 38476 24142 38528 24148
rect 38108 21956 38160 21962
rect 38108 21898 38160 21904
rect 38016 21004 38068 21010
rect 38016 20946 38068 20952
rect 37844 20594 37964 20622
rect 37648 17060 37700 17066
rect 37648 17002 37700 17008
rect 37464 16584 37516 16590
rect 37464 16526 37516 16532
rect 37556 16584 37608 16590
rect 37556 16526 37608 16532
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 36820 14952 36872 14958
rect 36820 14894 36872 14900
rect 36832 14346 36860 14894
rect 37004 14476 37056 14482
rect 37004 14418 37056 14424
rect 36820 14340 36872 14346
rect 36820 14282 36872 14288
rect 36820 4480 36872 4486
rect 36820 4422 36872 4428
rect 36832 4078 36860 4422
rect 37016 4282 37044 14418
rect 37004 4276 37056 4282
rect 37004 4218 37056 4224
rect 37476 4078 37504 16526
rect 37568 16114 37596 16526
rect 37556 16108 37608 16114
rect 37556 16050 37608 16056
rect 37660 4758 37688 17002
rect 37844 15706 37872 20594
rect 38028 19922 38056 20946
rect 38016 19916 38068 19922
rect 38016 19858 38068 19864
rect 37832 15700 37884 15706
rect 37832 15642 37884 15648
rect 38120 15638 38148 21898
rect 38384 21548 38436 21554
rect 38384 21490 38436 21496
rect 38396 20602 38424 21490
rect 38384 20596 38436 20602
rect 38384 20538 38436 20544
rect 38200 16448 38252 16454
rect 38200 16390 38252 16396
rect 38212 16114 38240 16390
rect 38200 16108 38252 16114
rect 38200 16050 38252 16056
rect 38384 15972 38436 15978
rect 38384 15914 38436 15920
rect 38108 15632 38160 15638
rect 38108 15574 38160 15580
rect 38120 14958 38148 15574
rect 38108 14952 38160 14958
rect 38108 14894 38160 14900
rect 37648 4752 37700 4758
rect 37648 4694 37700 4700
rect 36820 4072 36872 4078
rect 36820 4014 36872 4020
rect 37464 4072 37516 4078
rect 37464 4014 37516 4020
rect 36636 3596 36688 3602
rect 36636 3538 36688 3544
rect 36360 3460 36412 3466
rect 36360 3402 36412 3408
rect 36176 3052 36228 3058
rect 36176 2994 36228 3000
rect 36268 2916 36320 2922
rect 36268 2858 36320 2864
rect 36280 2514 36308 2858
rect 35360 2468 35480 2496
rect 36084 2508 36136 2514
rect 35360 2310 35388 2468
rect 36084 2450 36136 2456
rect 36268 2508 36320 2514
rect 36268 2450 36320 2456
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 35348 2304 35400 2310
rect 35348 2246 35400 2252
rect 35452 800 35480 2314
rect 36372 800 36400 3402
rect 36452 3392 36504 3398
rect 36452 3334 36504 3340
rect 36464 2990 36492 3334
rect 36544 3120 36596 3126
rect 36544 3062 36596 3068
rect 36452 2984 36504 2990
rect 36452 2926 36504 2932
rect 36464 2378 36492 2926
rect 36556 2514 36584 3062
rect 36544 2508 36596 2514
rect 36544 2450 36596 2456
rect 36452 2372 36504 2378
rect 36452 2314 36504 2320
rect 36832 800 36860 4014
rect 37372 4004 37424 4010
rect 37372 3946 37424 3952
rect 37384 3602 37412 3946
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 37660 2990 37688 4694
rect 38200 3936 38252 3942
rect 38200 3878 38252 3884
rect 38212 3602 38240 3878
rect 38200 3596 38252 3602
rect 38200 3538 38252 3544
rect 37832 3120 37884 3126
rect 37832 3062 37884 3068
rect 37648 2984 37700 2990
rect 37648 2926 37700 2932
rect 37372 2644 37424 2650
rect 37372 2586 37424 2592
rect 37280 2304 37332 2310
rect 37280 2246 37332 2252
rect 37292 800 37320 2246
rect 37384 2106 37412 2586
rect 37844 2514 37872 3062
rect 37832 2508 37884 2514
rect 37832 2450 37884 2456
rect 37372 2100 37424 2106
rect 37372 2042 37424 2048
rect 38212 800 38240 3538
rect 38292 3392 38344 3398
rect 38292 3334 38344 3340
rect 38304 2990 38332 3334
rect 38396 3126 38424 15914
rect 38488 4622 38516 24142
rect 38580 21962 38608 25298
rect 38568 21956 38620 21962
rect 38568 21898 38620 21904
rect 38660 15496 38712 15502
rect 38660 15438 38712 15444
rect 38672 8362 38700 15438
rect 38660 8356 38712 8362
rect 38660 8298 38712 8304
rect 38476 4616 38528 4622
rect 38476 4558 38528 4564
rect 38660 3936 38712 3942
rect 38660 3878 38712 3884
rect 38672 3602 38700 3878
rect 38764 3738 38792 25434
rect 38856 21010 38884 26182
rect 39132 25294 39160 27270
rect 39316 27062 39344 27474
rect 39764 27464 39816 27470
rect 39764 27406 39816 27412
rect 39304 27056 39356 27062
rect 39304 26998 39356 27004
rect 39776 26874 39804 27406
rect 39868 27062 39896 27934
rect 39856 27056 39908 27062
rect 39856 26998 39908 27004
rect 40052 26926 40080 29200
rect 40132 27600 40184 27606
rect 40132 27542 40184 27548
rect 39856 26920 39908 26926
rect 39776 26868 39856 26874
rect 39776 26862 39908 26868
rect 40040 26920 40092 26926
rect 40040 26862 40092 26868
rect 39776 26846 39896 26862
rect 39484 26684 39780 26704
rect 39540 26682 39564 26684
rect 39620 26682 39644 26684
rect 39700 26682 39724 26684
rect 39562 26630 39564 26682
rect 39626 26630 39638 26682
rect 39700 26630 39702 26682
rect 39540 26628 39564 26630
rect 39620 26628 39644 26630
rect 39700 26628 39724 26630
rect 39484 26608 39780 26628
rect 39868 26518 39896 26846
rect 39396 26512 39448 26518
rect 39396 26454 39448 26460
rect 39856 26512 39908 26518
rect 39856 26454 39908 26460
rect 39408 25362 39436 26454
rect 40144 26042 40172 27542
rect 40224 27532 40276 27538
rect 40224 27474 40276 27480
rect 40132 26036 40184 26042
rect 40132 25978 40184 25984
rect 39856 25832 39908 25838
rect 39856 25774 39908 25780
rect 39948 25832 40000 25838
rect 39948 25774 40000 25780
rect 39484 25596 39780 25616
rect 39540 25594 39564 25596
rect 39620 25594 39644 25596
rect 39700 25594 39724 25596
rect 39562 25542 39564 25594
rect 39626 25542 39638 25594
rect 39700 25542 39702 25594
rect 39540 25540 39564 25542
rect 39620 25540 39644 25542
rect 39700 25540 39724 25542
rect 39484 25520 39780 25540
rect 39304 25356 39356 25362
rect 39304 25298 39356 25304
rect 39396 25356 39448 25362
rect 39396 25298 39448 25304
rect 39120 25288 39172 25294
rect 39120 25230 39172 25236
rect 39212 24268 39264 24274
rect 39212 24210 39264 24216
rect 39224 23866 39252 24210
rect 39316 24206 39344 25298
rect 39408 25158 39436 25298
rect 39396 25152 39448 25158
rect 39396 25094 39448 25100
rect 39408 24818 39436 25094
rect 39396 24812 39448 24818
rect 39396 24754 39448 24760
rect 39868 24682 39896 25774
rect 39960 24886 39988 25774
rect 39948 24880 40000 24886
rect 39948 24822 40000 24828
rect 39856 24676 39908 24682
rect 39856 24618 39908 24624
rect 39484 24508 39780 24528
rect 39540 24506 39564 24508
rect 39620 24506 39644 24508
rect 39700 24506 39724 24508
rect 39562 24454 39564 24506
rect 39626 24454 39638 24506
rect 39700 24454 39702 24506
rect 39540 24452 39564 24454
rect 39620 24452 39644 24454
rect 39700 24452 39724 24454
rect 39484 24432 39780 24452
rect 39304 24200 39356 24206
rect 39304 24142 39356 24148
rect 39212 23860 39264 23866
rect 39212 23802 39264 23808
rect 39948 23520 40000 23526
rect 39948 23462 40000 23468
rect 39484 23420 39780 23440
rect 39540 23418 39564 23420
rect 39620 23418 39644 23420
rect 39700 23418 39724 23420
rect 39562 23366 39564 23418
rect 39626 23366 39638 23418
rect 39700 23366 39702 23418
rect 39540 23364 39564 23366
rect 39620 23364 39644 23366
rect 39700 23364 39724 23366
rect 39484 23344 39780 23364
rect 39484 22332 39780 22352
rect 39540 22330 39564 22332
rect 39620 22330 39644 22332
rect 39700 22330 39724 22332
rect 39562 22278 39564 22330
rect 39626 22278 39638 22330
rect 39700 22278 39702 22330
rect 39540 22276 39564 22278
rect 39620 22276 39644 22278
rect 39700 22276 39724 22278
rect 39484 22256 39780 22276
rect 39484 21244 39780 21264
rect 39540 21242 39564 21244
rect 39620 21242 39644 21244
rect 39700 21242 39724 21244
rect 39562 21190 39564 21242
rect 39626 21190 39638 21242
rect 39700 21190 39702 21242
rect 39540 21188 39564 21190
rect 39620 21188 39644 21190
rect 39700 21188 39724 21190
rect 39484 21168 39780 21188
rect 38844 21004 38896 21010
rect 38844 20946 38896 20952
rect 38936 20256 38988 20262
rect 38936 20198 38988 20204
rect 38948 12646 38976 20198
rect 39484 20156 39780 20176
rect 39540 20154 39564 20156
rect 39620 20154 39644 20156
rect 39700 20154 39724 20156
rect 39562 20102 39564 20154
rect 39626 20102 39638 20154
rect 39700 20102 39702 20154
rect 39540 20100 39564 20102
rect 39620 20100 39644 20102
rect 39700 20100 39724 20102
rect 39484 20080 39780 20100
rect 39484 19068 39780 19088
rect 39540 19066 39564 19068
rect 39620 19066 39644 19068
rect 39700 19066 39724 19068
rect 39562 19014 39564 19066
rect 39626 19014 39638 19066
rect 39700 19014 39702 19066
rect 39540 19012 39564 19014
rect 39620 19012 39644 19014
rect 39700 19012 39724 19014
rect 39484 18992 39780 19012
rect 39484 17980 39780 18000
rect 39540 17978 39564 17980
rect 39620 17978 39644 17980
rect 39700 17978 39724 17980
rect 39562 17926 39564 17978
rect 39626 17926 39638 17978
rect 39700 17926 39702 17978
rect 39540 17924 39564 17926
rect 39620 17924 39644 17926
rect 39700 17924 39724 17926
rect 39484 17904 39780 17924
rect 39484 16892 39780 16912
rect 39540 16890 39564 16892
rect 39620 16890 39644 16892
rect 39700 16890 39724 16892
rect 39562 16838 39564 16890
rect 39626 16838 39638 16890
rect 39700 16838 39702 16890
rect 39540 16836 39564 16838
rect 39620 16836 39644 16838
rect 39700 16836 39724 16838
rect 39484 16816 39780 16836
rect 39856 15904 39908 15910
rect 39856 15846 39908 15852
rect 39484 15804 39780 15824
rect 39540 15802 39564 15804
rect 39620 15802 39644 15804
rect 39700 15802 39724 15804
rect 39562 15750 39564 15802
rect 39626 15750 39638 15802
rect 39700 15750 39702 15802
rect 39540 15748 39564 15750
rect 39620 15748 39644 15750
rect 39700 15748 39724 15750
rect 39484 15728 39780 15748
rect 39868 15570 39896 15846
rect 39856 15564 39908 15570
rect 39856 15506 39908 15512
rect 39484 14716 39780 14736
rect 39540 14714 39564 14716
rect 39620 14714 39644 14716
rect 39700 14714 39724 14716
rect 39562 14662 39564 14714
rect 39626 14662 39638 14714
rect 39700 14662 39702 14714
rect 39540 14660 39564 14662
rect 39620 14660 39644 14662
rect 39700 14660 39724 14662
rect 39484 14640 39780 14660
rect 39484 13628 39780 13648
rect 39540 13626 39564 13628
rect 39620 13626 39644 13628
rect 39700 13626 39724 13628
rect 39562 13574 39564 13626
rect 39626 13574 39638 13626
rect 39700 13574 39702 13626
rect 39540 13572 39564 13574
rect 39620 13572 39644 13574
rect 39700 13572 39724 13574
rect 39484 13552 39780 13572
rect 38936 12640 38988 12646
rect 38936 12582 38988 12588
rect 39484 12540 39780 12560
rect 39540 12538 39564 12540
rect 39620 12538 39644 12540
rect 39700 12538 39724 12540
rect 39562 12486 39564 12538
rect 39626 12486 39638 12538
rect 39700 12486 39702 12538
rect 39540 12484 39564 12486
rect 39620 12484 39644 12486
rect 39700 12484 39724 12486
rect 39484 12464 39780 12484
rect 39484 11452 39780 11472
rect 39540 11450 39564 11452
rect 39620 11450 39644 11452
rect 39700 11450 39724 11452
rect 39562 11398 39564 11450
rect 39626 11398 39638 11450
rect 39700 11398 39702 11450
rect 39540 11396 39564 11398
rect 39620 11396 39644 11398
rect 39700 11396 39724 11398
rect 39484 11376 39780 11396
rect 39484 10364 39780 10384
rect 39540 10362 39564 10364
rect 39620 10362 39644 10364
rect 39700 10362 39724 10364
rect 39562 10310 39564 10362
rect 39626 10310 39638 10362
rect 39700 10310 39702 10362
rect 39540 10308 39564 10310
rect 39620 10308 39644 10310
rect 39700 10308 39724 10310
rect 39484 10288 39780 10308
rect 39484 9276 39780 9296
rect 39540 9274 39564 9276
rect 39620 9274 39644 9276
rect 39700 9274 39724 9276
rect 39562 9222 39564 9274
rect 39626 9222 39638 9274
rect 39700 9222 39702 9274
rect 39540 9220 39564 9222
rect 39620 9220 39644 9222
rect 39700 9220 39724 9222
rect 39484 9200 39780 9220
rect 39484 8188 39780 8208
rect 39540 8186 39564 8188
rect 39620 8186 39644 8188
rect 39700 8186 39724 8188
rect 39562 8134 39564 8186
rect 39626 8134 39638 8186
rect 39700 8134 39702 8186
rect 39540 8132 39564 8134
rect 39620 8132 39644 8134
rect 39700 8132 39724 8134
rect 39484 8112 39780 8132
rect 39484 7100 39780 7120
rect 39540 7098 39564 7100
rect 39620 7098 39644 7100
rect 39700 7098 39724 7100
rect 39562 7046 39564 7098
rect 39626 7046 39638 7098
rect 39700 7046 39702 7098
rect 39540 7044 39564 7046
rect 39620 7044 39644 7046
rect 39700 7044 39724 7046
rect 39484 7024 39780 7044
rect 39484 6012 39780 6032
rect 39540 6010 39564 6012
rect 39620 6010 39644 6012
rect 39700 6010 39724 6012
rect 39562 5958 39564 6010
rect 39626 5958 39638 6010
rect 39700 5958 39702 6010
rect 39540 5956 39564 5958
rect 39620 5956 39644 5958
rect 39700 5956 39724 5958
rect 39484 5936 39780 5956
rect 39484 4924 39780 4944
rect 39540 4922 39564 4924
rect 39620 4922 39644 4924
rect 39700 4922 39724 4924
rect 39562 4870 39564 4922
rect 39626 4870 39638 4922
rect 39700 4870 39702 4922
rect 39540 4868 39564 4870
rect 39620 4868 39644 4870
rect 39700 4868 39724 4870
rect 39484 4848 39780 4868
rect 39868 4554 39896 15506
rect 39120 4548 39172 4554
rect 39120 4490 39172 4496
rect 39856 4548 39908 4554
rect 39856 4490 39908 4496
rect 38752 3732 38804 3738
rect 38752 3674 38804 3680
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 38384 3120 38436 3126
rect 38384 3062 38436 3068
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 38672 800 38700 3538
rect 39132 2514 39160 4490
rect 39304 4480 39356 4486
rect 39304 4422 39356 4428
rect 39316 2514 39344 4422
rect 39868 4078 39896 4490
rect 39396 4072 39448 4078
rect 39396 4014 39448 4020
rect 39856 4072 39908 4078
rect 39856 4014 39908 4020
rect 39408 3942 39436 4014
rect 39396 3936 39448 3942
rect 39396 3878 39448 3884
rect 39408 3618 39436 3878
rect 39484 3836 39780 3856
rect 39540 3834 39564 3836
rect 39620 3834 39644 3836
rect 39700 3834 39724 3836
rect 39562 3782 39564 3834
rect 39626 3782 39638 3834
rect 39700 3782 39702 3834
rect 39540 3780 39564 3782
rect 39620 3780 39644 3782
rect 39700 3780 39724 3782
rect 39484 3760 39780 3780
rect 39408 3590 39528 3618
rect 39396 3460 39448 3466
rect 39396 3402 39448 3408
rect 39120 2508 39172 2514
rect 39120 2450 39172 2456
rect 39304 2508 39356 2514
rect 39304 2450 39356 2456
rect 39408 1714 39436 3402
rect 39500 2990 39528 3590
rect 39488 2984 39540 2990
rect 39488 2926 39540 2932
rect 39484 2748 39780 2768
rect 39540 2746 39564 2748
rect 39620 2746 39644 2748
rect 39700 2746 39724 2748
rect 39562 2694 39564 2746
rect 39626 2694 39638 2746
rect 39700 2694 39702 2746
rect 39540 2692 39564 2694
rect 39620 2692 39644 2694
rect 39700 2692 39724 2694
rect 39484 2672 39780 2692
rect 39764 2508 39816 2514
rect 39764 2450 39816 2456
rect 39408 1686 39620 1714
rect 39592 800 39620 1686
rect 39776 1630 39804 2450
rect 39868 2446 39896 4014
rect 39960 2854 39988 23462
rect 40236 22778 40264 27474
rect 40512 26450 40540 29200
rect 41432 27538 41460 29200
rect 41420 27532 41472 27538
rect 41420 27474 41472 27480
rect 40960 26920 41012 26926
rect 40960 26862 41012 26868
rect 40592 26852 40644 26858
rect 40592 26794 40644 26800
rect 40500 26444 40552 26450
rect 40500 26386 40552 26392
rect 40604 26382 40632 26794
rect 40592 26376 40644 26382
rect 40592 26318 40644 26324
rect 40972 26042 41000 26862
rect 41328 26784 41380 26790
rect 41328 26726 41380 26732
rect 41144 26444 41196 26450
rect 41144 26386 41196 26392
rect 41156 26042 41184 26386
rect 40316 26036 40368 26042
rect 40316 25978 40368 25984
rect 40960 26036 41012 26042
rect 40960 25978 41012 25984
rect 41144 26036 41196 26042
rect 41144 25978 41196 25984
rect 40224 22772 40276 22778
rect 40224 22714 40276 22720
rect 40132 3936 40184 3942
rect 40132 3878 40184 3884
rect 40144 3602 40172 3878
rect 40132 3596 40184 3602
rect 40132 3538 40184 3544
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 39948 2848 40000 2854
rect 39948 2790 40000 2796
rect 39856 2440 39908 2446
rect 39856 2382 39908 2388
rect 39764 1624 39816 1630
rect 39764 1566 39816 1572
rect 40052 800 40080 2994
rect 40132 2916 40184 2922
rect 40132 2858 40184 2864
rect 40144 2650 40172 2858
rect 40132 2644 40184 2650
rect 40132 2586 40184 2592
rect 40328 2106 40356 25978
rect 40684 24064 40736 24070
rect 40684 24006 40736 24012
rect 40696 23866 40724 24006
rect 40684 23860 40736 23866
rect 40684 23802 40736 23808
rect 40868 16516 40920 16522
rect 40868 16458 40920 16464
rect 40880 16114 40908 16458
rect 40868 16108 40920 16114
rect 40868 16050 40920 16056
rect 41144 16040 41196 16046
rect 41144 15982 41196 15988
rect 40408 5568 40460 5574
rect 40408 5510 40460 5516
rect 40420 2514 40448 5510
rect 40500 5024 40552 5030
rect 40500 4966 40552 4972
rect 40512 4690 40540 4966
rect 40500 4684 40552 4690
rect 40500 4626 40552 4632
rect 40408 2508 40460 2514
rect 40408 2450 40460 2456
rect 40316 2100 40368 2106
rect 40316 2042 40368 2048
rect 40512 800 40540 4626
rect 41156 4622 41184 15982
rect 41340 6454 41368 26726
rect 41432 26586 41460 27474
rect 41788 27328 41840 27334
rect 41788 27270 41840 27276
rect 41696 26988 41748 26994
rect 41696 26930 41748 26936
rect 41708 26586 41736 26930
rect 41420 26580 41472 26586
rect 41420 26522 41472 26528
rect 41696 26580 41748 26586
rect 41696 26522 41748 26528
rect 41604 26036 41656 26042
rect 41604 25978 41656 25984
rect 41616 25838 41644 25978
rect 41604 25832 41656 25838
rect 41604 25774 41656 25780
rect 41420 15496 41472 15502
rect 41420 15438 41472 15444
rect 41432 11218 41460 15438
rect 41420 11212 41472 11218
rect 41420 11154 41472 11160
rect 41800 8430 41828 27270
rect 41892 27062 41920 29200
rect 42812 27606 42840 29200
rect 43272 27674 43300 29200
rect 43260 27668 43312 27674
rect 43260 27610 43312 27616
rect 42800 27600 42852 27606
rect 43732 27588 43760 29200
rect 43812 27600 43864 27606
rect 43732 27560 43812 27588
rect 42800 27542 42852 27548
rect 43812 27542 43864 27548
rect 43536 27532 43588 27538
rect 43536 27474 43588 27480
rect 44088 27532 44140 27538
rect 44088 27474 44140 27480
rect 41880 27056 41932 27062
rect 41880 26998 41932 27004
rect 41880 26920 41932 26926
rect 41880 26862 41932 26868
rect 41892 26518 41920 26862
rect 42340 26852 42392 26858
rect 42340 26794 42392 26800
rect 41880 26512 41932 26518
rect 41880 26454 41932 26460
rect 42352 26246 42380 26794
rect 42340 26240 42392 26246
rect 42340 26182 42392 26188
rect 42352 18698 42380 26182
rect 42340 18692 42392 18698
rect 42340 18634 42392 18640
rect 43548 16114 43576 27474
rect 44100 27062 44128 27474
rect 44652 27062 44680 29200
rect 44088 27056 44140 27062
rect 44086 27024 44088 27033
rect 44640 27056 44692 27062
rect 44140 27024 44142 27033
rect 44640 26998 44692 27004
rect 44086 26959 44142 26968
rect 45112 26926 45140 29200
rect 45376 28008 45428 28014
rect 45376 27950 45428 27956
rect 45388 27062 45416 27950
rect 45572 27606 45600 29200
rect 46492 27606 46520 29200
rect 46952 27606 46980 29200
rect 47032 27872 47084 27878
rect 47032 27814 47084 27820
rect 47044 27674 47072 27814
rect 47032 27668 47084 27674
rect 47032 27610 47084 27616
rect 45560 27600 45612 27606
rect 45560 27542 45612 27548
rect 46480 27600 46532 27606
rect 46480 27542 46532 27548
rect 46940 27600 46992 27606
rect 46940 27542 46992 27548
rect 45836 27532 45888 27538
rect 45836 27474 45888 27480
rect 45376 27056 45428 27062
rect 45376 26998 45428 27004
rect 45100 26920 45152 26926
rect 45100 26862 45152 26868
rect 44456 26852 44508 26858
rect 44456 26794 44508 26800
rect 44468 26246 44496 26794
rect 45848 26246 45876 27474
rect 47872 27062 47900 29200
rect 48332 27606 48360 29200
rect 48320 27600 48372 27606
rect 48792 27588 48820 29200
rect 48964 27600 49016 27606
rect 48792 27560 48964 27588
rect 48320 27542 48372 27548
rect 48964 27542 49016 27548
rect 48332 27130 48360 27542
rect 49516 27532 49568 27538
rect 49516 27474 49568 27480
rect 48412 27328 48464 27334
rect 48412 27270 48464 27276
rect 48320 27124 48372 27130
rect 48320 27066 48372 27072
rect 47860 27056 47912 27062
rect 47860 26998 47912 27004
rect 47768 26852 47820 26858
rect 47768 26794 47820 26800
rect 47400 26580 47452 26586
rect 47400 26522 47452 26528
rect 44456 26240 44508 26246
rect 44456 26182 44508 26188
rect 45836 26240 45888 26246
rect 45836 26182 45888 26188
rect 44468 18766 44496 26182
rect 45744 19168 45796 19174
rect 45744 19110 45796 19116
rect 44456 18760 44508 18766
rect 44456 18702 44508 18708
rect 44548 16448 44600 16454
rect 44548 16390 44600 16396
rect 43536 16108 43588 16114
rect 43536 16050 43588 16056
rect 44560 16046 44588 16390
rect 43628 16040 43680 16046
rect 43628 15982 43680 15988
rect 44548 16040 44600 16046
rect 44548 15982 44600 15988
rect 42340 9920 42392 9926
rect 42340 9862 42392 9868
rect 41788 8424 41840 8430
rect 41788 8366 41840 8372
rect 41248 6426 41368 6454
rect 41248 4758 41276 6426
rect 41328 5228 41380 5234
rect 41328 5170 41380 5176
rect 41512 5228 41564 5234
rect 41512 5170 41564 5176
rect 41236 4752 41288 4758
rect 41236 4694 41288 4700
rect 41144 4616 41196 4622
rect 41144 4558 41196 4564
rect 41052 4548 41104 4554
rect 41052 4490 41104 4496
rect 41064 4078 41092 4490
rect 41144 4480 41196 4486
rect 41144 4422 41196 4428
rect 41052 4072 41104 4078
rect 41052 4014 41104 4020
rect 41156 3602 41184 4422
rect 41144 3596 41196 3602
rect 41144 3538 41196 3544
rect 40592 3392 40644 3398
rect 40592 3334 40644 3340
rect 40604 2990 40632 3334
rect 41248 3058 41276 4694
rect 41340 4554 41368 5170
rect 41420 4616 41472 4622
rect 41420 4558 41472 4564
rect 41328 4548 41380 4554
rect 41328 4490 41380 4496
rect 41052 3052 41104 3058
rect 41052 2994 41104 3000
rect 41236 3052 41288 3058
rect 41236 2994 41288 3000
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 41064 2938 41092 2994
rect 41340 2938 41368 4490
rect 41432 4078 41460 4558
rect 41420 4072 41472 4078
rect 41420 4014 41472 4020
rect 41420 3732 41472 3738
rect 41420 3674 41472 3680
rect 41064 2916 41368 2938
rect 41064 2910 41236 2916
rect 41288 2910 41368 2916
rect 41236 2858 41288 2864
rect 41248 2446 41276 2858
rect 41236 2440 41288 2446
rect 41236 2382 41288 2388
rect 41432 800 41460 3674
rect 41524 3058 41552 5170
rect 41604 3936 41656 3942
rect 41604 3878 41656 3884
rect 41616 3602 41644 3878
rect 41604 3596 41656 3602
rect 41604 3538 41656 3544
rect 41880 3460 41932 3466
rect 41880 3402 41932 3408
rect 41788 3392 41840 3398
rect 41788 3334 41840 3340
rect 41604 3120 41656 3126
rect 41604 3062 41656 3068
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 41524 1970 41552 2994
rect 41616 2650 41644 3062
rect 41604 2644 41656 2650
rect 41604 2586 41656 2592
rect 41616 2514 41644 2586
rect 41800 2514 41828 3334
rect 41604 2508 41656 2514
rect 41604 2450 41656 2456
rect 41788 2508 41840 2514
rect 41788 2450 41840 2456
rect 41512 1964 41564 1970
rect 41512 1906 41564 1912
rect 41892 800 41920 3402
rect 42352 3126 42380 9862
rect 42432 4480 42484 4486
rect 42432 4422 42484 4428
rect 42444 4078 42472 4422
rect 43640 4282 43668 15982
rect 44560 15570 44588 15982
rect 44548 15564 44600 15570
rect 44548 15506 44600 15512
rect 44088 4548 44140 4554
rect 44088 4490 44140 4496
rect 43628 4276 43680 4282
rect 43628 4218 43680 4224
rect 43996 4276 44048 4282
rect 43996 4218 44048 4224
rect 42432 4072 42484 4078
rect 42432 4014 42484 4020
rect 42444 3738 42472 4014
rect 43444 3936 43496 3942
rect 43444 3878 43496 3884
rect 42432 3732 42484 3738
rect 42432 3674 42484 3680
rect 43456 3602 43484 3878
rect 43640 3738 43668 4218
rect 43812 4072 43864 4078
rect 43812 4014 43864 4020
rect 43628 3732 43680 3738
rect 43628 3674 43680 3680
rect 43444 3596 43496 3602
rect 43444 3538 43496 3544
rect 42800 3392 42852 3398
rect 42800 3334 42852 3340
rect 43168 3392 43220 3398
rect 43168 3334 43220 3340
rect 42340 3120 42392 3126
rect 42340 3062 42392 3068
rect 42812 2922 42840 3334
rect 42064 2916 42116 2922
rect 42064 2858 42116 2864
rect 42800 2916 42852 2922
rect 42800 2858 42852 2864
rect 42076 2446 42104 2858
rect 42064 2440 42116 2446
rect 42064 2382 42116 2388
rect 42524 2304 42576 2310
rect 42524 2246 42576 2252
rect 42708 2304 42760 2310
rect 42708 2246 42760 2252
rect 42536 1970 42564 2246
rect 42720 2038 42748 2246
rect 42708 2032 42760 2038
rect 42708 1974 42760 1980
rect 42524 1964 42576 1970
rect 42524 1906 42576 1912
rect 42812 800 42840 2858
rect 43180 2650 43208 3334
rect 43076 2644 43128 2650
rect 43076 2586 43128 2592
rect 43168 2644 43220 2650
rect 43168 2586 43220 2592
rect 43352 2644 43404 2650
rect 43352 2586 43404 2592
rect 43088 2530 43116 2586
rect 43364 2530 43392 2586
rect 43088 2502 43392 2530
rect 43456 2428 43484 3538
rect 43720 3528 43772 3534
rect 43720 3470 43772 3476
rect 43628 3120 43680 3126
rect 43628 3062 43680 3068
rect 43640 2961 43668 3062
rect 43626 2952 43682 2961
rect 43626 2887 43682 2896
rect 43272 2400 43484 2428
rect 43272 800 43300 2400
rect 43732 800 43760 3470
rect 43824 2446 43852 4014
rect 44008 3602 44036 4218
rect 44100 4078 44128 4490
rect 44640 4480 44692 4486
rect 44640 4422 44692 4428
rect 44272 4140 44324 4146
rect 44272 4082 44324 4088
rect 44088 4072 44140 4078
rect 44088 4014 44140 4020
rect 43996 3596 44048 3602
rect 43996 3538 44048 3544
rect 43996 3460 44048 3466
rect 43996 3402 44048 3408
rect 44008 2854 44036 3402
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 44100 3058 44128 3334
rect 44088 3052 44140 3058
rect 44088 2994 44140 3000
rect 44180 2916 44232 2922
rect 44180 2858 44232 2864
rect 43996 2848 44048 2854
rect 43996 2790 44048 2796
rect 44192 2446 44220 2858
rect 44284 2854 44312 4082
rect 44652 3942 44680 4422
rect 45468 4004 45520 4010
rect 45468 3946 45520 3952
rect 45560 4004 45612 4010
rect 45560 3946 45612 3952
rect 44548 3936 44600 3942
rect 44548 3878 44600 3884
rect 44640 3936 44692 3942
rect 44640 3878 44692 3884
rect 44272 2848 44324 2854
rect 44272 2790 44324 2796
rect 44364 2848 44416 2854
rect 44364 2790 44416 2796
rect 44376 2650 44404 2790
rect 44364 2644 44416 2650
rect 44364 2586 44416 2592
rect 44560 2514 44588 3878
rect 45480 3126 45508 3946
rect 45468 3120 45520 3126
rect 45468 3062 45520 3068
rect 45100 2984 45152 2990
rect 45100 2926 45152 2932
rect 44640 2916 44692 2922
rect 44640 2858 44692 2864
rect 44916 2916 44968 2922
rect 44916 2858 44968 2864
rect 44548 2508 44600 2514
rect 44548 2450 44600 2456
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 44180 2440 44232 2446
rect 44180 2382 44232 2388
rect 44652 800 44680 2858
rect 44928 2650 44956 2858
rect 44916 2644 44968 2650
rect 44916 2586 44968 2592
rect 44916 2508 44968 2514
rect 44916 2450 44968 2456
rect 44928 1562 44956 2450
rect 44916 1556 44968 1562
rect 44916 1498 44968 1504
rect 45112 800 45140 2926
rect 45572 2514 45600 3946
rect 45756 2514 45784 19110
rect 45848 15910 45876 26182
rect 47216 21004 47268 21010
rect 47216 20946 47268 20952
rect 47228 20806 47256 20946
rect 47412 20942 47440 26522
rect 47400 20936 47452 20942
rect 47400 20878 47452 20884
rect 47216 20800 47268 20806
rect 47216 20742 47268 20748
rect 45836 15904 45888 15910
rect 45836 15846 45888 15852
rect 47228 15609 47256 20742
rect 47412 20602 47440 20878
rect 47780 20806 47808 26794
rect 47860 26784 47912 26790
rect 47860 26726 47912 26732
rect 47872 25226 47900 26726
rect 47860 25220 47912 25226
rect 47860 25162 47912 25168
rect 47768 20800 47820 20806
rect 47768 20742 47820 20748
rect 47400 20596 47452 20602
rect 47400 20538 47452 20544
rect 47214 15600 47270 15609
rect 47214 15535 47270 15544
rect 48424 4146 48452 27270
rect 49116 27228 49412 27248
rect 49172 27226 49196 27228
rect 49252 27226 49276 27228
rect 49332 27226 49356 27228
rect 49194 27174 49196 27226
rect 49258 27174 49270 27226
rect 49332 27174 49334 27226
rect 49172 27172 49196 27174
rect 49252 27172 49276 27174
rect 49332 27172 49356 27174
rect 49116 27152 49412 27172
rect 49422 26344 49478 26353
rect 49528 26330 49556 27474
rect 49712 27062 49740 29200
rect 50172 27062 50200 29200
rect 50436 27532 50488 27538
rect 50436 27474 50488 27480
rect 49700 27056 49752 27062
rect 49700 26998 49752 27004
rect 50160 27056 50212 27062
rect 50160 26998 50212 27004
rect 49976 26852 50028 26858
rect 49976 26794 50028 26800
rect 49478 26302 49556 26330
rect 49422 26279 49424 26288
rect 49476 26279 49478 26288
rect 49424 26250 49476 26256
rect 49988 26246 50016 26794
rect 49976 26240 50028 26246
rect 49976 26182 50028 26188
rect 49116 26140 49412 26160
rect 49172 26138 49196 26140
rect 49252 26138 49276 26140
rect 49332 26138 49356 26140
rect 49194 26086 49196 26138
rect 49258 26086 49270 26138
rect 49332 26086 49334 26138
rect 49172 26084 49196 26086
rect 49252 26084 49276 26086
rect 49332 26084 49356 26086
rect 49116 26064 49412 26084
rect 49116 25052 49412 25072
rect 49172 25050 49196 25052
rect 49252 25050 49276 25052
rect 49332 25050 49356 25052
rect 49194 24998 49196 25050
rect 49258 24998 49270 25050
rect 49332 24998 49334 25050
rect 49172 24996 49196 24998
rect 49252 24996 49276 24998
rect 49332 24996 49356 24998
rect 49116 24976 49412 24996
rect 49116 23964 49412 23984
rect 49172 23962 49196 23964
rect 49252 23962 49276 23964
rect 49332 23962 49356 23964
rect 49194 23910 49196 23962
rect 49258 23910 49270 23962
rect 49332 23910 49334 23962
rect 49172 23908 49196 23910
rect 49252 23908 49276 23910
rect 49332 23908 49356 23910
rect 49116 23888 49412 23908
rect 49116 22876 49412 22896
rect 49172 22874 49196 22876
rect 49252 22874 49276 22876
rect 49332 22874 49356 22876
rect 49194 22822 49196 22874
rect 49258 22822 49270 22874
rect 49332 22822 49334 22874
rect 49172 22820 49196 22822
rect 49252 22820 49276 22822
rect 49332 22820 49356 22822
rect 49116 22800 49412 22820
rect 49116 21788 49412 21808
rect 49172 21786 49196 21788
rect 49252 21786 49276 21788
rect 49332 21786 49356 21788
rect 49194 21734 49196 21786
rect 49258 21734 49270 21786
rect 49332 21734 49334 21786
rect 49172 21732 49196 21734
rect 49252 21732 49276 21734
rect 49332 21732 49356 21734
rect 49116 21712 49412 21732
rect 49116 20700 49412 20720
rect 49172 20698 49196 20700
rect 49252 20698 49276 20700
rect 49332 20698 49356 20700
rect 49194 20646 49196 20698
rect 49258 20646 49270 20698
rect 49332 20646 49334 20698
rect 49172 20644 49196 20646
rect 49252 20644 49276 20646
rect 49332 20644 49356 20646
rect 49116 20624 49412 20644
rect 49116 19612 49412 19632
rect 49172 19610 49196 19612
rect 49252 19610 49276 19612
rect 49332 19610 49356 19612
rect 49194 19558 49196 19610
rect 49258 19558 49270 19610
rect 49332 19558 49334 19610
rect 49172 19556 49196 19558
rect 49252 19556 49276 19558
rect 49332 19556 49356 19558
rect 49116 19536 49412 19556
rect 49116 18524 49412 18544
rect 49172 18522 49196 18524
rect 49252 18522 49276 18524
rect 49332 18522 49356 18524
rect 49194 18470 49196 18522
rect 49258 18470 49270 18522
rect 49332 18470 49334 18522
rect 49172 18468 49196 18470
rect 49252 18468 49276 18470
rect 49332 18468 49356 18470
rect 49116 18448 49412 18468
rect 49116 17436 49412 17456
rect 49172 17434 49196 17436
rect 49252 17434 49276 17436
rect 49332 17434 49356 17436
rect 49194 17382 49196 17434
rect 49258 17382 49270 17434
rect 49332 17382 49334 17434
rect 49172 17380 49196 17382
rect 49252 17380 49276 17382
rect 49332 17380 49356 17382
rect 49116 17360 49412 17380
rect 49116 16348 49412 16368
rect 49172 16346 49196 16348
rect 49252 16346 49276 16348
rect 49332 16346 49356 16348
rect 49194 16294 49196 16346
rect 49258 16294 49270 16346
rect 49332 16294 49334 16346
rect 49172 16292 49196 16294
rect 49252 16292 49276 16294
rect 49332 16292 49356 16294
rect 49116 16272 49412 16292
rect 49116 15260 49412 15280
rect 49172 15258 49196 15260
rect 49252 15258 49276 15260
rect 49332 15258 49356 15260
rect 49194 15206 49196 15258
rect 49258 15206 49270 15258
rect 49332 15206 49334 15258
rect 49172 15204 49196 15206
rect 49252 15204 49276 15206
rect 49332 15204 49356 15206
rect 49116 15184 49412 15204
rect 49116 14172 49412 14192
rect 49172 14170 49196 14172
rect 49252 14170 49276 14172
rect 49332 14170 49356 14172
rect 49194 14118 49196 14170
rect 49258 14118 49270 14170
rect 49332 14118 49334 14170
rect 49172 14116 49196 14118
rect 49252 14116 49276 14118
rect 49332 14116 49356 14118
rect 49116 14096 49412 14116
rect 49116 13084 49412 13104
rect 49172 13082 49196 13084
rect 49252 13082 49276 13084
rect 49332 13082 49356 13084
rect 49194 13030 49196 13082
rect 49258 13030 49270 13082
rect 49332 13030 49334 13082
rect 49172 13028 49196 13030
rect 49252 13028 49276 13030
rect 49332 13028 49356 13030
rect 49116 13008 49412 13028
rect 49116 11996 49412 12016
rect 49172 11994 49196 11996
rect 49252 11994 49276 11996
rect 49332 11994 49356 11996
rect 49194 11942 49196 11994
rect 49258 11942 49270 11994
rect 49332 11942 49334 11994
rect 49172 11940 49196 11942
rect 49252 11940 49276 11942
rect 49332 11940 49356 11942
rect 49116 11920 49412 11940
rect 49116 10908 49412 10928
rect 49172 10906 49196 10908
rect 49252 10906 49276 10908
rect 49332 10906 49356 10908
rect 49194 10854 49196 10906
rect 49258 10854 49270 10906
rect 49332 10854 49334 10906
rect 49172 10852 49196 10854
rect 49252 10852 49276 10854
rect 49332 10852 49356 10854
rect 49116 10832 49412 10852
rect 49116 9820 49412 9840
rect 49172 9818 49196 9820
rect 49252 9818 49276 9820
rect 49332 9818 49356 9820
rect 49194 9766 49196 9818
rect 49258 9766 49270 9818
rect 49332 9766 49334 9818
rect 49172 9764 49196 9766
rect 49252 9764 49276 9766
rect 49332 9764 49356 9766
rect 49116 9744 49412 9764
rect 49988 9722 50016 26182
rect 50448 25974 50476 27474
rect 51092 27062 51120 29200
rect 51552 27606 51580 29200
rect 52012 27606 52040 29200
rect 52932 27674 52960 29200
rect 52920 27668 52972 27674
rect 52920 27610 52972 27616
rect 53392 27606 53420 29200
rect 54312 27606 54340 29200
rect 54772 27674 54800 29200
rect 54760 27668 54812 27674
rect 54760 27610 54812 27616
rect 55232 27606 55260 29200
rect 51540 27600 51592 27606
rect 51540 27542 51592 27548
rect 52000 27600 52052 27606
rect 52000 27542 52052 27548
rect 53380 27600 53432 27606
rect 53380 27542 53432 27548
rect 54300 27600 54352 27606
rect 54300 27542 54352 27548
rect 55220 27600 55272 27606
rect 55220 27542 55272 27548
rect 51172 27328 51224 27334
rect 51172 27270 51224 27276
rect 51080 27056 51132 27062
rect 51080 26998 51132 27004
rect 50436 25968 50488 25974
rect 50436 25910 50488 25916
rect 51184 24486 51212 27270
rect 51552 26586 51580 27542
rect 52012 27130 52040 27542
rect 52368 27328 52420 27334
rect 52368 27270 52420 27276
rect 52000 27124 52052 27130
rect 52000 27066 52052 27072
rect 51540 26580 51592 26586
rect 51540 26522 51592 26528
rect 51092 24458 51212 24486
rect 49976 9716 50028 9722
rect 49976 9658 50028 9664
rect 49116 8732 49412 8752
rect 49172 8730 49196 8732
rect 49252 8730 49276 8732
rect 49332 8730 49356 8732
rect 49194 8678 49196 8730
rect 49258 8678 49270 8730
rect 49332 8678 49334 8730
rect 49172 8676 49196 8678
rect 49252 8676 49276 8678
rect 49332 8676 49356 8678
rect 49116 8656 49412 8676
rect 49116 7644 49412 7664
rect 49172 7642 49196 7644
rect 49252 7642 49276 7644
rect 49332 7642 49356 7644
rect 49194 7590 49196 7642
rect 49258 7590 49270 7642
rect 49332 7590 49334 7642
rect 49172 7588 49196 7590
rect 49252 7588 49276 7590
rect 49332 7588 49356 7590
rect 49116 7568 49412 7588
rect 49116 6556 49412 6576
rect 49172 6554 49196 6556
rect 49252 6554 49276 6556
rect 49332 6554 49356 6556
rect 49194 6502 49196 6554
rect 49258 6502 49270 6554
rect 49332 6502 49334 6554
rect 49172 6500 49196 6502
rect 49252 6500 49276 6502
rect 49332 6500 49356 6502
rect 49116 6480 49412 6500
rect 49116 5468 49412 5488
rect 49172 5466 49196 5468
rect 49252 5466 49276 5468
rect 49332 5466 49356 5468
rect 49194 5414 49196 5466
rect 49258 5414 49270 5466
rect 49332 5414 49334 5466
rect 49172 5412 49196 5414
rect 49252 5412 49276 5414
rect 49332 5412 49356 5414
rect 49116 5392 49412 5412
rect 49116 4380 49412 4400
rect 49172 4378 49196 4380
rect 49252 4378 49276 4380
rect 49332 4378 49356 4380
rect 49194 4326 49196 4378
rect 49258 4326 49270 4378
rect 49332 4326 49334 4378
rect 49172 4324 49196 4326
rect 49252 4324 49276 4326
rect 49332 4324 49356 4326
rect 49116 4304 49412 4324
rect 48412 4140 48464 4146
rect 48412 4082 48464 4088
rect 47124 4072 47176 4078
rect 47124 4014 47176 4020
rect 46296 3936 46348 3942
rect 46296 3878 46348 3884
rect 45836 3392 45888 3398
rect 45836 3334 45888 3340
rect 46020 3392 46072 3398
rect 46020 3334 46072 3340
rect 45848 2990 45876 3334
rect 45836 2984 45888 2990
rect 45836 2926 45888 2932
rect 46032 2514 46060 3334
rect 45560 2508 45612 2514
rect 45560 2450 45612 2456
rect 45744 2508 45796 2514
rect 45744 2450 45796 2456
rect 46020 2508 46072 2514
rect 46020 2450 46072 2456
rect 46032 800 46060 2450
rect 46308 2310 46336 3878
rect 47032 3392 47084 3398
rect 47032 3334 47084 3340
rect 47044 2990 47072 3334
rect 47136 3194 47164 4014
rect 51092 4010 51120 24458
rect 52380 4554 52408 27270
rect 53392 27130 53420 27542
rect 54392 27532 54444 27538
rect 54392 27474 54444 27480
rect 56048 27532 56100 27538
rect 56048 27474 56100 27480
rect 53472 27328 53524 27334
rect 53472 27270 53524 27276
rect 53380 27124 53432 27130
rect 53380 27066 53432 27072
rect 52460 23044 52512 23050
rect 52460 22986 52512 22992
rect 52472 14550 52500 22986
rect 52460 14544 52512 14550
rect 52460 14486 52512 14492
rect 53104 14476 53156 14482
rect 53104 14418 53156 14424
rect 52368 4548 52420 4554
rect 52368 4490 52420 4496
rect 51080 4004 51132 4010
rect 51080 3946 51132 3952
rect 47308 3936 47360 3942
rect 47308 3878 47360 3884
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 47124 3188 47176 3194
rect 47124 3130 47176 3136
rect 46940 2984 46992 2990
rect 46940 2926 46992 2932
rect 47032 2984 47084 2990
rect 47032 2926 47084 2932
rect 46480 2916 46532 2922
rect 46480 2858 46532 2864
rect 46296 2304 46348 2310
rect 46296 2246 46348 2252
rect 46492 800 46520 2858
rect 46952 2650 46980 2926
rect 46940 2644 46992 2650
rect 46940 2586 46992 2592
rect 47044 2530 47072 2926
rect 46952 2502 47072 2530
rect 47320 2514 47348 3878
rect 47596 2990 47624 3878
rect 47860 3528 47912 3534
rect 47860 3470 47912 3476
rect 47584 2984 47636 2990
rect 47584 2926 47636 2932
rect 47308 2508 47360 2514
rect 46952 800 46980 2502
rect 47308 2450 47360 2456
rect 47320 1766 47348 2450
rect 47400 2440 47452 2446
rect 47400 2382 47452 2388
rect 47412 2038 47440 2382
rect 47400 2032 47452 2038
rect 47400 1974 47452 1980
rect 47308 1760 47360 1766
rect 47308 1702 47360 1708
rect 47872 800 47900 3470
rect 49608 3392 49660 3398
rect 49608 3334 49660 3340
rect 50068 3392 50120 3398
rect 50068 3334 50120 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52552 3392 52604 3398
rect 52552 3334 52604 3340
rect 49116 3292 49412 3312
rect 49172 3290 49196 3292
rect 49252 3290 49276 3292
rect 49332 3290 49356 3292
rect 49194 3238 49196 3290
rect 49258 3238 49270 3290
rect 49332 3238 49334 3290
rect 49172 3236 49196 3238
rect 49252 3236 49276 3238
rect 49332 3236 49356 3238
rect 49116 3216 49412 3236
rect 48320 2916 48372 2922
rect 48320 2858 48372 2864
rect 48332 800 48360 2858
rect 49620 2650 49648 3334
rect 49700 3120 49752 3126
rect 49698 3088 49700 3097
rect 49752 3088 49754 3097
rect 49698 3023 49754 3032
rect 50080 2990 50108 3334
rect 50804 3120 50856 3126
rect 50804 3062 50856 3068
rect 49700 2984 49752 2990
rect 49700 2926 49752 2932
rect 50068 2984 50120 2990
rect 50068 2926 50120 2932
rect 49608 2644 49660 2650
rect 49608 2586 49660 2592
rect 48412 2508 48464 2514
rect 48412 2450 48464 2456
rect 49516 2508 49568 2514
rect 49516 2450 49568 2456
rect 48424 1970 48452 2450
rect 49528 2310 49556 2450
rect 48504 2304 48556 2310
rect 48504 2246 48556 2252
rect 49516 2304 49568 2310
rect 49516 2246 49568 2252
rect 48516 2106 48544 2246
rect 49116 2204 49412 2224
rect 49172 2202 49196 2204
rect 49252 2202 49276 2204
rect 49332 2202 49356 2204
rect 49194 2150 49196 2202
rect 49258 2150 49270 2202
rect 49332 2150 49334 2202
rect 49172 2148 49196 2150
rect 49252 2148 49276 2150
rect 49332 2148 49356 2150
rect 49116 2128 49412 2148
rect 48504 2100 48556 2106
rect 48504 2042 48556 2048
rect 48412 1964 48464 1970
rect 48412 1906 48464 1912
rect 49528 1578 49556 2246
rect 49252 1550 49556 1578
rect 49252 800 49280 1550
rect 49712 800 49740 2926
rect 50160 2916 50212 2922
rect 50160 2858 50212 2864
rect 50620 2916 50672 2922
rect 50620 2858 50672 2864
rect 50172 800 50200 2858
rect 50528 2508 50580 2514
rect 50528 2450 50580 2456
rect 50540 1698 50568 2450
rect 50632 2310 50660 2858
rect 50816 2650 50844 3062
rect 51540 2916 51592 2922
rect 51540 2858 51592 2864
rect 50804 2644 50856 2650
rect 50804 2586 50856 2592
rect 51080 2644 51132 2650
rect 51080 2586 51132 2592
rect 50816 2446 50844 2586
rect 50804 2440 50856 2446
rect 50804 2382 50856 2388
rect 50620 2304 50672 2310
rect 50620 2246 50672 2252
rect 50528 1692 50580 1698
rect 50528 1634 50580 1640
rect 51092 800 51120 2586
rect 51552 800 51580 2858
rect 52276 2848 52328 2854
rect 52276 2790 52328 2796
rect 52288 2582 52316 2790
rect 52276 2576 52328 2582
rect 52276 2518 52328 2524
rect 52380 2514 52408 3334
rect 52564 2990 52592 3334
rect 53116 3194 53144 14418
rect 53484 5574 53512 27270
rect 54404 26926 54432 27474
rect 55128 27396 55180 27402
rect 55128 27338 55180 27344
rect 54392 26920 54444 26926
rect 54390 26888 54392 26897
rect 54444 26888 54446 26897
rect 54390 26823 54446 26832
rect 54668 26852 54720 26858
rect 54668 26794 54720 26800
rect 54680 26586 54708 26794
rect 54668 26580 54720 26586
rect 54668 26522 54720 26528
rect 54392 24948 54444 24954
rect 54392 24890 54444 24896
rect 54404 21010 54432 24890
rect 54680 24486 54708 26522
rect 55140 26518 55168 27338
rect 55496 26784 55548 26790
rect 55496 26726 55548 26732
rect 55680 26784 55732 26790
rect 55680 26726 55732 26732
rect 55128 26512 55180 26518
rect 55126 26480 55128 26489
rect 55180 26480 55182 26489
rect 55036 26444 55088 26450
rect 55126 26415 55182 26424
rect 55036 26386 55088 26392
rect 55048 25974 55076 26386
rect 55508 26042 55536 26726
rect 55496 26036 55548 26042
rect 55496 25978 55548 25984
rect 55036 25968 55088 25974
rect 55036 25910 55088 25916
rect 55048 24486 55076 25910
rect 55692 25158 55720 26726
rect 56060 25906 56088 27474
rect 56152 27062 56180 29200
rect 56140 27056 56192 27062
rect 56140 26998 56192 27004
rect 56612 26518 56640 29200
rect 57532 27062 57560 29200
rect 57992 27606 58020 29200
rect 58162 28656 58218 28665
rect 58162 28591 58218 28600
rect 57980 27600 58032 27606
rect 57980 27542 58032 27548
rect 57612 27328 57664 27334
rect 57612 27270 57664 27276
rect 57520 27056 57572 27062
rect 57520 26998 57572 27004
rect 56600 26512 56652 26518
rect 56600 26454 56652 26460
rect 56968 26444 57020 26450
rect 56968 26386 57020 26392
rect 56048 25900 56100 25906
rect 56048 25842 56100 25848
rect 56692 25764 56744 25770
rect 56692 25706 56744 25712
rect 55680 25152 55732 25158
rect 55680 25094 55732 25100
rect 55692 24886 55720 25094
rect 56704 24954 56732 25706
rect 56876 25424 56928 25430
rect 56876 25366 56928 25372
rect 56692 24948 56744 24954
rect 56692 24890 56744 24896
rect 56784 24948 56836 24954
rect 56784 24890 56836 24896
rect 55680 24880 55732 24886
rect 55680 24822 55732 24828
rect 54588 24458 54708 24486
rect 54956 24458 55076 24486
rect 54588 21146 54616 24458
rect 54576 21140 54628 21146
rect 54576 21082 54628 21088
rect 54392 21004 54444 21010
rect 54392 20946 54444 20952
rect 54404 17678 54432 20946
rect 54956 19854 54984 24458
rect 56796 21350 56824 24890
rect 56888 24410 56916 25366
rect 56980 24954 57008 26386
rect 57244 26376 57296 26382
rect 57244 26318 57296 26324
rect 57256 26042 57284 26318
rect 57244 26036 57296 26042
rect 57244 25978 57296 25984
rect 57242 25936 57298 25945
rect 57242 25871 57298 25880
rect 57256 25362 57284 25871
rect 57428 25696 57480 25702
rect 57428 25638 57480 25644
rect 57440 25498 57468 25638
rect 57428 25492 57480 25498
rect 57428 25434 57480 25440
rect 57244 25356 57296 25362
rect 57244 25298 57296 25304
rect 56968 24948 57020 24954
rect 56968 24890 57020 24896
rect 57624 24486 57652 27270
rect 57704 26852 57756 26858
rect 57704 26794 57756 26800
rect 57532 24458 57652 24486
rect 56876 24404 56928 24410
rect 56876 24346 56928 24352
rect 57336 21956 57388 21962
rect 57336 21898 57388 21904
rect 56784 21344 56836 21350
rect 56784 21286 56836 21292
rect 57348 20874 57376 21898
rect 57336 20868 57388 20874
rect 57336 20810 57388 20816
rect 54944 19848 54996 19854
rect 54944 19790 54996 19796
rect 57336 19168 57388 19174
rect 57336 19110 57388 19116
rect 57152 18692 57204 18698
rect 57152 18634 57204 18640
rect 54392 17672 54444 17678
rect 54392 17614 54444 17620
rect 54404 17338 54432 17614
rect 54944 17536 54996 17542
rect 54944 17478 54996 17484
rect 54392 17332 54444 17338
rect 54392 17274 54444 17280
rect 54404 14550 54432 17274
rect 54392 14544 54444 14550
rect 54392 14486 54444 14492
rect 54404 14278 54432 14486
rect 54392 14272 54444 14278
rect 54392 14214 54444 14220
rect 54024 6656 54076 6662
rect 54024 6598 54076 6604
rect 53472 5568 53524 5574
rect 53472 5510 53524 5516
rect 53196 3392 53248 3398
rect 53196 3334 53248 3340
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 53104 3188 53156 3194
rect 53104 3130 53156 3136
rect 53208 2990 53236 3334
rect 52552 2984 52604 2990
rect 52552 2926 52604 2932
rect 52920 2984 52972 2990
rect 52920 2926 52972 2932
rect 53196 2984 53248 2990
rect 53196 2926 53248 2932
rect 52564 2590 52592 2926
rect 52472 2562 52592 2590
rect 52368 2508 52420 2514
rect 52368 2450 52420 2456
rect 52380 1834 52408 2450
rect 52368 1828 52420 1834
rect 52368 1770 52420 1776
rect 52472 800 52500 2562
rect 52932 800 52960 2926
rect 53392 2514 53420 3334
rect 54036 2990 54064 6598
rect 54208 3460 54260 3466
rect 54208 3402 54260 3408
rect 54220 2990 54248 3402
rect 54956 2990 54984 17478
rect 56324 14272 56376 14278
rect 56324 14214 56376 14220
rect 55128 13728 55180 13734
rect 55128 13670 55180 13676
rect 55140 4146 55168 13670
rect 56336 11606 56364 14214
rect 56336 11578 56456 11606
rect 56428 11150 56456 11578
rect 56416 11144 56468 11150
rect 56416 11086 56468 11092
rect 56428 10470 56456 11086
rect 56416 10464 56468 10470
rect 56416 10406 56468 10412
rect 56428 5234 56456 10406
rect 56876 5772 56928 5778
rect 56876 5714 56928 5720
rect 56416 5228 56468 5234
rect 56416 5170 56468 5176
rect 55128 4140 55180 4146
rect 55128 4082 55180 4088
rect 55588 3936 55640 3942
rect 55588 3878 55640 3884
rect 55600 3126 55628 3878
rect 55680 3392 55732 3398
rect 55680 3334 55732 3340
rect 56324 3392 56376 3398
rect 56324 3334 56376 3340
rect 55588 3120 55640 3126
rect 55588 3062 55640 3068
rect 54024 2984 54076 2990
rect 54024 2926 54076 2932
rect 54208 2984 54260 2990
rect 54208 2926 54260 2932
rect 54944 2984 54996 2990
rect 54944 2926 54996 2932
rect 54760 2916 54812 2922
rect 54760 2858 54812 2864
rect 54116 2848 54168 2854
rect 54116 2790 54168 2796
rect 54128 2582 54156 2790
rect 54116 2576 54168 2582
rect 54116 2518 54168 2524
rect 53380 2508 53432 2514
rect 53380 2450 53432 2456
rect 53392 800 53420 2450
rect 54300 2372 54352 2378
rect 54300 2314 54352 2320
rect 53472 2304 53524 2310
rect 53472 2246 53524 2252
rect 53484 1902 53512 2246
rect 53472 1896 53524 1902
rect 53472 1838 53524 1844
rect 54312 800 54340 2314
rect 54772 800 54800 2858
rect 55600 2582 55628 3062
rect 55588 2576 55640 2582
rect 55588 2518 55640 2524
rect 55692 2514 55720 3334
rect 56336 2990 56364 3334
rect 56428 3194 56456 5170
rect 56692 5092 56744 5098
rect 56692 5034 56744 5040
rect 56416 3188 56468 3194
rect 56416 3130 56468 3136
rect 56324 2984 56376 2990
rect 56324 2926 56376 2932
rect 56336 2590 56364 2926
rect 56508 2916 56560 2922
rect 56508 2858 56560 2864
rect 56336 2562 56456 2590
rect 55680 2508 55732 2514
rect 55680 2450 55732 2456
rect 55692 800 55720 2450
rect 56140 2372 56192 2378
rect 56140 2314 56192 2320
rect 55864 2304 55916 2310
rect 55864 2246 55916 2252
rect 55876 1970 55904 2246
rect 55864 1964 55916 1970
rect 55864 1906 55916 1912
rect 56152 800 56180 2314
rect 56428 2145 56456 2562
rect 56414 2136 56470 2145
rect 56414 2071 56470 2080
rect 56520 1766 56548 2858
rect 56600 2848 56652 2854
rect 56600 2790 56652 2796
rect 56508 1760 56560 1766
rect 56508 1702 56560 1708
rect 56612 800 56640 2790
rect 56704 2038 56732 5034
rect 56888 4826 56916 5714
rect 57060 5568 57112 5574
rect 57060 5510 57112 5516
rect 56876 4820 56928 4826
rect 56876 4762 56928 4768
rect 57072 3602 57100 5510
rect 57060 3596 57112 3602
rect 57060 3538 57112 3544
rect 57164 3194 57192 18634
rect 57348 16182 57376 19110
rect 57336 16176 57388 16182
rect 57336 16118 57388 16124
rect 57532 6730 57560 24458
rect 57716 16454 57744 26794
rect 57886 26616 57942 26625
rect 57886 26551 57942 26560
rect 57900 24750 57928 26551
rect 57992 25974 58020 27542
rect 58070 27296 58126 27305
rect 58070 27231 58126 27240
rect 58084 26926 58112 27231
rect 58072 26920 58124 26926
rect 58072 26862 58124 26868
rect 58084 26586 58112 26862
rect 58072 26580 58124 26586
rect 58072 26522 58124 26528
rect 58176 26518 58204 28591
rect 58164 26512 58216 26518
rect 58164 26454 58216 26460
rect 57980 25968 58032 25974
rect 57980 25910 58032 25916
rect 58072 25900 58124 25906
rect 58072 25842 58124 25848
rect 57888 24744 57940 24750
rect 57888 24686 57940 24692
rect 57886 24576 57942 24585
rect 57886 24511 57942 24520
rect 57900 24274 57928 24511
rect 57888 24268 57940 24274
rect 57888 24210 57940 24216
rect 57796 24200 57848 24206
rect 57796 24142 57848 24148
rect 57808 23526 57836 24142
rect 57980 24064 58032 24070
rect 57980 24006 58032 24012
rect 57992 23866 58020 24006
rect 57980 23860 58032 23866
rect 57980 23802 58032 23808
rect 57796 23520 57848 23526
rect 57796 23462 57848 23468
rect 57888 21956 57940 21962
rect 57888 21898 57940 21904
rect 57900 21865 57928 21898
rect 57886 21856 57942 21865
rect 57886 21791 57942 21800
rect 57796 20052 57848 20058
rect 57796 19994 57848 20000
rect 57704 16448 57756 16454
rect 57704 16390 57756 16396
rect 57808 10198 57836 19994
rect 58084 17218 58112 25842
rect 58452 25430 58480 29200
rect 59372 26994 59400 29200
rect 59360 26988 59412 26994
rect 59360 26930 59412 26936
rect 58440 25424 58492 25430
rect 58440 25366 58492 25372
rect 58162 23896 58218 23905
rect 58162 23831 58218 23840
rect 58176 23662 58204 23831
rect 58164 23656 58216 23662
rect 58164 23598 58216 23604
rect 58164 22568 58216 22574
rect 58162 22536 58164 22545
rect 58216 22536 58218 22545
rect 58162 22471 58218 22480
rect 58256 22432 58308 22438
rect 58256 22374 58308 22380
rect 58162 21176 58218 21185
rect 58162 21111 58218 21120
rect 58176 21010 58204 21111
rect 58164 21004 58216 21010
rect 58164 20946 58216 20952
rect 58162 19816 58218 19825
rect 58162 19751 58164 19760
rect 58216 19751 58218 19760
rect 58164 19722 58216 19728
rect 58164 19236 58216 19242
rect 58164 19178 58216 19184
rect 58176 19145 58204 19178
rect 58162 19136 58218 19145
rect 58162 19071 58218 19080
rect 58162 17776 58218 17785
rect 58162 17711 58164 17720
rect 58216 17711 58218 17720
rect 58164 17682 58216 17688
rect 57992 17190 58112 17218
rect 57888 17128 57940 17134
rect 57888 17070 57940 17076
rect 57900 16726 57928 17070
rect 57992 16946 58020 17190
rect 58070 17096 58126 17105
rect 58070 17031 58072 17040
rect 58124 17031 58126 17040
rect 58072 17002 58124 17008
rect 57992 16918 58112 16946
rect 57888 16720 57940 16726
rect 57888 16662 57940 16668
rect 57980 16652 58032 16658
rect 57980 16594 58032 16600
rect 57992 15978 58020 16594
rect 57980 15972 58032 15978
rect 57980 15914 58032 15920
rect 57980 14816 58032 14822
rect 57980 14758 58032 14764
rect 57992 14618 58020 14758
rect 57980 14612 58032 14618
rect 57980 14554 58032 14560
rect 57886 13016 57942 13025
rect 57886 12951 57942 12960
rect 57900 12850 57928 12951
rect 57888 12844 57940 12850
rect 57888 12786 57940 12792
rect 57888 11620 57940 11626
rect 57888 11562 57940 11568
rect 57900 11354 57928 11562
rect 57888 11348 57940 11354
rect 57888 11290 57940 11296
rect 58084 10962 58112 16918
rect 58164 16516 58216 16522
rect 58164 16458 58216 16464
rect 58176 16425 58204 16458
rect 58162 16416 58218 16425
rect 58162 16351 58218 16360
rect 58162 15056 58218 15065
rect 58162 14991 58218 15000
rect 58176 14958 58204 14991
rect 58164 14952 58216 14958
rect 58164 14894 58216 14900
rect 58164 14476 58216 14482
rect 58164 14418 58216 14424
rect 58176 14385 58204 14418
rect 58162 14376 58218 14385
rect 58162 14311 58218 14320
rect 58162 12336 58218 12345
rect 58162 12271 58164 12280
rect 58216 12271 58218 12280
rect 58164 12242 58216 12248
rect 58162 11656 58218 11665
rect 58162 11591 58164 11600
rect 58216 11591 58218 11600
rect 58164 11562 58216 11568
rect 58268 11286 58296 22374
rect 58256 11280 58308 11286
rect 58256 11222 58308 11228
rect 58084 10934 58296 10962
rect 58162 10296 58218 10305
rect 58162 10231 58218 10240
rect 58176 10198 58204 10231
rect 57796 10192 57848 10198
rect 57796 10134 57848 10140
rect 58164 10192 58216 10198
rect 58164 10134 58216 10140
rect 58162 9616 58218 9625
rect 58162 9551 58164 9560
rect 58216 9551 58218 9560
rect 58164 9522 58216 9528
rect 58164 8356 58216 8362
rect 58164 8298 58216 8304
rect 58176 8265 58204 8298
rect 58162 8256 58218 8265
rect 58162 8191 58218 8200
rect 58162 7576 58218 7585
rect 58162 7511 58218 7520
rect 58176 7342 58204 7511
rect 58164 7336 58216 7342
rect 58164 7278 58216 7284
rect 57888 7268 57940 7274
rect 57888 7210 57940 7216
rect 57900 6934 57928 7210
rect 57980 7200 58032 7206
rect 57980 7142 58032 7148
rect 57888 6928 57940 6934
rect 57888 6870 57940 6876
rect 57992 6866 58020 7142
rect 58070 6896 58126 6905
rect 57980 6860 58032 6866
rect 58070 6831 58072 6840
rect 57980 6802 58032 6808
rect 58124 6831 58126 6840
rect 58072 6802 58124 6808
rect 57520 6724 57572 6730
rect 57520 6666 57572 6672
rect 57704 6112 57756 6118
rect 57704 6054 57756 6060
rect 57716 5778 57744 6054
rect 57704 5772 57756 5778
rect 57704 5714 57756 5720
rect 58164 5636 58216 5642
rect 58164 5578 58216 5584
rect 58176 5545 58204 5578
rect 58162 5536 58218 5545
rect 58162 5471 58218 5480
rect 57796 5160 57848 5166
rect 57796 5102 57848 5108
rect 57612 5024 57664 5030
rect 57612 4966 57664 4972
rect 57624 4690 57652 4966
rect 57612 4684 57664 4690
rect 57612 4626 57664 4632
rect 57244 4480 57296 4486
rect 57244 4422 57296 4428
rect 57256 4282 57284 4422
rect 57244 4276 57296 4282
rect 57244 4218 57296 4224
rect 57520 3936 57572 3942
rect 57520 3878 57572 3884
rect 57244 3596 57296 3602
rect 57244 3538 57296 3544
rect 57152 3188 57204 3194
rect 57152 3130 57204 3136
rect 57256 2310 57284 3538
rect 57428 3460 57480 3466
rect 57428 3402 57480 3408
rect 57244 2304 57296 2310
rect 57244 2246 57296 2252
rect 56692 2032 56744 2038
rect 56692 1974 56744 1980
rect 57440 1714 57468 3402
rect 57532 2990 57560 3878
rect 57520 2984 57572 2990
rect 57520 2926 57572 2932
rect 57440 1686 57560 1714
rect 57532 800 57560 1686
rect 478 0 534 800
rect 938 0 994 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9678 0 9734 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11978 0 12034 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14278 0 14334 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 18418 0 18474 800
rect 18878 0 18934 800
rect 19338 0 19394 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22098 0 22154 800
rect 22558 0 22614 800
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25318 0 25374 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27158 0 27214 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29918 0 29974 800
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 33598 0 33654 800
rect 34058 0 34114 800
rect 34978 0 35034 800
rect 35438 0 35494 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 38658 0 38714 800
rect 39578 0 39634 800
rect 40038 0 40094 800
rect 40498 0 40554 800
rect 41418 0 41474 800
rect 41878 0 41934 800
rect 42798 0 42854 800
rect 43258 0 43314 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 46018 0 46074 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47858 0 47914 800
rect 48318 0 48374 800
rect 49238 0 49294 800
rect 49698 0 49754 800
rect 50158 0 50214 800
rect 51078 0 51134 800
rect 51538 0 51594 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 54758 0 54814 800
rect 55678 0 55734 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 57518 0 57574 800
rect 57624 785 57652 4626
rect 57808 4185 57836 5102
rect 58070 4856 58126 4865
rect 58070 4791 58126 4800
rect 58084 4758 58112 4791
rect 58072 4752 58124 4758
rect 58072 4694 58124 4700
rect 57888 4548 57940 4554
rect 57888 4490 57940 4496
rect 57900 4214 57928 4490
rect 58268 4282 58296 10934
rect 58256 4276 58308 4282
rect 58256 4218 58308 4224
rect 57888 4208 57940 4214
rect 57794 4176 57850 4185
rect 57888 4150 57940 4156
rect 57794 4111 57850 4120
rect 57980 4140 58032 4146
rect 57980 4082 58032 4088
rect 57796 4072 57848 4078
rect 57796 4014 57848 4020
rect 57888 4072 57940 4078
rect 57888 4014 57940 4020
rect 57808 2666 57836 4014
rect 57900 2825 57928 4014
rect 57992 3670 58020 4082
rect 57980 3664 58032 3670
rect 57980 3606 58032 3612
rect 58072 3528 58124 3534
rect 58072 3470 58124 3476
rect 57886 2816 57942 2825
rect 57886 2751 57942 2760
rect 57808 2638 58020 2666
rect 57704 2508 57756 2514
rect 57704 2450 57756 2456
rect 57716 2417 57744 2450
rect 57702 2408 57758 2417
rect 57702 2343 57758 2352
rect 57992 800 58020 2638
rect 58084 2514 58112 3470
rect 58900 3460 58952 3466
rect 58900 3402 58952 3408
rect 58072 2508 58124 2514
rect 58072 2450 58124 2456
rect 58912 800 58940 3402
rect 59360 2508 59412 2514
rect 59360 2450 59412 2456
rect 59372 800 59400 2450
rect 57610 776 57666 785
rect 57610 711 57666 720
rect 57978 0 58034 800
rect 58898 0 58954 800
rect 59358 0 59414 800
<< via2 >>
rect 1582 27376 1638 27432
rect 1490 27240 1546 27296
rect 1398 25900 1454 25936
rect 1398 25880 1400 25900
rect 1400 25880 1452 25900
rect 1452 25880 1454 25900
rect 1398 25220 1454 25256
rect 1398 25200 1400 25220
rect 1400 25200 1452 25220
rect 1452 25200 1454 25220
rect 1490 23860 1546 23896
rect 1490 23840 1492 23860
rect 1492 23840 1544 23860
rect 1544 23840 1546 23860
rect 1398 23180 1454 23216
rect 1398 23160 1400 23180
rect 1400 23160 1452 23180
rect 1452 23160 1454 23180
rect 1398 22500 1454 22536
rect 1398 22480 1400 22500
rect 1400 22480 1452 22500
rect 1452 22480 1454 22500
rect 1490 21140 1546 21176
rect 1490 21120 1492 21140
rect 1492 21120 1544 21140
rect 1544 21120 1546 21140
rect 1398 20440 1454 20496
rect 1398 19080 1454 19136
rect 1398 18400 1454 18456
rect 1398 17740 1454 17776
rect 1398 17720 1400 17740
rect 1400 17720 1452 17740
rect 1452 17720 1454 17740
rect 1398 16360 1454 16416
rect 1398 15680 1454 15736
rect 1582 15544 1638 15600
rect 1398 14320 1454 14376
rect 1398 13640 1454 13696
rect 1398 12960 1454 13016
rect 1398 11620 1454 11656
rect 1398 11600 1400 11620
rect 1400 11600 1452 11620
rect 1452 11600 1454 11620
rect 1490 10956 1492 10976
rect 1492 10956 1544 10976
rect 1544 10956 1546 10976
rect 1490 10920 1546 10956
rect 1490 9560 1546 9616
rect 1398 8900 1454 8936
rect 1398 8880 1400 8900
rect 1400 8880 1452 8900
rect 1452 8880 1454 8900
rect 1490 8236 1492 8256
rect 1492 8236 1544 8256
rect 1544 8236 1546 8256
rect 1490 8200 1546 8236
rect 1398 6840 1454 6896
rect 1398 6180 1454 6216
rect 1398 6160 1400 6180
rect 1400 6160 1452 6180
rect 1452 6160 1454 6180
rect 1398 4800 1454 4856
rect 1398 4140 1454 4176
rect 1398 4120 1400 4140
rect 1400 4120 1452 4140
rect 1452 4120 1454 4140
rect 1398 3440 1454 3496
rect 2594 28600 2650 28656
rect 2870 27920 2926 27976
rect 3330 26424 3386 26480
rect 1490 1400 1546 1456
rect 2594 2080 2650 2136
rect 5722 2916 5778 2952
rect 5722 2896 5724 2916
rect 5724 2896 5776 2916
rect 5776 2896 5778 2916
rect 5170 2352 5226 2408
rect 10588 27226 10644 27228
rect 10668 27226 10724 27228
rect 10748 27226 10804 27228
rect 10828 27226 10884 27228
rect 10588 27174 10614 27226
rect 10614 27174 10644 27226
rect 10668 27174 10678 27226
rect 10678 27174 10724 27226
rect 10748 27174 10794 27226
rect 10794 27174 10804 27226
rect 10828 27174 10858 27226
rect 10858 27174 10884 27226
rect 10588 27172 10644 27174
rect 10668 27172 10724 27174
rect 10748 27172 10804 27174
rect 10828 27172 10884 27174
rect 11058 26968 11114 27024
rect 10588 26138 10644 26140
rect 10668 26138 10724 26140
rect 10748 26138 10804 26140
rect 10828 26138 10884 26140
rect 10588 26086 10614 26138
rect 10614 26086 10644 26138
rect 10668 26086 10678 26138
rect 10678 26086 10724 26138
rect 10748 26086 10794 26138
rect 10794 26086 10804 26138
rect 10828 26086 10858 26138
rect 10858 26086 10884 26138
rect 10588 26084 10644 26086
rect 10668 26084 10724 26086
rect 10748 26084 10804 26086
rect 10828 26084 10884 26086
rect 10588 25050 10644 25052
rect 10668 25050 10724 25052
rect 10748 25050 10804 25052
rect 10828 25050 10884 25052
rect 10588 24998 10614 25050
rect 10614 24998 10644 25050
rect 10668 24998 10678 25050
rect 10678 24998 10724 25050
rect 10748 24998 10794 25050
rect 10794 24998 10804 25050
rect 10828 24998 10858 25050
rect 10858 24998 10884 25050
rect 10588 24996 10644 24998
rect 10668 24996 10724 24998
rect 10748 24996 10804 24998
rect 10828 24996 10884 24998
rect 10588 23962 10644 23964
rect 10668 23962 10724 23964
rect 10748 23962 10804 23964
rect 10828 23962 10884 23964
rect 10588 23910 10614 23962
rect 10614 23910 10644 23962
rect 10668 23910 10678 23962
rect 10678 23910 10724 23962
rect 10748 23910 10794 23962
rect 10794 23910 10804 23962
rect 10828 23910 10858 23962
rect 10858 23910 10884 23962
rect 10588 23908 10644 23910
rect 10668 23908 10724 23910
rect 10748 23908 10804 23910
rect 10828 23908 10884 23910
rect 10588 22874 10644 22876
rect 10668 22874 10724 22876
rect 10748 22874 10804 22876
rect 10828 22874 10884 22876
rect 10588 22822 10614 22874
rect 10614 22822 10644 22874
rect 10668 22822 10678 22874
rect 10678 22822 10724 22874
rect 10748 22822 10794 22874
rect 10794 22822 10804 22874
rect 10828 22822 10858 22874
rect 10858 22822 10884 22874
rect 10588 22820 10644 22822
rect 10668 22820 10724 22822
rect 10748 22820 10804 22822
rect 10828 22820 10884 22822
rect 10588 21786 10644 21788
rect 10668 21786 10724 21788
rect 10748 21786 10804 21788
rect 10828 21786 10884 21788
rect 10588 21734 10614 21786
rect 10614 21734 10644 21786
rect 10668 21734 10678 21786
rect 10678 21734 10724 21786
rect 10748 21734 10794 21786
rect 10794 21734 10804 21786
rect 10828 21734 10858 21786
rect 10858 21734 10884 21786
rect 10588 21732 10644 21734
rect 10668 21732 10724 21734
rect 10748 21732 10804 21734
rect 10828 21732 10884 21734
rect 10588 20698 10644 20700
rect 10668 20698 10724 20700
rect 10748 20698 10804 20700
rect 10828 20698 10884 20700
rect 10588 20646 10614 20698
rect 10614 20646 10644 20698
rect 10668 20646 10678 20698
rect 10678 20646 10724 20698
rect 10748 20646 10794 20698
rect 10794 20646 10804 20698
rect 10828 20646 10858 20698
rect 10858 20646 10884 20698
rect 10588 20644 10644 20646
rect 10668 20644 10724 20646
rect 10748 20644 10804 20646
rect 10828 20644 10884 20646
rect 10588 19610 10644 19612
rect 10668 19610 10724 19612
rect 10748 19610 10804 19612
rect 10828 19610 10884 19612
rect 10588 19558 10614 19610
rect 10614 19558 10644 19610
rect 10668 19558 10678 19610
rect 10678 19558 10724 19610
rect 10748 19558 10794 19610
rect 10794 19558 10804 19610
rect 10828 19558 10858 19610
rect 10858 19558 10884 19610
rect 10588 19556 10644 19558
rect 10668 19556 10724 19558
rect 10748 19556 10804 19558
rect 10828 19556 10884 19558
rect 10588 18522 10644 18524
rect 10668 18522 10724 18524
rect 10748 18522 10804 18524
rect 10828 18522 10884 18524
rect 10588 18470 10614 18522
rect 10614 18470 10644 18522
rect 10668 18470 10678 18522
rect 10678 18470 10724 18522
rect 10748 18470 10794 18522
rect 10794 18470 10804 18522
rect 10828 18470 10858 18522
rect 10858 18470 10884 18522
rect 10588 18468 10644 18470
rect 10668 18468 10724 18470
rect 10748 18468 10804 18470
rect 10828 18468 10884 18470
rect 10588 17434 10644 17436
rect 10668 17434 10724 17436
rect 10748 17434 10804 17436
rect 10828 17434 10884 17436
rect 10588 17382 10614 17434
rect 10614 17382 10644 17434
rect 10668 17382 10678 17434
rect 10678 17382 10724 17434
rect 10748 17382 10794 17434
rect 10794 17382 10804 17434
rect 10828 17382 10858 17434
rect 10858 17382 10884 17434
rect 10588 17380 10644 17382
rect 10668 17380 10724 17382
rect 10748 17380 10804 17382
rect 10828 17380 10884 17382
rect 10588 16346 10644 16348
rect 10668 16346 10724 16348
rect 10748 16346 10804 16348
rect 10828 16346 10884 16348
rect 10588 16294 10614 16346
rect 10614 16294 10644 16346
rect 10668 16294 10678 16346
rect 10678 16294 10724 16346
rect 10748 16294 10794 16346
rect 10794 16294 10804 16346
rect 10828 16294 10858 16346
rect 10858 16294 10884 16346
rect 10588 16292 10644 16294
rect 10668 16292 10724 16294
rect 10748 16292 10804 16294
rect 10828 16292 10884 16294
rect 10588 15258 10644 15260
rect 10668 15258 10724 15260
rect 10748 15258 10804 15260
rect 10828 15258 10884 15260
rect 10588 15206 10614 15258
rect 10614 15206 10644 15258
rect 10668 15206 10678 15258
rect 10678 15206 10724 15258
rect 10748 15206 10794 15258
rect 10794 15206 10804 15258
rect 10828 15206 10858 15258
rect 10858 15206 10884 15258
rect 10588 15204 10644 15206
rect 10668 15204 10724 15206
rect 10748 15204 10804 15206
rect 10828 15204 10884 15206
rect 10588 14170 10644 14172
rect 10668 14170 10724 14172
rect 10748 14170 10804 14172
rect 10828 14170 10884 14172
rect 10588 14118 10614 14170
rect 10614 14118 10644 14170
rect 10668 14118 10678 14170
rect 10678 14118 10724 14170
rect 10748 14118 10794 14170
rect 10794 14118 10804 14170
rect 10828 14118 10858 14170
rect 10858 14118 10884 14170
rect 10588 14116 10644 14118
rect 10668 14116 10724 14118
rect 10748 14116 10804 14118
rect 10828 14116 10884 14118
rect 10588 13082 10644 13084
rect 10668 13082 10724 13084
rect 10748 13082 10804 13084
rect 10828 13082 10884 13084
rect 10588 13030 10614 13082
rect 10614 13030 10644 13082
rect 10668 13030 10678 13082
rect 10678 13030 10724 13082
rect 10748 13030 10794 13082
rect 10794 13030 10804 13082
rect 10828 13030 10858 13082
rect 10858 13030 10884 13082
rect 10588 13028 10644 13030
rect 10668 13028 10724 13030
rect 10748 13028 10804 13030
rect 10828 13028 10884 13030
rect 10588 11994 10644 11996
rect 10668 11994 10724 11996
rect 10748 11994 10804 11996
rect 10828 11994 10884 11996
rect 10588 11942 10614 11994
rect 10614 11942 10644 11994
rect 10668 11942 10678 11994
rect 10678 11942 10724 11994
rect 10748 11942 10794 11994
rect 10794 11942 10804 11994
rect 10828 11942 10858 11994
rect 10858 11942 10884 11994
rect 10588 11940 10644 11942
rect 10668 11940 10724 11942
rect 10748 11940 10804 11942
rect 10828 11940 10884 11942
rect 10588 10906 10644 10908
rect 10668 10906 10724 10908
rect 10748 10906 10804 10908
rect 10828 10906 10884 10908
rect 10588 10854 10614 10906
rect 10614 10854 10644 10906
rect 10668 10854 10678 10906
rect 10678 10854 10724 10906
rect 10748 10854 10794 10906
rect 10794 10854 10804 10906
rect 10828 10854 10858 10906
rect 10858 10854 10884 10906
rect 10588 10852 10644 10854
rect 10668 10852 10724 10854
rect 10748 10852 10804 10854
rect 10828 10852 10884 10854
rect 10588 9818 10644 9820
rect 10668 9818 10724 9820
rect 10748 9818 10804 9820
rect 10828 9818 10884 9820
rect 10588 9766 10614 9818
rect 10614 9766 10644 9818
rect 10668 9766 10678 9818
rect 10678 9766 10724 9818
rect 10748 9766 10794 9818
rect 10794 9766 10804 9818
rect 10828 9766 10858 9818
rect 10858 9766 10884 9818
rect 10588 9764 10644 9766
rect 10668 9764 10724 9766
rect 10748 9764 10804 9766
rect 10828 9764 10884 9766
rect 10588 8730 10644 8732
rect 10668 8730 10724 8732
rect 10748 8730 10804 8732
rect 10828 8730 10884 8732
rect 10588 8678 10614 8730
rect 10614 8678 10644 8730
rect 10668 8678 10678 8730
rect 10678 8678 10724 8730
rect 10748 8678 10794 8730
rect 10794 8678 10804 8730
rect 10828 8678 10858 8730
rect 10858 8678 10884 8730
rect 10588 8676 10644 8678
rect 10668 8676 10724 8678
rect 10748 8676 10804 8678
rect 10828 8676 10884 8678
rect 10588 7642 10644 7644
rect 10668 7642 10724 7644
rect 10748 7642 10804 7644
rect 10828 7642 10884 7644
rect 10588 7590 10614 7642
rect 10614 7590 10644 7642
rect 10668 7590 10678 7642
rect 10678 7590 10724 7642
rect 10748 7590 10794 7642
rect 10794 7590 10804 7642
rect 10828 7590 10858 7642
rect 10858 7590 10884 7642
rect 10588 7588 10644 7590
rect 10668 7588 10724 7590
rect 10748 7588 10804 7590
rect 10828 7588 10884 7590
rect 10588 6554 10644 6556
rect 10668 6554 10724 6556
rect 10748 6554 10804 6556
rect 10828 6554 10884 6556
rect 10588 6502 10614 6554
rect 10614 6502 10644 6554
rect 10668 6502 10678 6554
rect 10678 6502 10724 6554
rect 10748 6502 10794 6554
rect 10794 6502 10804 6554
rect 10828 6502 10858 6554
rect 10858 6502 10884 6554
rect 10588 6500 10644 6502
rect 10668 6500 10724 6502
rect 10748 6500 10804 6502
rect 10828 6500 10884 6502
rect 10588 5466 10644 5468
rect 10668 5466 10724 5468
rect 10748 5466 10804 5468
rect 10828 5466 10884 5468
rect 10588 5414 10614 5466
rect 10614 5414 10644 5466
rect 10668 5414 10678 5466
rect 10678 5414 10724 5466
rect 10748 5414 10794 5466
rect 10794 5414 10804 5466
rect 10828 5414 10858 5466
rect 10858 5414 10884 5466
rect 10588 5412 10644 5414
rect 10668 5412 10724 5414
rect 10748 5412 10804 5414
rect 10828 5412 10884 5414
rect 10588 4378 10644 4380
rect 10668 4378 10724 4380
rect 10748 4378 10804 4380
rect 10828 4378 10884 4380
rect 10588 4326 10614 4378
rect 10614 4326 10644 4378
rect 10668 4326 10678 4378
rect 10678 4326 10724 4378
rect 10748 4326 10794 4378
rect 10794 4326 10804 4378
rect 10828 4326 10858 4378
rect 10858 4326 10884 4378
rect 10588 4324 10644 4326
rect 10668 4324 10724 4326
rect 10748 4324 10804 4326
rect 10828 4324 10884 4326
rect 12898 26288 12954 26344
rect 14186 26152 14242 26208
rect 10588 3290 10644 3292
rect 10668 3290 10724 3292
rect 10748 3290 10804 3292
rect 10828 3290 10884 3292
rect 10588 3238 10614 3290
rect 10614 3238 10644 3290
rect 10668 3238 10678 3290
rect 10678 3238 10724 3290
rect 10748 3238 10794 3290
rect 10794 3238 10804 3290
rect 10828 3238 10858 3290
rect 10858 3238 10884 3290
rect 10588 3236 10644 3238
rect 10668 3236 10724 3238
rect 10748 3236 10804 3238
rect 10828 3236 10884 3238
rect 10588 2202 10644 2204
rect 10668 2202 10724 2204
rect 10748 2202 10804 2204
rect 10828 2202 10884 2204
rect 10588 2150 10614 2202
rect 10614 2150 10644 2202
rect 10668 2150 10678 2202
rect 10678 2150 10724 2202
rect 10748 2150 10794 2202
rect 10794 2150 10804 2202
rect 10828 2150 10858 2202
rect 10858 2150 10884 2202
rect 10588 2148 10644 2150
rect 10668 2148 10724 2150
rect 10748 2148 10804 2150
rect 10828 2148 10884 2150
rect 12162 2624 12218 2680
rect 20220 27770 20276 27772
rect 20300 27770 20356 27772
rect 20380 27770 20436 27772
rect 20460 27770 20516 27772
rect 20220 27718 20246 27770
rect 20246 27718 20276 27770
rect 20300 27718 20310 27770
rect 20310 27718 20356 27770
rect 20380 27718 20426 27770
rect 20426 27718 20436 27770
rect 20460 27718 20490 27770
rect 20490 27718 20516 27770
rect 20220 27716 20276 27718
rect 20300 27716 20356 27718
rect 20380 27716 20436 27718
rect 20460 27716 20516 27718
rect 20220 26682 20276 26684
rect 20300 26682 20356 26684
rect 20380 26682 20436 26684
rect 20460 26682 20516 26684
rect 20220 26630 20246 26682
rect 20246 26630 20276 26682
rect 20300 26630 20310 26682
rect 20310 26630 20356 26682
rect 20380 26630 20426 26682
rect 20426 26630 20436 26682
rect 20460 26630 20490 26682
rect 20490 26630 20516 26682
rect 20220 26628 20276 26630
rect 20300 26628 20356 26630
rect 20380 26628 20436 26630
rect 20460 26628 20516 26630
rect 20994 26832 21050 26888
rect 21086 26288 21142 26344
rect 20220 25594 20276 25596
rect 20300 25594 20356 25596
rect 20380 25594 20436 25596
rect 20460 25594 20516 25596
rect 20220 25542 20246 25594
rect 20246 25542 20276 25594
rect 20300 25542 20310 25594
rect 20310 25542 20356 25594
rect 20380 25542 20426 25594
rect 20426 25542 20436 25594
rect 20460 25542 20490 25594
rect 20490 25542 20516 25594
rect 20220 25540 20276 25542
rect 20300 25540 20356 25542
rect 20380 25540 20436 25542
rect 20460 25540 20516 25542
rect 20220 24506 20276 24508
rect 20300 24506 20356 24508
rect 20380 24506 20436 24508
rect 20460 24506 20516 24508
rect 20220 24454 20246 24506
rect 20246 24454 20276 24506
rect 20300 24454 20310 24506
rect 20310 24454 20356 24506
rect 20380 24454 20426 24506
rect 20426 24454 20436 24506
rect 20460 24454 20490 24506
rect 20490 24454 20516 24506
rect 20220 24452 20276 24454
rect 20300 24452 20356 24454
rect 20380 24452 20436 24454
rect 20460 24452 20516 24454
rect 20220 23418 20276 23420
rect 20300 23418 20356 23420
rect 20380 23418 20436 23420
rect 20460 23418 20516 23420
rect 20220 23366 20246 23418
rect 20246 23366 20276 23418
rect 20300 23366 20310 23418
rect 20310 23366 20356 23418
rect 20380 23366 20426 23418
rect 20426 23366 20436 23418
rect 20460 23366 20490 23418
rect 20490 23366 20516 23418
rect 20220 23364 20276 23366
rect 20300 23364 20356 23366
rect 20380 23364 20436 23366
rect 20460 23364 20516 23366
rect 20220 22330 20276 22332
rect 20300 22330 20356 22332
rect 20380 22330 20436 22332
rect 20460 22330 20516 22332
rect 20220 22278 20246 22330
rect 20246 22278 20276 22330
rect 20300 22278 20310 22330
rect 20310 22278 20356 22330
rect 20380 22278 20426 22330
rect 20426 22278 20436 22330
rect 20460 22278 20490 22330
rect 20490 22278 20516 22330
rect 20220 22276 20276 22278
rect 20300 22276 20356 22278
rect 20380 22276 20436 22278
rect 20460 22276 20516 22278
rect 20220 21242 20276 21244
rect 20300 21242 20356 21244
rect 20380 21242 20436 21244
rect 20460 21242 20516 21244
rect 20220 21190 20246 21242
rect 20246 21190 20276 21242
rect 20300 21190 20310 21242
rect 20310 21190 20356 21242
rect 20380 21190 20426 21242
rect 20426 21190 20436 21242
rect 20460 21190 20490 21242
rect 20490 21190 20516 21242
rect 20220 21188 20276 21190
rect 20300 21188 20356 21190
rect 20380 21188 20436 21190
rect 20460 21188 20516 21190
rect 16026 3032 16082 3088
rect 15290 2644 15346 2680
rect 15290 2624 15292 2644
rect 15292 2624 15344 2644
rect 15344 2624 15346 2644
rect 20220 20154 20276 20156
rect 20300 20154 20356 20156
rect 20380 20154 20436 20156
rect 20460 20154 20516 20156
rect 20220 20102 20246 20154
rect 20246 20102 20276 20154
rect 20300 20102 20310 20154
rect 20310 20102 20356 20154
rect 20380 20102 20426 20154
rect 20426 20102 20436 20154
rect 20460 20102 20490 20154
rect 20490 20102 20516 20154
rect 20220 20100 20276 20102
rect 20300 20100 20356 20102
rect 20380 20100 20436 20102
rect 20460 20100 20516 20102
rect 20220 19066 20276 19068
rect 20300 19066 20356 19068
rect 20380 19066 20436 19068
rect 20460 19066 20516 19068
rect 20220 19014 20246 19066
rect 20246 19014 20276 19066
rect 20300 19014 20310 19066
rect 20310 19014 20356 19066
rect 20380 19014 20426 19066
rect 20426 19014 20436 19066
rect 20460 19014 20490 19066
rect 20490 19014 20516 19066
rect 20220 19012 20276 19014
rect 20300 19012 20356 19014
rect 20380 19012 20436 19014
rect 20460 19012 20516 19014
rect 20220 17978 20276 17980
rect 20300 17978 20356 17980
rect 20380 17978 20436 17980
rect 20460 17978 20516 17980
rect 20220 17926 20246 17978
rect 20246 17926 20276 17978
rect 20300 17926 20310 17978
rect 20310 17926 20356 17978
rect 20380 17926 20426 17978
rect 20426 17926 20436 17978
rect 20460 17926 20490 17978
rect 20490 17926 20516 17978
rect 20220 17924 20276 17926
rect 20300 17924 20356 17926
rect 20380 17924 20436 17926
rect 20460 17924 20516 17926
rect 20220 16890 20276 16892
rect 20300 16890 20356 16892
rect 20380 16890 20436 16892
rect 20460 16890 20516 16892
rect 20220 16838 20246 16890
rect 20246 16838 20276 16890
rect 20300 16838 20310 16890
rect 20310 16838 20356 16890
rect 20380 16838 20426 16890
rect 20426 16838 20436 16890
rect 20460 16838 20490 16890
rect 20490 16838 20516 16890
rect 20220 16836 20276 16838
rect 20300 16836 20356 16838
rect 20380 16836 20436 16838
rect 20460 16836 20516 16838
rect 20220 15802 20276 15804
rect 20300 15802 20356 15804
rect 20380 15802 20436 15804
rect 20460 15802 20516 15804
rect 20220 15750 20246 15802
rect 20246 15750 20276 15802
rect 20300 15750 20310 15802
rect 20310 15750 20356 15802
rect 20380 15750 20426 15802
rect 20426 15750 20436 15802
rect 20460 15750 20490 15802
rect 20490 15750 20516 15802
rect 20220 15748 20276 15750
rect 20300 15748 20356 15750
rect 20380 15748 20436 15750
rect 20460 15748 20516 15750
rect 20220 14714 20276 14716
rect 20300 14714 20356 14716
rect 20380 14714 20436 14716
rect 20460 14714 20516 14716
rect 20220 14662 20246 14714
rect 20246 14662 20276 14714
rect 20300 14662 20310 14714
rect 20310 14662 20356 14714
rect 20380 14662 20426 14714
rect 20426 14662 20436 14714
rect 20460 14662 20490 14714
rect 20490 14662 20516 14714
rect 20220 14660 20276 14662
rect 20300 14660 20356 14662
rect 20380 14660 20436 14662
rect 20460 14660 20516 14662
rect 20220 13626 20276 13628
rect 20300 13626 20356 13628
rect 20380 13626 20436 13628
rect 20460 13626 20516 13628
rect 20220 13574 20246 13626
rect 20246 13574 20276 13626
rect 20300 13574 20310 13626
rect 20310 13574 20356 13626
rect 20380 13574 20426 13626
rect 20426 13574 20436 13626
rect 20460 13574 20490 13626
rect 20490 13574 20516 13626
rect 20220 13572 20276 13574
rect 20300 13572 20356 13574
rect 20380 13572 20436 13574
rect 20460 13572 20516 13574
rect 20220 12538 20276 12540
rect 20300 12538 20356 12540
rect 20380 12538 20436 12540
rect 20460 12538 20516 12540
rect 20220 12486 20246 12538
rect 20246 12486 20276 12538
rect 20300 12486 20310 12538
rect 20310 12486 20356 12538
rect 20380 12486 20426 12538
rect 20426 12486 20436 12538
rect 20460 12486 20490 12538
rect 20490 12486 20516 12538
rect 20220 12484 20276 12486
rect 20300 12484 20356 12486
rect 20380 12484 20436 12486
rect 20460 12484 20516 12486
rect 20220 11450 20276 11452
rect 20300 11450 20356 11452
rect 20380 11450 20436 11452
rect 20460 11450 20516 11452
rect 20220 11398 20246 11450
rect 20246 11398 20276 11450
rect 20300 11398 20310 11450
rect 20310 11398 20356 11450
rect 20380 11398 20426 11450
rect 20426 11398 20436 11450
rect 20460 11398 20490 11450
rect 20490 11398 20516 11450
rect 20220 11396 20276 11398
rect 20300 11396 20356 11398
rect 20380 11396 20436 11398
rect 20460 11396 20516 11398
rect 20220 10362 20276 10364
rect 20300 10362 20356 10364
rect 20380 10362 20436 10364
rect 20460 10362 20516 10364
rect 20220 10310 20246 10362
rect 20246 10310 20276 10362
rect 20300 10310 20310 10362
rect 20310 10310 20356 10362
rect 20380 10310 20426 10362
rect 20426 10310 20436 10362
rect 20460 10310 20490 10362
rect 20490 10310 20516 10362
rect 20220 10308 20276 10310
rect 20300 10308 20356 10310
rect 20380 10308 20436 10310
rect 20460 10308 20516 10310
rect 20220 9274 20276 9276
rect 20300 9274 20356 9276
rect 20380 9274 20436 9276
rect 20460 9274 20516 9276
rect 20220 9222 20246 9274
rect 20246 9222 20276 9274
rect 20300 9222 20310 9274
rect 20310 9222 20356 9274
rect 20380 9222 20426 9274
rect 20426 9222 20436 9274
rect 20460 9222 20490 9274
rect 20490 9222 20516 9274
rect 20220 9220 20276 9222
rect 20300 9220 20356 9222
rect 20380 9220 20436 9222
rect 20460 9220 20516 9222
rect 20220 8186 20276 8188
rect 20300 8186 20356 8188
rect 20380 8186 20436 8188
rect 20460 8186 20516 8188
rect 20220 8134 20246 8186
rect 20246 8134 20276 8186
rect 20300 8134 20310 8186
rect 20310 8134 20356 8186
rect 20380 8134 20426 8186
rect 20426 8134 20436 8186
rect 20460 8134 20490 8186
rect 20490 8134 20516 8186
rect 20220 8132 20276 8134
rect 20300 8132 20356 8134
rect 20380 8132 20436 8134
rect 20460 8132 20516 8134
rect 20220 7098 20276 7100
rect 20300 7098 20356 7100
rect 20380 7098 20436 7100
rect 20460 7098 20516 7100
rect 20220 7046 20246 7098
rect 20246 7046 20276 7098
rect 20300 7046 20310 7098
rect 20310 7046 20356 7098
rect 20380 7046 20426 7098
rect 20426 7046 20436 7098
rect 20460 7046 20490 7098
rect 20490 7046 20516 7098
rect 20220 7044 20276 7046
rect 20300 7044 20356 7046
rect 20380 7044 20436 7046
rect 20460 7044 20516 7046
rect 20220 6010 20276 6012
rect 20300 6010 20356 6012
rect 20380 6010 20436 6012
rect 20460 6010 20516 6012
rect 20220 5958 20246 6010
rect 20246 5958 20276 6010
rect 20300 5958 20310 6010
rect 20310 5958 20356 6010
rect 20380 5958 20426 6010
rect 20426 5958 20436 6010
rect 20460 5958 20490 6010
rect 20490 5958 20516 6010
rect 20220 5956 20276 5958
rect 20300 5956 20356 5958
rect 20380 5956 20436 5958
rect 20460 5956 20516 5958
rect 20220 4922 20276 4924
rect 20300 4922 20356 4924
rect 20380 4922 20436 4924
rect 20460 4922 20516 4924
rect 20220 4870 20246 4922
rect 20246 4870 20276 4922
rect 20300 4870 20310 4922
rect 20310 4870 20356 4922
rect 20380 4870 20426 4922
rect 20426 4870 20436 4922
rect 20460 4870 20490 4922
rect 20490 4870 20516 4922
rect 20220 4868 20276 4870
rect 20300 4868 20356 4870
rect 20380 4868 20436 4870
rect 20460 4868 20516 4870
rect 20220 3834 20276 3836
rect 20300 3834 20356 3836
rect 20380 3834 20436 3836
rect 20460 3834 20516 3836
rect 20220 3782 20246 3834
rect 20246 3782 20276 3834
rect 20300 3782 20310 3834
rect 20310 3782 20356 3834
rect 20380 3782 20426 3834
rect 20426 3782 20436 3834
rect 20460 3782 20490 3834
rect 20490 3782 20516 3834
rect 20220 3780 20276 3782
rect 20300 3780 20356 3782
rect 20380 3780 20436 3782
rect 20460 3780 20516 3782
rect 20220 2746 20276 2748
rect 20300 2746 20356 2748
rect 20380 2746 20436 2748
rect 20460 2746 20516 2748
rect 20220 2694 20246 2746
rect 20246 2694 20276 2746
rect 20300 2694 20310 2746
rect 20310 2694 20356 2746
rect 20380 2694 20426 2746
rect 20426 2694 20436 2746
rect 20460 2694 20490 2746
rect 20490 2694 20516 2746
rect 20220 2692 20276 2694
rect 20300 2692 20356 2694
rect 20380 2692 20436 2694
rect 20460 2692 20516 2694
rect 24490 26152 24546 26208
rect 27986 26580 28042 26616
rect 27986 26560 27988 26580
rect 27988 26560 28040 26580
rect 28040 26560 28042 26580
rect 28170 26288 28226 26344
rect 29852 27226 29908 27228
rect 29932 27226 29988 27228
rect 30012 27226 30068 27228
rect 30092 27226 30148 27228
rect 29852 27174 29878 27226
rect 29878 27174 29908 27226
rect 29932 27174 29942 27226
rect 29942 27174 29988 27226
rect 30012 27174 30058 27226
rect 30058 27174 30068 27226
rect 30092 27174 30122 27226
rect 30122 27174 30148 27226
rect 29852 27172 29908 27174
rect 29932 27172 29988 27174
rect 30012 27172 30068 27174
rect 30092 27172 30148 27174
rect 29550 26424 29606 26480
rect 29852 26138 29908 26140
rect 29932 26138 29988 26140
rect 30012 26138 30068 26140
rect 30092 26138 30148 26140
rect 29852 26086 29878 26138
rect 29878 26086 29908 26138
rect 29932 26086 29942 26138
rect 29942 26086 29988 26138
rect 30012 26086 30058 26138
rect 30058 26086 30068 26138
rect 30092 26086 30122 26138
rect 30122 26086 30148 26138
rect 29852 26084 29908 26086
rect 29932 26084 29988 26086
rect 30012 26084 30068 26086
rect 30092 26084 30148 26086
rect 29852 25050 29908 25052
rect 29932 25050 29988 25052
rect 30012 25050 30068 25052
rect 30092 25050 30148 25052
rect 29852 24998 29878 25050
rect 29878 24998 29908 25050
rect 29932 24998 29942 25050
rect 29942 24998 29988 25050
rect 30012 24998 30058 25050
rect 30058 24998 30068 25050
rect 30092 24998 30122 25050
rect 30122 24998 30148 25050
rect 29852 24996 29908 24998
rect 29932 24996 29988 24998
rect 30012 24996 30068 24998
rect 30092 24996 30148 24998
rect 29852 23962 29908 23964
rect 29932 23962 29988 23964
rect 30012 23962 30068 23964
rect 30092 23962 30148 23964
rect 29852 23910 29878 23962
rect 29878 23910 29908 23962
rect 29932 23910 29942 23962
rect 29942 23910 29988 23962
rect 30012 23910 30058 23962
rect 30058 23910 30068 23962
rect 30092 23910 30122 23962
rect 30122 23910 30148 23962
rect 29852 23908 29908 23910
rect 29932 23908 29988 23910
rect 30012 23908 30068 23910
rect 30092 23908 30148 23910
rect 29852 22874 29908 22876
rect 29932 22874 29988 22876
rect 30012 22874 30068 22876
rect 30092 22874 30148 22876
rect 29852 22822 29878 22874
rect 29878 22822 29908 22874
rect 29932 22822 29942 22874
rect 29942 22822 29988 22874
rect 30012 22822 30058 22874
rect 30058 22822 30068 22874
rect 30092 22822 30122 22874
rect 30122 22822 30148 22874
rect 29852 22820 29908 22822
rect 29932 22820 29988 22822
rect 30012 22820 30068 22822
rect 30092 22820 30148 22822
rect 29852 21786 29908 21788
rect 29932 21786 29988 21788
rect 30012 21786 30068 21788
rect 30092 21786 30148 21788
rect 29852 21734 29878 21786
rect 29878 21734 29908 21786
rect 29932 21734 29942 21786
rect 29942 21734 29988 21786
rect 30012 21734 30058 21786
rect 30058 21734 30068 21786
rect 30092 21734 30122 21786
rect 30122 21734 30148 21786
rect 29852 21732 29908 21734
rect 29932 21732 29988 21734
rect 30012 21732 30068 21734
rect 30092 21732 30148 21734
rect 29852 20698 29908 20700
rect 29932 20698 29988 20700
rect 30012 20698 30068 20700
rect 30092 20698 30148 20700
rect 29852 20646 29878 20698
rect 29878 20646 29908 20698
rect 29932 20646 29942 20698
rect 29942 20646 29988 20698
rect 30012 20646 30058 20698
rect 30058 20646 30068 20698
rect 30092 20646 30122 20698
rect 30122 20646 30148 20698
rect 29852 20644 29908 20646
rect 29932 20644 29988 20646
rect 30012 20644 30068 20646
rect 30092 20644 30148 20646
rect 29852 19610 29908 19612
rect 29932 19610 29988 19612
rect 30012 19610 30068 19612
rect 30092 19610 30148 19612
rect 29852 19558 29878 19610
rect 29878 19558 29908 19610
rect 29932 19558 29942 19610
rect 29942 19558 29988 19610
rect 30012 19558 30058 19610
rect 30058 19558 30068 19610
rect 30092 19558 30122 19610
rect 30122 19558 30148 19610
rect 29852 19556 29908 19558
rect 29932 19556 29988 19558
rect 30012 19556 30068 19558
rect 30092 19556 30148 19558
rect 29852 18522 29908 18524
rect 29932 18522 29988 18524
rect 30012 18522 30068 18524
rect 30092 18522 30148 18524
rect 29852 18470 29878 18522
rect 29878 18470 29908 18522
rect 29932 18470 29942 18522
rect 29942 18470 29988 18522
rect 30012 18470 30058 18522
rect 30058 18470 30068 18522
rect 30092 18470 30122 18522
rect 30122 18470 30148 18522
rect 29852 18468 29908 18470
rect 29932 18468 29988 18470
rect 30012 18468 30068 18470
rect 30092 18468 30148 18470
rect 29852 17434 29908 17436
rect 29932 17434 29988 17436
rect 30012 17434 30068 17436
rect 30092 17434 30148 17436
rect 29852 17382 29878 17434
rect 29878 17382 29908 17434
rect 29932 17382 29942 17434
rect 29942 17382 29988 17434
rect 30012 17382 30058 17434
rect 30058 17382 30068 17434
rect 30092 17382 30122 17434
rect 30122 17382 30148 17434
rect 29852 17380 29908 17382
rect 29932 17380 29988 17382
rect 30012 17380 30068 17382
rect 30092 17380 30148 17382
rect 29852 16346 29908 16348
rect 29932 16346 29988 16348
rect 30012 16346 30068 16348
rect 30092 16346 30148 16348
rect 29852 16294 29878 16346
rect 29878 16294 29908 16346
rect 29932 16294 29942 16346
rect 29942 16294 29988 16346
rect 30012 16294 30058 16346
rect 30058 16294 30068 16346
rect 30092 16294 30122 16346
rect 30122 16294 30148 16346
rect 29852 16292 29908 16294
rect 29932 16292 29988 16294
rect 30012 16292 30068 16294
rect 30092 16292 30148 16294
rect 29852 15258 29908 15260
rect 29932 15258 29988 15260
rect 30012 15258 30068 15260
rect 30092 15258 30148 15260
rect 29852 15206 29878 15258
rect 29878 15206 29908 15258
rect 29932 15206 29942 15258
rect 29942 15206 29988 15258
rect 30012 15206 30058 15258
rect 30058 15206 30068 15258
rect 30092 15206 30122 15258
rect 30122 15206 30148 15258
rect 29852 15204 29908 15206
rect 29932 15204 29988 15206
rect 30012 15204 30068 15206
rect 30092 15204 30148 15206
rect 29852 14170 29908 14172
rect 29932 14170 29988 14172
rect 30012 14170 30068 14172
rect 30092 14170 30148 14172
rect 29852 14118 29878 14170
rect 29878 14118 29908 14170
rect 29932 14118 29942 14170
rect 29942 14118 29988 14170
rect 30012 14118 30058 14170
rect 30058 14118 30068 14170
rect 30092 14118 30122 14170
rect 30122 14118 30148 14170
rect 29852 14116 29908 14118
rect 29932 14116 29988 14118
rect 30012 14116 30068 14118
rect 30092 14116 30148 14118
rect 29852 13082 29908 13084
rect 29932 13082 29988 13084
rect 30012 13082 30068 13084
rect 30092 13082 30148 13084
rect 29852 13030 29878 13082
rect 29878 13030 29908 13082
rect 29932 13030 29942 13082
rect 29942 13030 29988 13082
rect 30012 13030 30058 13082
rect 30058 13030 30068 13082
rect 30092 13030 30122 13082
rect 30122 13030 30148 13082
rect 29852 13028 29908 13030
rect 29932 13028 29988 13030
rect 30012 13028 30068 13030
rect 30092 13028 30148 13030
rect 29852 11994 29908 11996
rect 29932 11994 29988 11996
rect 30012 11994 30068 11996
rect 30092 11994 30148 11996
rect 29852 11942 29878 11994
rect 29878 11942 29908 11994
rect 29932 11942 29942 11994
rect 29942 11942 29988 11994
rect 30012 11942 30058 11994
rect 30058 11942 30068 11994
rect 30092 11942 30122 11994
rect 30122 11942 30148 11994
rect 29852 11940 29908 11942
rect 29932 11940 29988 11942
rect 30012 11940 30068 11942
rect 30092 11940 30148 11942
rect 29852 10906 29908 10908
rect 29932 10906 29988 10908
rect 30012 10906 30068 10908
rect 30092 10906 30148 10908
rect 29852 10854 29878 10906
rect 29878 10854 29908 10906
rect 29932 10854 29942 10906
rect 29942 10854 29988 10906
rect 30012 10854 30058 10906
rect 30058 10854 30068 10906
rect 30092 10854 30122 10906
rect 30122 10854 30148 10906
rect 29852 10852 29908 10854
rect 29932 10852 29988 10854
rect 30012 10852 30068 10854
rect 30092 10852 30148 10854
rect 29852 9818 29908 9820
rect 29932 9818 29988 9820
rect 30012 9818 30068 9820
rect 30092 9818 30148 9820
rect 29852 9766 29878 9818
rect 29878 9766 29908 9818
rect 29932 9766 29942 9818
rect 29942 9766 29988 9818
rect 30012 9766 30058 9818
rect 30058 9766 30068 9818
rect 30092 9766 30122 9818
rect 30122 9766 30148 9818
rect 29852 9764 29908 9766
rect 29932 9764 29988 9766
rect 30012 9764 30068 9766
rect 30092 9764 30148 9766
rect 29852 8730 29908 8732
rect 29932 8730 29988 8732
rect 30012 8730 30068 8732
rect 30092 8730 30148 8732
rect 29852 8678 29878 8730
rect 29878 8678 29908 8730
rect 29932 8678 29942 8730
rect 29942 8678 29988 8730
rect 30012 8678 30058 8730
rect 30058 8678 30068 8730
rect 30092 8678 30122 8730
rect 30122 8678 30148 8730
rect 29852 8676 29908 8678
rect 29932 8676 29988 8678
rect 30012 8676 30068 8678
rect 30092 8676 30148 8678
rect 29852 7642 29908 7644
rect 29932 7642 29988 7644
rect 30012 7642 30068 7644
rect 30092 7642 30148 7644
rect 29852 7590 29878 7642
rect 29878 7590 29908 7642
rect 29932 7590 29942 7642
rect 29942 7590 29988 7642
rect 30012 7590 30058 7642
rect 30058 7590 30068 7642
rect 30092 7590 30122 7642
rect 30122 7590 30148 7642
rect 29852 7588 29908 7590
rect 29932 7588 29988 7590
rect 30012 7588 30068 7590
rect 30092 7588 30148 7590
rect 29852 6554 29908 6556
rect 29932 6554 29988 6556
rect 30012 6554 30068 6556
rect 30092 6554 30148 6556
rect 29852 6502 29878 6554
rect 29878 6502 29908 6554
rect 29932 6502 29942 6554
rect 29942 6502 29988 6554
rect 30012 6502 30058 6554
rect 30058 6502 30068 6554
rect 30092 6502 30122 6554
rect 30122 6502 30148 6554
rect 29852 6500 29908 6502
rect 29932 6500 29988 6502
rect 30012 6500 30068 6502
rect 30092 6500 30148 6502
rect 29852 5466 29908 5468
rect 29932 5466 29988 5468
rect 30012 5466 30068 5468
rect 30092 5466 30148 5468
rect 29852 5414 29878 5466
rect 29878 5414 29908 5466
rect 29932 5414 29942 5466
rect 29942 5414 29988 5466
rect 30012 5414 30058 5466
rect 30058 5414 30068 5466
rect 30092 5414 30122 5466
rect 30122 5414 30148 5466
rect 29852 5412 29908 5414
rect 29932 5412 29988 5414
rect 30012 5412 30068 5414
rect 30092 5412 30148 5414
rect 29852 4378 29908 4380
rect 29932 4378 29988 4380
rect 30012 4378 30068 4380
rect 30092 4378 30148 4380
rect 29852 4326 29878 4378
rect 29878 4326 29908 4378
rect 29932 4326 29942 4378
rect 29942 4326 29988 4378
rect 30012 4326 30058 4378
rect 30058 4326 30068 4378
rect 30092 4326 30122 4378
rect 30122 4326 30148 4378
rect 29852 4324 29908 4326
rect 29932 4324 29988 4326
rect 30012 4324 30068 4326
rect 30092 4324 30148 4326
rect 29852 3290 29908 3292
rect 29932 3290 29988 3292
rect 30012 3290 30068 3292
rect 30092 3290 30148 3292
rect 29852 3238 29878 3290
rect 29878 3238 29908 3290
rect 29932 3238 29942 3290
rect 29942 3238 29988 3290
rect 30012 3238 30058 3290
rect 30058 3238 30068 3290
rect 30092 3238 30122 3290
rect 30122 3238 30148 3290
rect 29852 3236 29908 3238
rect 29932 3236 29988 3238
rect 30012 3236 30068 3238
rect 30092 3236 30148 3238
rect 29852 2202 29908 2204
rect 29932 2202 29988 2204
rect 30012 2202 30068 2204
rect 30092 2202 30148 2204
rect 29852 2150 29878 2202
rect 29878 2150 29908 2202
rect 29932 2150 29942 2202
rect 29942 2150 29988 2202
rect 30012 2150 30058 2202
rect 30058 2150 30068 2202
rect 30092 2150 30122 2202
rect 30122 2150 30148 2202
rect 29852 2148 29908 2150
rect 29932 2148 29988 2150
rect 30012 2148 30068 2150
rect 30092 2148 30148 2150
rect 34518 26424 34574 26480
rect 35714 26560 35770 26616
rect 39484 27770 39540 27772
rect 39564 27770 39620 27772
rect 39644 27770 39700 27772
rect 39724 27770 39780 27772
rect 39484 27718 39510 27770
rect 39510 27718 39540 27770
rect 39564 27718 39574 27770
rect 39574 27718 39620 27770
rect 39644 27718 39690 27770
rect 39690 27718 39700 27770
rect 39724 27718 39754 27770
rect 39754 27718 39780 27770
rect 39484 27716 39540 27718
rect 39564 27716 39620 27718
rect 39644 27716 39700 27718
rect 39724 27716 39780 27718
rect 39026 27396 39082 27432
rect 39026 27376 39028 27396
rect 39028 27376 39080 27396
rect 39080 27376 39082 27396
rect 39484 26682 39540 26684
rect 39564 26682 39620 26684
rect 39644 26682 39700 26684
rect 39724 26682 39780 26684
rect 39484 26630 39510 26682
rect 39510 26630 39540 26682
rect 39564 26630 39574 26682
rect 39574 26630 39620 26682
rect 39644 26630 39690 26682
rect 39690 26630 39700 26682
rect 39724 26630 39754 26682
rect 39754 26630 39780 26682
rect 39484 26628 39540 26630
rect 39564 26628 39620 26630
rect 39644 26628 39700 26630
rect 39724 26628 39780 26630
rect 39484 25594 39540 25596
rect 39564 25594 39620 25596
rect 39644 25594 39700 25596
rect 39724 25594 39780 25596
rect 39484 25542 39510 25594
rect 39510 25542 39540 25594
rect 39564 25542 39574 25594
rect 39574 25542 39620 25594
rect 39644 25542 39690 25594
rect 39690 25542 39700 25594
rect 39724 25542 39754 25594
rect 39754 25542 39780 25594
rect 39484 25540 39540 25542
rect 39564 25540 39620 25542
rect 39644 25540 39700 25542
rect 39724 25540 39780 25542
rect 39484 24506 39540 24508
rect 39564 24506 39620 24508
rect 39644 24506 39700 24508
rect 39724 24506 39780 24508
rect 39484 24454 39510 24506
rect 39510 24454 39540 24506
rect 39564 24454 39574 24506
rect 39574 24454 39620 24506
rect 39644 24454 39690 24506
rect 39690 24454 39700 24506
rect 39724 24454 39754 24506
rect 39754 24454 39780 24506
rect 39484 24452 39540 24454
rect 39564 24452 39620 24454
rect 39644 24452 39700 24454
rect 39724 24452 39780 24454
rect 39484 23418 39540 23420
rect 39564 23418 39620 23420
rect 39644 23418 39700 23420
rect 39724 23418 39780 23420
rect 39484 23366 39510 23418
rect 39510 23366 39540 23418
rect 39564 23366 39574 23418
rect 39574 23366 39620 23418
rect 39644 23366 39690 23418
rect 39690 23366 39700 23418
rect 39724 23366 39754 23418
rect 39754 23366 39780 23418
rect 39484 23364 39540 23366
rect 39564 23364 39620 23366
rect 39644 23364 39700 23366
rect 39724 23364 39780 23366
rect 39484 22330 39540 22332
rect 39564 22330 39620 22332
rect 39644 22330 39700 22332
rect 39724 22330 39780 22332
rect 39484 22278 39510 22330
rect 39510 22278 39540 22330
rect 39564 22278 39574 22330
rect 39574 22278 39620 22330
rect 39644 22278 39690 22330
rect 39690 22278 39700 22330
rect 39724 22278 39754 22330
rect 39754 22278 39780 22330
rect 39484 22276 39540 22278
rect 39564 22276 39620 22278
rect 39644 22276 39700 22278
rect 39724 22276 39780 22278
rect 39484 21242 39540 21244
rect 39564 21242 39620 21244
rect 39644 21242 39700 21244
rect 39724 21242 39780 21244
rect 39484 21190 39510 21242
rect 39510 21190 39540 21242
rect 39564 21190 39574 21242
rect 39574 21190 39620 21242
rect 39644 21190 39690 21242
rect 39690 21190 39700 21242
rect 39724 21190 39754 21242
rect 39754 21190 39780 21242
rect 39484 21188 39540 21190
rect 39564 21188 39620 21190
rect 39644 21188 39700 21190
rect 39724 21188 39780 21190
rect 39484 20154 39540 20156
rect 39564 20154 39620 20156
rect 39644 20154 39700 20156
rect 39724 20154 39780 20156
rect 39484 20102 39510 20154
rect 39510 20102 39540 20154
rect 39564 20102 39574 20154
rect 39574 20102 39620 20154
rect 39644 20102 39690 20154
rect 39690 20102 39700 20154
rect 39724 20102 39754 20154
rect 39754 20102 39780 20154
rect 39484 20100 39540 20102
rect 39564 20100 39620 20102
rect 39644 20100 39700 20102
rect 39724 20100 39780 20102
rect 39484 19066 39540 19068
rect 39564 19066 39620 19068
rect 39644 19066 39700 19068
rect 39724 19066 39780 19068
rect 39484 19014 39510 19066
rect 39510 19014 39540 19066
rect 39564 19014 39574 19066
rect 39574 19014 39620 19066
rect 39644 19014 39690 19066
rect 39690 19014 39700 19066
rect 39724 19014 39754 19066
rect 39754 19014 39780 19066
rect 39484 19012 39540 19014
rect 39564 19012 39620 19014
rect 39644 19012 39700 19014
rect 39724 19012 39780 19014
rect 39484 17978 39540 17980
rect 39564 17978 39620 17980
rect 39644 17978 39700 17980
rect 39724 17978 39780 17980
rect 39484 17926 39510 17978
rect 39510 17926 39540 17978
rect 39564 17926 39574 17978
rect 39574 17926 39620 17978
rect 39644 17926 39690 17978
rect 39690 17926 39700 17978
rect 39724 17926 39754 17978
rect 39754 17926 39780 17978
rect 39484 17924 39540 17926
rect 39564 17924 39620 17926
rect 39644 17924 39700 17926
rect 39724 17924 39780 17926
rect 39484 16890 39540 16892
rect 39564 16890 39620 16892
rect 39644 16890 39700 16892
rect 39724 16890 39780 16892
rect 39484 16838 39510 16890
rect 39510 16838 39540 16890
rect 39564 16838 39574 16890
rect 39574 16838 39620 16890
rect 39644 16838 39690 16890
rect 39690 16838 39700 16890
rect 39724 16838 39754 16890
rect 39754 16838 39780 16890
rect 39484 16836 39540 16838
rect 39564 16836 39620 16838
rect 39644 16836 39700 16838
rect 39724 16836 39780 16838
rect 39484 15802 39540 15804
rect 39564 15802 39620 15804
rect 39644 15802 39700 15804
rect 39724 15802 39780 15804
rect 39484 15750 39510 15802
rect 39510 15750 39540 15802
rect 39564 15750 39574 15802
rect 39574 15750 39620 15802
rect 39644 15750 39690 15802
rect 39690 15750 39700 15802
rect 39724 15750 39754 15802
rect 39754 15750 39780 15802
rect 39484 15748 39540 15750
rect 39564 15748 39620 15750
rect 39644 15748 39700 15750
rect 39724 15748 39780 15750
rect 39484 14714 39540 14716
rect 39564 14714 39620 14716
rect 39644 14714 39700 14716
rect 39724 14714 39780 14716
rect 39484 14662 39510 14714
rect 39510 14662 39540 14714
rect 39564 14662 39574 14714
rect 39574 14662 39620 14714
rect 39644 14662 39690 14714
rect 39690 14662 39700 14714
rect 39724 14662 39754 14714
rect 39754 14662 39780 14714
rect 39484 14660 39540 14662
rect 39564 14660 39620 14662
rect 39644 14660 39700 14662
rect 39724 14660 39780 14662
rect 39484 13626 39540 13628
rect 39564 13626 39620 13628
rect 39644 13626 39700 13628
rect 39724 13626 39780 13628
rect 39484 13574 39510 13626
rect 39510 13574 39540 13626
rect 39564 13574 39574 13626
rect 39574 13574 39620 13626
rect 39644 13574 39690 13626
rect 39690 13574 39700 13626
rect 39724 13574 39754 13626
rect 39754 13574 39780 13626
rect 39484 13572 39540 13574
rect 39564 13572 39620 13574
rect 39644 13572 39700 13574
rect 39724 13572 39780 13574
rect 39484 12538 39540 12540
rect 39564 12538 39620 12540
rect 39644 12538 39700 12540
rect 39724 12538 39780 12540
rect 39484 12486 39510 12538
rect 39510 12486 39540 12538
rect 39564 12486 39574 12538
rect 39574 12486 39620 12538
rect 39644 12486 39690 12538
rect 39690 12486 39700 12538
rect 39724 12486 39754 12538
rect 39754 12486 39780 12538
rect 39484 12484 39540 12486
rect 39564 12484 39620 12486
rect 39644 12484 39700 12486
rect 39724 12484 39780 12486
rect 39484 11450 39540 11452
rect 39564 11450 39620 11452
rect 39644 11450 39700 11452
rect 39724 11450 39780 11452
rect 39484 11398 39510 11450
rect 39510 11398 39540 11450
rect 39564 11398 39574 11450
rect 39574 11398 39620 11450
rect 39644 11398 39690 11450
rect 39690 11398 39700 11450
rect 39724 11398 39754 11450
rect 39754 11398 39780 11450
rect 39484 11396 39540 11398
rect 39564 11396 39620 11398
rect 39644 11396 39700 11398
rect 39724 11396 39780 11398
rect 39484 10362 39540 10364
rect 39564 10362 39620 10364
rect 39644 10362 39700 10364
rect 39724 10362 39780 10364
rect 39484 10310 39510 10362
rect 39510 10310 39540 10362
rect 39564 10310 39574 10362
rect 39574 10310 39620 10362
rect 39644 10310 39690 10362
rect 39690 10310 39700 10362
rect 39724 10310 39754 10362
rect 39754 10310 39780 10362
rect 39484 10308 39540 10310
rect 39564 10308 39620 10310
rect 39644 10308 39700 10310
rect 39724 10308 39780 10310
rect 39484 9274 39540 9276
rect 39564 9274 39620 9276
rect 39644 9274 39700 9276
rect 39724 9274 39780 9276
rect 39484 9222 39510 9274
rect 39510 9222 39540 9274
rect 39564 9222 39574 9274
rect 39574 9222 39620 9274
rect 39644 9222 39690 9274
rect 39690 9222 39700 9274
rect 39724 9222 39754 9274
rect 39754 9222 39780 9274
rect 39484 9220 39540 9222
rect 39564 9220 39620 9222
rect 39644 9220 39700 9222
rect 39724 9220 39780 9222
rect 39484 8186 39540 8188
rect 39564 8186 39620 8188
rect 39644 8186 39700 8188
rect 39724 8186 39780 8188
rect 39484 8134 39510 8186
rect 39510 8134 39540 8186
rect 39564 8134 39574 8186
rect 39574 8134 39620 8186
rect 39644 8134 39690 8186
rect 39690 8134 39700 8186
rect 39724 8134 39754 8186
rect 39754 8134 39780 8186
rect 39484 8132 39540 8134
rect 39564 8132 39620 8134
rect 39644 8132 39700 8134
rect 39724 8132 39780 8134
rect 39484 7098 39540 7100
rect 39564 7098 39620 7100
rect 39644 7098 39700 7100
rect 39724 7098 39780 7100
rect 39484 7046 39510 7098
rect 39510 7046 39540 7098
rect 39564 7046 39574 7098
rect 39574 7046 39620 7098
rect 39644 7046 39690 7098
rect 39690 7046 39700 7098
rect 39724 7046 39754 7098
rect 39754 7046 39780 7098
rect 39484 7044 39540 7046
rect 39564 7044 39620 7046
rect 39644 7044 39700 7046
rect 39724 7044 39780 7046
rect 39484 6010 39540 6012
rect 39564 6010 39620 6012
rect 39644 6010 39700 6012
rect 39724 6010 39780 6012
rect 39484 5958 39510 6010
rect 39510 5958 39540 6010
rect 39564 5958 39574 6010
rect 39574 5958 39620 6010
rect 39644 5958 39690 6010
rect 39690 5958 39700 6010
rect 39724 5958 39754 6010
rect 39754 5958 39780 6010
rect 39484 5956 39540 5958
rect 39564 5956 39620 5958
rect 39644 5956 39700 5958
rect 39724 5956 39780 5958
rect 39484 4922 39540 4924
rect 39564 4922 39620 4924
rect 39644 4922 39700 4924
rect 39724 4922 39780 4924
rect 39484 4870 39510 4922
rect 39510 4870 39540 4922
rect 39564 4870 39574 4922
rect 39574 4870 39620 4922
rect 39644 4870 39690 4922
rect 39690 4870 39700 4922
rect 39724 4870 39754 4922
rect 39754 4870 39780 4922
rect 39484 4868 39540 4870
rect 39564 4868 39620 4870
rect 39644 4868 39700 4870
rect 39724 4868 39780 4870
rect 39484 3834 39540 3836
rect 39564 3834 39620 3836
rect 39644 3834 39700 3836
rect 39724 3834 39780 3836
rect 39484 3782 39510 3834
rect 39510 3782 39540 3834
rect 39564 3782 39574 3834
rect 39574 3782 39620 3834
rect 39644 3782 39690 3834
rect 39690 3782 39700 3834
rect 39724 3782 39754 3834
rect 39754 3782 39780 3834
rect 39484 3780 39540 3782
rect 39564 3780 39620 3782
rect 39644 3780 39700 3782
rect 39724 3780 39780 3782
rect 39484 2746 39540 2748
rect 39564 2746 39620 2748
rect 39644 2746 39700 2748
rect 39724 2746 39780 2748
rect 39484 2694 39510 2746
rect 39510 2694 39540 2746
rect 39564 2694 39574 2746
rect 39574 2694 39620 2746
rect 39644 2694 39690 2746
rect 39690 2694 39700 2746
rect 39724 2694 39754 2746
rect 39754 2694 39780 2746
rect 39484 2692 39540 2694
rect 39564 2692 39620 2694
rect 39644 2692 39700 2694
rect 39724 2692 39780 2694
rect 44086 27004 44088 27024
rect 44088 27004 44140 27024
rect 44140 27004 44142 27024
rect 44086 26968 44142 27004
rect 43626 2896 43682 2952
rect 47214 15544 47270 15600
rect 49116 27226 49172 27228
rect 49196 27226 49252 27228
rect 49276 27226 49332 27228
rect 49356 27226 49412 27228
rect 49116 27174 49142 27226
rect 49142 27174 49172 27226
rect 49196 27174 49206 27226
rect 49206 27174 49252 27226
rect 49276 27174 49322 27226
rect 49322 27174 49332 27226
rect 49356 27174 49386 27226
rect 49386 27174 49412 27226
rect 49116 27172 49172 27174
rect 49196 27172 49252 27174
rect 49276 27172 49332 27174
rect 49356 27172 49412 27174
rect 49422 26308 49478 26344
rect 49422 26288 49424 26308
rect 49424 26288 49476 26308
rect 49476 26288 49478 26308
rect 49116 26138 49172 26140
rect 49196 26138 49252 26140
rect 49276 26138 49332 26140
rect 49356 26138 49412 26140
rect 49116 26086 49142 26138
rect 49142 26086 49172 26138
rect 49196 26086 49206 26138
rect 49206 26086 49252 26138
rect 49276 26086 49322 26138
rect 49322 26086 49332 26138
rect 49356 26086 49386 26138
rect 49386 26086 49412 26138
rect 49116 26084 49172 26086
rect 49196 26084 49252 26086
rect 49276 26084 49332 26086
rect 49356 26084 49412 26086
rect 49116 25050 49172 25052
rect 49196 25050 49252 25052
rect 49276 25050 49332 25052
rect 49356 25050 49412 25052
rect 49116 24998 49142 25050
rect 49142 24998 49172 25050
rect 49196 24998 49206 25050
rect 49206 24998 49252 25050
rect 49276 24998 49322 25050
rect 49322 24998 49332 25050
rect 49356 24998 49386 25050
rect 49386 24998 49412 25050
rect 49116 24996 49172 24998
rect 49196 24996 49252 24998
rect 49276 24996 49332 24998
rect 49356 24996 49412 24998
rect 49116 23962 49172 23964
rect 49196 23962 49252 23964
rect 49276 23962 49332 23964
rect 49356 23962 49412 23964
rect 49116 23910 49142 23962
rect 49142 23910 49172 23962
rect 49196 23910 49206 23962
rect 49206 23910 49252 23962
rect 49276 23910 49322 23962
rect 49322 23910 49332 23962
rect 49356 23910 49386 23962
rect 49386 23910 49412 23962
rect 49116 23908 49172 23910
rect 49196 23908 49252 23910
rect 49276 23908 49332 23910
rect 49356 23908 49412 23910
rect 49116 22874 49172 22876
rect 49196 22874 49252 22876
rect 49276 22874 49332 22876
rect 49356 22874 49412 22876
rect 49116 22822 49142 22874
rect 49142 22822 49172 22874
rect 49196 22822 49206 22874
rect 49206 22822 49252 22874
rect 49276 22822 49322 22874
rect 49322 22822 49332 22874
rect 49356 22822 49386 22874
rect 49386 22822 49412 22874
rect 49116 22820 49172 22822
rect 49196 22820 49252 22822
rect 49276 22820 49332 22822
rect 49356 22820 49412 22822
rect 49116 21786 49172 21788
rect 49196 21786 49252 21788
rect 49276 21786 49332 21788
rect 49356 21786 49412 21788
rect 49116 21734 49142 21786
rect 49142 21734 49172 21786
rect 49196 21734 49206 21786
rect 49206 21734 49252 21786
rect 49276 21734 49322 21786
rect 49322 21734 49332 21786
rect 49356 21734 49386 21786
rect 49386 21734 49412 21786
rect 49116 21732 49172 21734
rect 49196 21732 49252 21734
rect 49276 21732 49332 21734
rect 49356 21732 49412 21734
rect 49116 20698 49172 20700
rect 49196 20698 49252 20700
rect 49276 20698 49332 20700
rect 49356 20698 49412 20700
rect 49116 20646 49142 20698
rect 49142 20646 49172 20698
rect 49196 20646 49206 20698
rect 49206 20646 49252 20698
rect 49276 20646 49322 20698
rect 49322 20646 49332 20698
rect 49356 20646 49386 20698
rect 49386 20646 49412 20698
rect 49116 20644 49172 20646
rect 49196 20644 49252 20646
rect 49276 20644 49332 20646
rect 49356 20644 49412 20646
rect 49116 19610 49172 19612
rect 49196 19610 49252 19612
rect 49276 19610 49332 19612
rect 49356 19610 49412 19612
rect 49116 19558 49142 19610
rect 49142 19558 49172 19610
rect 49196 19558 49206 19610
rect 49206 19558 49252 19610
rect 49276 19558 49322 19610
rect 49322 19558 49332 19610
rect 49356 19558 49386 19610
rect 49386 19558 49412 19610
rect 49116 19556 49172 19558
rect 49196 19556 49252 19558
rect 49276 19556 49332 19558
rect 49356 19556 49412 19558
rect 49116 18522 49172 18524
rect 49196 18522 49252 18524
rect 49276 18522 49332 18524
rect 49356 18522 49412 18524
rect 49116 18470 49142 18522
rect 49142 18470 49172 18522
rect 49196 18470 49206 18522
rect 49206 18470 49252 18522
rect 49276 18470 49322 18522
rect 49322 18470 49332 18522
rect 49356 18470 49386 18522
rect 49386 18470 49412 18522
rect 49116 18468 49172 18470
rect 49196 18468 49252 18470
rect 49276 18468 49332 18470
rect 49356 18468 49412 18470
rect 49116 17434 49172 17436
rect 49196 17434 49252 17436
rect 49276 17434 49332 17436
rect 49356 17434 49412 17436
rect 49116 17382 49142 17434
rect 49142 17382 49172 17434
rect 49196 17382 49206 17434
rect 49206 17382 49252 17434
rect 49276 17382 49322 17434
rect 49322 17382 49332 17434
rect 49356 17382 49386 17434
rect 49386 17382 49412 17434
rect 49116 17380 49172 17382
rect 49196 17380 49252 17382
rect 49276 17380 49332 17382
rect 49356 17380 49412 17382
rect 49116 16346 49172 16348
rect 49196 16346 49252 16348
rect 49276 16346 49332 16348
rect 49356 16346 49412 16348
rect 49116 16294 49142 16346
rect 49142 16294 49172 16346
rect 49196 16294 49206 16346
rect 49206 16294 49252 16346
rect 49276 16294 49322 16346
rect 49322 16294 49332 16346
rect 49356 16294 49386 16346
rect 49386 16294 49412 16346
rect 49116 16292 49172 16294
rect 49196 16292 49252 16294
rect 49276 16292 49332 16294
rect 49356 16292 49412 16294
rect 49116 15258 49172 15260
rect 49196 15258 49252 15260
rect 49276 15258 49332 15260
rect 49356 15258 49412 15260
rect 49116 15206 49142 15258
rect 49142 15206 49172 15258
rect 49196 15206 49206 15258
rect 49206 15206 49252 15258
rect 49276 15206 49322 15258
rect 49322 15206 49332 15258
rect 49356 15206 49386 15258
rect 49386 15206 49412 15258
rect 49116 15204 49172 15206
rect 49196 15204 49252 15206
rect 49276 15204 49332 15206
rect 49356 15204 49412 15206
rect 49116 14170 49172 14172
rect 49196 14170 49252 14172
rect 49276 14170 49332 14172
rect 49356 14170 49412 14172
rect 49116 14118 49142 14170
rect 49142 14118 49172 14170
rect 49196 14118 49206 14170
rect 49206 14118 49252 14170
rect 49276 14118 49322 14170
rect 49322 14118 49332 14170
rect 49356 14118 49386 14170
rect 49386 14118 49412 14170
rect 49116 14116 49172 14118
rect 49196 14116 49252 14118
rect 49276 14116 49332 14118
rect 49356 14116 49412 14118
rect 49116 13082 49172 13084
rect 49196 13082 49252 13084
rect 49276 13082 49332 13084
rect 49356 13082 49412 13084
rect 49116 13030 49142 13082
rect 49142 13030 49172 13082
rect 49196 13030 49206 13082
rect 49206 13030 49252 13082
rect 49276 13030 49322 13082
rect 49322 13030 49332 13082
rect 49356 13030 49386 13082
rect 49386 13030 49412 13082
rect 49116 13028 49172 13030
rect 49196 13028 49252 13030
rect 49276 13028 49332 13030
rect 49356 13028 49412 13030
rect 49116 11994 49172 11996
rect 49196 11994 49252 11996
rect 49276 11994 49332 11996
rect 49356 11994 49412 11996
rect 49116 11942 49142 11994
rect 49142 11942 49172 11994
rect 49196 11942 49206 11994
rect 49206 11942 49252 11994
rect 49276 11942 49322 11994
rect 49322 11942 49332 11994
rect 49356 11942 49386 11994
rect 49386 11942 49412 11994
rect 49116 11940 49172 11942
rect 49196 11940 49252 11942
rect 49276 11940 49332 11942
rect 49356 11940 49412 11942
rect 49116 10906 49172 10908
rect 49196 10906 49252 10908
rect 49276 10906 49332 10908
rect 49356 10906 49412 10908
rect 49116 10854 49142 10906
rect 49142 10854 49172 10906
rect 49196 10854 49206 10906
rect 49206 10854 49252 10906
rect 49276 10854 49322 10906
rect 49322 10854 49332 10906
rect 49356 10854 49386 10906
rect 49386 10854 49412 10906
rect 49116 10852 49172 10854
rect 49196 10852 49252 10854
rect 49276 10852 49332 10854
rect 49356 10852 49412 10854
rect 49116 9818 49172 9820
rect 49196 9818 49252 9820
rect 49276 9818 49332 9820
rect 49356 9818 49412 9820
rect 49116 9766 49142 9818
rect 49142 9766 49172 9818
rect 49196 9766 49206 9818
rect 49206 9766 49252 9818
rect 49276 9766 49322 9818
rect 49322 9766 49332 9818
rect 49356 9766 49386 9818
rect 49386 9766 49412 9818
rect 49116 9764 49172 9766
rect 49196 9764 49252 9766
rect 49276 9764 49332 9766
rect 49356 9764 49412 9766
rect 49116 8730 49172 8732
rect 49196 8730 49252 8732
rect 49276 8730 49332 8732
rect 49356 8730 49412 8732
rect 49116 8678 49142 8730
rect 49142 8678 49172 8730
rect 49196 8678 49206 8730
rect 49206 8678 49252 8730
rect 49276 8678 49322 8730
rect 49322 8678 49332 8730
rect 49356 8678 49386 8730
rect 49386 8678 49412 8730
rect 49116 8676 49172 8678
rect 49196 8676 49252 8678
rect 49276 8676 49332 8678
rect 49356 8676 49412 8678
rect 49116 7642 49172 7644
rect 49196 7642 49252 7644
rect 49276 7642 49332 7644
rect 49356 7642 49412 7644
rect 49116 7590 49142 7642
rect 49142 7590 49172 7642
rect 49196 7590 49206 7642
rect 49206 7590 49252 7642
rect 49276 7590 49322 7642
rect 49322 7590 49332 7642
rect 49356 7590 49386 7642
rect 49386 7590 49412 7642
rect 49116 7588 49172 7590
rect 49196 7588 49252 7590
rect 49276 7588 49332 7590
rect 49356 7588 49412 7590
rect 49116 6554 49172 6556
rect 49196 6554 49252 6556
rect 49276 6554 49332 6556
rect 49356 6554 49412 6556
rect 49116 6502 49142 6554
rect 49142 6502 49172 6554
rect 49196 6502 49206 6554
rect 49206 6502 49252 6554
rect 49276 6502 49322 6554
rect 49322 6502 49332 6554
rect 49356 6502 49386 6554
rect 49386 6502 49412 6554
rect 49116 6500 49172 6502
rect 49196 6500 49252 6502
rect 49276 6500 49332 6502
rect 49356 6500 49412 6502
rect 49116 5466 49172 5468
rect 49196 5466 49252 5468
rect 49276 5466 49332 5468
rect 49356 5466 49412 5468
rect 49116 5414 49142 5466
rect 49142 5414 49172 5466
rect 49196 5414 49206 5466
rect 49206 5414 49252 5466
rect 49276 5414 49322 5466
rect 49322 5414 49332 5466
rect 49356 5414 49386 5466
rect 49386 5414 49412 5466
rect 49116 5412 49172 5414
rect 49196 5412 49252 5414
rect 49276 5412 49332 5414
rect 49356 5412 49412 5414
rect 49116 4378 49172 4380
rect 49196 4378 49252 4380
rect 49276 4378 49332 4380
rect 49356 4378 49412 4380
rect 49116 4326 49142 4378
rect 49142 4326 49172 4378
rect 49196 4326 49206 4378
rect 49206 4326 49252 4378
rect 49276 4326 49322 4378
rect 49322 4326 49332 4378
rect 49356 4326 49386 4378
rect 49386 4326 49412 4378
rect 49116 4324 49172 4326
rect 49196 4324 49252 4326
rect 49276 4324 49332 4326
rect 49356 4324 49412 4326
rect 49116 3290 49172 3292
rect 49196 3290 49252 3292
rect 49276 3290 49332 3292
rect 49356 3290 49412 3292
rect 49116 3238 49142 3290
rect 49142 3238 49172 3290
rect 49196 3238 49206 3290
rect 49206 3238 49252 3290
rect 49276 3238 49322 3290
rect 49322 3238 49332 3290
rect 49356 3238 49386 3290
rect 49386 3238 49412 3290
rect 49116 3236 49172 3238
rect 49196 3236 49252 3238
rect 49276 3236 49332 3238
rect 49356 3236 49412 3238
rect 49698 3068 49700 3088
rect 49700 3068 49752 3088
rect 49752 3068 49754 3088
rect 49698 3032 49754 3068
rect 49116 2202 49172 2204
rect 49196 2202 49252 2204
rect 49276 2202 49332 2204
rect 49356 2202 49412 2204
rect 49116 2150 49142 2202
rect 49142 2150 49172 2202
rect 49196 2150 49206 2202
rect 49206 2150 49252 2202
rect 49276 2150 49322 2202
rect 49322 2150 49332 2202
rect 49356 2150 49386 2202
rect 49386 2150 49412 2202
rect 49116 2148 49172 2150
rect 49196 2148 49252 2150
rect 49276 2148 49332 2150
rect 49356 2148 49412 2150
rect 54390 26868 54392 26888
rect 54392 26868 54444 26888
rect 54444 26868 54446 26888
rect 54390 26832 54446 26868
rect 55126 26460 55128 26480
rect 55128 26460 55180 26480
rect 55180 26460 55182 26480
rect 55126 26424 55182 26460
rect 58162 28600 58218 28656
rect 57242 25880 57298 25936
rect 56414 2080 56470 2136
rect 57886 26560 57942 26616
rect 58070 27240 58126 27296
rect 57886 24520 57942 24576
rect 57886 21800 57942 21856
rect 58162 23840 58218 23896
rect 58162 22516 58164 22536
rect 58164 22516 58216 22536
rect 58216 22516 58218 22536
rect 58162 22480 58218 22516
rect 58162 21120 58218 21176
rect 58162 19780 58218 19816
rect 58162 19760 58164 19780
rect 58164 19760 58216 19780
rect 58216 19760 58218 19780
rect 58162 19080 58218 19136
rect 58162 17740 58218 17776
rect 58162 17720 58164 17740
rect 58164 17720 58216 17740
rect 58216 17720 58218 17740
rect 58070 17060 58126 17096
rect 58070 17040 58072 17060
rect 58072 17040 58124 17060
rect 58124 17040 58126 17060
rect 57886 12960 57942 13016
rect 58162 16360 58218 16416
rect 58162 15000 58218 15056
rect 58162 14320 58218 14376
rect 58162 12300 58218 12336
rect 58162 12280 58164 12300
rect 58164 12280 58216 12300
rect 58216 12280 58218 12300
rect 58162 11620 58218 11656
rect 58162 11600 58164 11620
rect 58164 11600 58216 11620
rect 58216 11600 58218 11620
rect 58162 10240 58218 10296
rect 58162 9580 58218 9616
rect 58162 9560 58164 9580
rect 58164 9560 58216 9580
rect 58216 9560 58218 9580
rect 58162 8200 58218 8256
rect 58162 7520 58218 7576
rect 58070 6860 58126 6896
rect 58070 6840 58072 6860
rect 58072 6840 58124 6860
rect 58124 6840 58126 6860
rect 58162 5480 58218 5536
rect 58070 4800 58126 4856
rect 57794 4120 57850 4176
rect 57886 2760 57942 2816
rect 57702 2352 57758 2408
rect 57610 720 57666 776
<< metal3 >>
rect 0 28658 800 28688
rect 2589 28658 2655 28661
rect 0 28656 2655 28658
rect 0 28600 2594 28656
rect 2650 28600 2655 28656
rect 0 28598 2655 28600
rect 0 28568 800 28598
rect 2589 28595 2655 28598
rect 58157 28658 58223 28661
rect 59200 28658 60000 28688
rect 58157 28656 60000 28658
rect 58157 28600 58162 28656
rect 58218 28600 60000 28656
rect 58157 28598 60000 28600
rect 58157 28595 58223 28598
rect 59200 28568 60000 28598
rect 0 27978 800 28008
rect 2865 27978 2931 27981
rect 0 27976 2931 27978
rect 0 27920 2870 27976
rect 2926 27920 2931 27976
rect 0 27918 2931 27920
rect 0 27888 800 27918
rect 2865 27915 2931 27918
rect 20208 27776 20528 27777
rect 20208 27712 20216 27776
rect 20280 27712 20296 27776
rect 20360 27712 20376 27776
rect 20440 27712 20456 27776
rect 20520 27712 20528 27776
rect 20208 27711 20528 27712
rect 39472 27776 39792 27777
rect 39472 27712 39480 27776
rect 39544 27712 39560 27776
rect 39624 27712 39640 27776
rect 39704 27712 39720 27776
rect 39784 27712 39792 27776
rect 39472 27711 39792 27712
rect 1577 27434 1643 27437
rect 39021 27434 39087 27437
rect 1577 27432 39087 27434
rect 1577 27376 1582 27432
rect 1638 27376 39026 27432
rect 39082 27376 39087 27432
rect 1577 27374 39087 27376
rect 1577 27371 1643 27374
rect 39021 27371 39087 27374
rect 0 27298 800 27328
rect 1485 27298 1551 27301
rect 0 27296 1551 27298
rect 0 27240 1490 27296
rect 1546 27240 1551 27296
rect 0 27238 1551 27240
rect 0 27208 800 27238
rect 1485 27235 1551 27238
rect 58065 27298 58131 27301
rect 59200 27298 60000 27328
rect 58065 27296 60000 27298
rect 58065 27240 58070 27296
rect 58126 27240 60000 27296
rect 58065 27238 60000 27240
rect 58065 27235 58131 27238
rect 10576 27232 10896 27233
rect 10576 27168 10584 27232
rect 10648 27168 10664 27232
rect 10728 27168 10744 27232
rect 10808 27168 10824 27232
rect 10888 27168 10896 27232
rect 10576 27167 10896 27168
rect 29840 27232 30160 27233
rect 29840 27168 29848 27232
rect 29912 27168 29928 27232
rect 29992 27168 30008 27232
rect 30072 27168 30088 27232
rect 30152 27168 30160 27232
rect 29840 27167 30160 27168
rect 49104 27232 49424 27233
rect 49104 27168 49112 27232
rect 49176 27168 49192 27232
rect 49256 27168 49272 27232
rect 49336 27168 49352 27232
rect 49416 27168 49424 27232
rect 59200 27208 60000 27238
rect 49104 27167 49424 27168
rect 11053 27026 11119 27029
rect 44081 27026 44147 27029
rect 11053 27024 44147 27026
rect 11053 26968 11058 27024
rect 11114 26968 44086 27024
rect 44142 26968 44147 27024
rect 11053 26966 44147 26968
rect 11053 26963 11119 26966
rect 44081 26963 44147 26966
rect 20989 26890 21055 26893
rect 54385 26890 54451 26893
rect 20989 26888 54451 26890
rect 20989 26832 20994 26888
rect 21050 26832 54390 26888
rect 54446 26832 54451 26888
rect 20989 26830 54451 26832
rect 20989 26827 21055 26830
rect 54385 26827 54451 26830
rect 20208 26688 20528 26689
rect 20208 26624 20216 26688
rect 20280 26624 20296 26688
rect 20360 26624 20376 26688
rect 20440 26624 20456 26688
rect 20520 26624 20528 26688
rect 20208 26623 20528 26624
rect 39472 26688 39792 26689
rect 39472 26624 39480 26688
rect 39544 26624 39560 26688
rect 39624 26624 39640 26688
rect 39704 26624 39720 26688
rect 39784 26624 39792 26688
rect 39472 26623 39792 26624
rect 27981 26618 28047 26621
rect 35709 26618 35775 26621
rect 27981 26616 35775 26618
rect 27981 26560 27986 26616
rect 28042 26560 35714 26616
rect 35770 26560 35775 26616
rect 27981 26558 35775 26560
rect 27981 26555 28047 26558
rect 35709 26555 35775 26558
rect 57881 26618 57947 26621
rect 59200 26618 60000 26648
rect 57881 26616 60000 26618
rect 57881 26560 57886 26616
rect 57942 26560 60000 26616
rect 57881 26558 60000 26560
rect 57881 26555 57947 26558
rect 59200 26528 60000 26558
rect 3325 26482 3391 26485
rect 29545 26482 29611 26485
rect 3325 26480 29611 26482
rect 3325 26424 3330 26480
rect 3386 26424 29550 26480
rect 29606 26424 29611 26480
rect 3325 26422 29611 26424
rect 3325 26419 3391 26422
rect 29545 26419 29611 26422
rect 34513 26482 34579 26485
rect 55121 26482 55187 26485
rect 34513 26480 55187 26482
rect 34513 26424 34518 26480
rect 34574 26424 55126 26480
rect 55182 26424 55187 26480
rect 34513 26422 55187 26424
rect 34513 26419 34579 26422
rect 55121 26419 55187 26422
rect 12893 26346 12959 26349
rect 21081 26346 21147 26349
rect 12893 26344 21147 26346
rect 12893 26288 12898 26344
rect 12954 26288 21086 26344
rect 21142 26288 21147 26344
rect 12893 26286 21147 26288
rect 12893 26283 12959 26286
rect 21081 26283 21147 26286
rect 28165 26346 28231 26349
rect 49417 26346 49483 26349
rect 28165 26344 49483 26346
rect 28165 26288 28170 26344
rect 28226 26288 49422 26344
rect 49478 26288 49483 26344
rect 28165 26286 49483 26288
rect 28165 26283 28231 26286
rect 49417 26283 49483 26286
rect 14181 26210 14247 26213
rect 24485 26210 24551 26213
rect 14181 26208 24551 26210
rect 14181 26152 14186 26208
rect 14242 26152 24490 26208
rect 24546 26152 24551 26208
rect 14181 26150 24551 26152
rect 14181 26147 14247 26150
rect 24485 26147 24551 26150
rect 10576 26144 10896 26145
rect 10576 26080 10584 26144
rect 10648 26080 10664 26144
rect 10728 26080 10744 26144
rect 10808 26080 10824 26144
rect 10888 26080 10896 26144
rect 10576 26079 10896 26080
rect 29840 26144 30160 26145
rect 29840 26080 29848 26144
rect 29912 26080 29928 26144
rect 29992 26080 30008 26144
rect 30072 26080 30088 26144
rect 30152 26080 30160 26144
rect 29840 26079 30160 26080
rect 49104 26144 49424 26145
rect 49104 26080 49112 26144
rect 49176 26080 49192 26144
rect 49256 26080 49272 26144
rect 49336 26080 49352 26144
rect 49416 26080 49424 26144
rect 49104 26079 49424 26080
rect 0 25938 800 25968
rect 1393 25938 1459 25941
rect 0 25936 1459 25938
rect 0 25880 1398 25936
rect 1454 25880 1459 25936
rect 0 25878 1459 25880
rect 0 25848 800 25878
rect 1393 25875 1459 25878
rect 57237 25938 57303 25941
rect 59200 25938 60000 25968
rect 57237 25936 60000 25938
rect 57237 25880 57242 25936
rect 57298 25880 60000 25936
rect 57237 25878 60000 25880
rect 57237 25875 57303 25878
rect 59200 25848 60000 25878
rect 20208 25600 20528 25601
rect 20208 25536 20216 25600
rect 20280 25536 20296 25600
rect 20360 25536 20376 25600
rect 20440 25536 20456 25600
rect 20520 25536 20528 25600
rect 20208 25535 20528 25536
rect 39472 25600 39792 25601
rect 39472 25536 39480 25600
rect 39544 25536 39560 25600
rect 39624 25536 39640 25600
rect 39704 25536 39720 25600
rect 39784 25536 39792 25600
rect 39472 25535 39792 25536
rect 0 25258 800 25288
rect 1393 25258 1459 25261
rect 0 25256 1459 25258
rect 0 25200 1398 25256
rect 1454 25200 1459 25256
rect 0 25198 1459 25200
rect 0 25168 800 25198
rect 1393 25195 1459 25198
rect 10576 25056 10896 25057
rect 10576 24992 10584 25056
rect 10648 24992 10664 25056
rect 10728 24992 10744 25056
rect 10808 24992 10824 25056
rect 10888 24992 10896 25056
rect 10576 24991 10896 24992
rect 29840 25056 30160 25057
rect 29840 24992 29848 25056
rect 29912 24992 29928 25056
rect 29992 24992 30008 25056
rect 30072 24992 30088 25056
rect 30152 24992 30160 25056
rect 29840 24991 30160 24992
rect 49104 25056 49424 25057
rect 49104 24992 49112 25056
rect 49176 24992 49192 25056
rect 49256 24992 49272 25056
rect 49336 24992 49352 25056
rect 49416 24992 49424 25056
rect 49104 24991 49424 24992
rect 57881 24578 57947 24581
rect 59200 24578 60000 24608
rect 57881 24576 60000 24578
rect 57881 24520 57886 24576
rect 57942 24520 60000 24576
rect 57881 24518 60000 24520
rect 57881 24515 57947 24518
rect 20208 24512 20528 24513
rect 20208 24448 20216 24512
rect 20280 24448 20296 24512
rect 20360 24448 20376 24512
rect 20440 24448 20456 24512
rect 20520 24448 20528 24512
rect 20208 24447 20528 24448
rect 39472 24512 39792 24513
rect 39472 24448 39480 24512
rect 39544 24448 39560 24512
rect 39624 24448 39640 24512
rect 39704 24448 39720 24512
rect 39784 24448 39792 24512
rect 59200 24488 60000 24518
rect 39472 24447 39792 24448
rect 10576 23968 10896 23969
rect 0 23898 800 23928
rect 10576 23904 10584 23968
rect 10648 23904 10664 23968
rect 10728 23904 10744 23968
rect 10808 23904 10824 23968
rect 10888 23904 10896 23968
rect 10576 23903 10896 23904
rect 29840 23968 30160 23969
rect 29840 23904 29848 23968
rect 29912 23904 29928 23968
rect 29992 23904 30008 23968
rect 30072 23904 30088 23968
rect 30152 23904 30160 23968
rect 29840 23903 30160 23904
rect 49104 23968 49424 23969
rect 49104 23904 49112 23968
rect 49176 23904 49192 23968
rect 49256 23904 49272 23968
rect 49336 23904 49352 23968
rect 49416 23904 49424 23968
rect 49104 23903 49424 23904
rect 1485 23898 1551 23901
rect 0 23896 1551 23898
rect 0 23840 1490 23896
rect 1546 23840 1551 23896
rect 0 23838 1551 23840
rect 0 23808 800 23838
rect 1485 23835 1551 23838
rect 58157 23898 58223 23901
rect 59200 23898 60000 23928
rect 58157 23896 60000 23898
rect 58157 23840 58162 23896
rect 58218 23840 60000 23896
rect 58157 23838 60000 23840
rect 58157 23835 58223 23838
rect 59200 23808 60000 23838
rect 20208 23424 20528 23425
rect 20208 23360 20216 23424
rect 20280 23360 20296 23424
rect 20360 23360 20376 23424
rect 20440 23360 20456 23424
rect 20520 23360 20528 23424
rect 20208 23359 20528 23360
rect 39472 23424 39792 23425
rect 39472 23360 39480 23424
rect 39544 23360 39560 23424
rect 39624 23360 39640 23424
rect 39704 23360 39720 23424
rect 39784 23360 39792 23424
rect 39472 23359 39792 23360
rect 0 23218 800 23248
rect 1393 23218 1459 23221
rect 0 23216 1459 23218
rect 0 23160 1398 23216
rect 1454 23160 1459 23216
rect 0 23158 1459 23160
rect 0 23128 800 23158
rect 1393 23155 1459 23158
rect 10576 22880 10896 22881
rect 10576 22816 10584 22880
rect 10648 22816 10664 22880
rect 10728 22816 10744 22880
rect 10808 22816 10824 22880
rect 10888 22816 10896 22880
rect 10576 22815 10896 22816
rect 29840 22880 30160 22881
rect 29840 22816 29848 22880
rect 29912 22816 29928 22880
rect 29992 22816 30008 22880
rect 30072 22816 30088 22880
rect 30152 22816 30160 22880
rect 29840 22815 30160 22816
rect 49104 22880 49424 22881
rect 49104 22816 49112 22880
rect 49176 22816 49192 22880
rect 49256 22816 49272 22880
rect 49336 22816 49352 22880
rect 49416 22816 49424 22880
rect 49104 22815 49424 22816
rect 0 22538 800 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 800 22478
rect 1393 22475 1459 22478
rect 58157 22538 58223 22541
rect 59200 22538 60000 22568
rect 58157 22536 60000 22538
rect 58157 22480 58162 22536
rect 58218 22480 60000 22536
rect 58157 22478 60000 22480
rect 58157 22475 58223 22478
rect 59200 22448 60000 22478
rect 20208 22336 20528 22337
rect 20208 22272 20216 22336
rect 20280 22272 20296 22336
rect 20360 22272 20376 22336
rect 20440 22272 20456 22336
rect 20520 22272 20528 22336
rect 20208 22271 20528 22272
rect 39472 22336 39792 22337
rect 39472 22272 39480 22336
rect 39544 22272 39560 22336
rect 39624 22272 39640 22336
rect 39704 22272 39720 22336
rect 39784 22272 39792 22336
rect 39472 22271 39792 22272
rect 57881 21858 57947 21861
rect 59200 21858 60000 21888
rect 57881 21856 60000 21858
rect 57881 21800 57886 21856
rect 57942 21800 60000 21856
rect 57881 21798 60000 21800
rect 57881 21795 57947 21798
rect 10576 21792 10896 21793
rect 10576 21728 10584 21792
rect 10648 21728 10664 21792
rect 10728 21728 10744 21792
rect 10808 21728 10824 21792
rect 10888 21728 10896 21792
rect 10576 21727 10896 21728
rect 29840 21792 30160 21793
rect 29840 21728 29848 21792
rect 29912 21728 29928 21792
rect 29992 21728 30008 21792
rect 30072 21728 30088 21792
rect 30152 21728 30160 21792
rect 29840 21727 30160 21728
rect 49104 21792 49424 21793
rect 49104 21728 49112 21792
rect 49176 21728 49192 21792
rect 49256 21728 49272 21792
rect 49336 21728 49352 21792
rect 49416 21728 49424 21792
rect 59200 21768 60000 21798
rect 49104 21727 49424 21728
rect 20208 21248 20528 21249
rect 0 21178 800 21208
rect 20208 21184 20216 21248
rect 20280 21184 20296 21248
rect 20360 21184 20376 21248
rect 20440 21184 20456 21248
rect 20520 21184 20528 21248
rect 20208 21183 20528 21184
rect 39472 21248 39792 21249
rect 39472 21184 39480 21248
rect 39544 21184 39560 21248
rect 39624 21184 39640 21248
rect 39704 21184 39720 21248
rect 39784 21184 39792 21248
rect 39472 21183 39792 21184
rect 1485 21178 1551 21181
rect 0 21176 1551 21178
rect 0 21120 1490 21176
rect 1546 21120 1551 21176
rect 0 21118 1551 21120
rect 0 21088 800 21118
rect 1485 21115 1551 21118
rect 58157 21178 58223 21181
rect 59200 21178 60000 21208
rect 58157 21176 60000 21178
rect 58157 21120 58162 21176
rect 58218 21120 60000 21176
rect 58157 21118 60000 21120
rect 58157 21115 58223 21118
rect 59200 21088 60000 21118
rect 10576 20704 10896 20705
rect 10576 20640 10584 20704
rect 10648 20640 10664 20704
rect 10728 20640 10744 20704
rect 10808 20640 10824 20704
rect 10888 20640 10896 20704
rect 10576 20639 10896 20640
rect 29840 20704 30160 20705
rect 29840 20640 29848 20704
rect 29912 20640 29928 20704
rect 29992 20640 30008 20704
rect 30072 20640 30088 20704
rect 30152 20640 30160 20704
rect 29840 20639 30160 20640
rect 49104 20704 49424 20705
rect 49104 20640 49112 20704
rect 49176 20640 49192 20704
rect 49256 20640 49272 20704
rect 49336 20640 49352 20704
rect 49416 20640 49424 20704
rect 49104 20639 49424 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 20208 20160 20528 20161
rect 20208 20096 20216 20160
rect 20280 20096 20296 20160
rect 20360 20096 20376 20160
rect 20440 20096 20456 20160
rect 20520 20096 20528 20160
rect 20208 20095 20528 20096
rect 39472 20160 39792 20161
rect 39472 20096 39480 20160
rect 39544 20096 39560 20160
rect 39624 20096 39640 20160
rect 39704 20096 39720 20160
rect 39784 20096 39792 20160
rect 39472 20095 39792 20096
rect 58157 19818 58223 19821
rect 59200 19818 60000 19848
rect 58157 19816 60000 19818
rect 58157 19760 58162 19816
rect 58218 19760 60000 19816
rect 58157 19758 60000 19760
rect 58157 19755 58223 19758
rect 59200 19728 60000 19758
rect 10576 19616 10896 19617
rect 10576 19552 10584 19616
rect 10648 19552 10664 19616
rect 10728 19552 10744 19616
rect 10808 19552 10824 19616
rect 10888 19552 10896 19616
rect 10576 19551 10896 19552
rect 29840 19616 30160 19617
rect 29840 19552 29848 19616
rect 29912 19552 29928 19616
rect 29992 19552 30008 19616
rect 30072 19552 30088 19616
rect 30152 19552 30160 19616
rect 29840 19551 30160 19552
rect 49104 19616 49424 19617
rect 49104 19552 49112 19616
rect 49176 19552 49192 19616
rect 49256 19552 49272 19616
rect 49336 19552 49352 19616
rect 49416 19552 49424 19616
rect 49104 19551 49424 19552
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 58157 19138 58223 19141
rect 59200 19138 60000 19168
rect 58157 19136 60000 19138
rect 58157 19080 58162 19136
rect 58218 19080 60000 19136
rect 58157 19078 60000 19080
rect 58157 19075 58223 19078
rect 20208 19072 20528 19073
rect 20208 19008 20216 19072
rect 20280 19008 20296 19072
rect 20360 19008 20376 19072
rect 20440 19008 20456 19072
rect 20520 19008 20528 19072
rect 20208 19007 20528 19008
rect 39472 19072 39792 19073
rect 39472 19008 39480 19072
rect 39544 19008 39560 19072
rect 39624 19008 39640 19072
rect 39704 19008 39720 19072
rect 39784 19008 39792 19072
rect 59200 19048 60000 19078
rect 39472 19007 39792 19008
rect 10576 18528 10896 18529
rect 0 18458 800 18488
rect 10576 18464 10584 18528
rect 10648 18464 10664 18528
rect 10728 18464 10744 18528
rect 10808 18464 10824 18528
rect 10888 18464 10896 18528
rect 10576 18463 10896 18464
rect 29840 18528 30160 18529
rect 29840 18464 29848 18528
rect 29912 18464 29928 18528
rect 29992 18464 30008 18528
rect 30072 18464 30088 18528
rect 30152 18464 30160 18528
rect 29840 18463 30160 18464
rect 49104 18528 49424 18529
rect 49104 18464 49112 18528
rect 49176 18464 49192 18528
rect 49256 18464 49272 18528
rect 49336 18464 49352 18528
rect 49416 18464 49424 18528
rect 49104 18463 49424 18464
rect 1393 18458 1459 18461
rect 0 18456 1459 18458
rect 0 18400 1398 18456
rect 1454 18400 1459 18456
rect 0 18398 1459 18400
rect 0 18368 800 18398
rect 1393 18395 1459 18398
rect 20208 17984 20528 17985
rect 20208 17920 20216 17984
rect 20280 17920 20296 17984
rect 20360 17920 20376 17984
rect 20440 17920 20456 17984
rect 20520 17920 20528 17984
rect 20208 17919 20528 17920
rect 39472 17984 39792 17985
rect 39472 17920 39480 17984
rect 39544 17920 39560 17984
rect 39624 17920 39640 17984
rect 39704 17920 39720 17984
rect 39784 17920 39792 17984
rect 39472 17919 39792 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 58157 17778 58223 17781
rect 59200 17778 60000 17808
rect 58157 17776 60000 17778
rect 58157 17720 58162 17776
rect 58218 17720 60000 17776
rect 58157 17718 60000 17720
rect 58157 17715 58223 17718
rect 59200 17688 60000 17718
rect 10576 17440 10896 17441
rect 10576 17376 10584 17440
rect 10648 17376 10664 17440
rect 10728 17376 10744 17440
rect 10808 17376 10824 17440
rect 10888 17376 10896 17440
rect 10576 17375 10896 17376
rect 29840 17440 30160 17441
rect 29840 17376 29848 17440
rect 29912 17376 29928 17440
rect 29992 17376 30008 17440
rect 30072 17376 30088 17440
rect 30152 17376 30160 17440
rect 29840 17375 30160 17376
rect 49104 17440 49424 17441
rect 49104 17376 49112 17440
rect 49176 17376 49192 17440
rect 49256 17376 49272 17440
rect 49336 17376 49352 17440
rect 49416 17376 49424 17440
rect 49104 17375 49424 17376
rect 58065 17098 58131 17101
rect 59200 17098 60000 17128
rect 58065 17096 60000 17098
rect 58065 17040 58070 17096
rect 58126 17040 60000 17096
rect 58065 17038 60000 17040
rect 58065 17035 58131 17038
rect 59200 17008 60000 17038
rect 20208 16896 20528 16897
rect 20208 16832 20216 16896
rect 20280 16832 20296 16896
rect 20360 16832 20376 16896
rect 20440 16832 20456 16896
rect 20520 16832 20528 16896
rect 20208 16831 20528 16832
rect 39472 16896 39792 16897
rect 39472 16832 39480 16896
rect 39544 16832 39560 16896
rect 39624 16832 39640 16896
rect 39704 16832 39720 16896
rect 39784 16832 39792 16896
rect 39472 16831 39792 16832
rect 0 16418 800 16448
rect 1393 16418 1459 16421
rect 0 16416 1459 16418
rect 0 16360 1398 16416
rect 1454 16360 1459 16416
rect 0 16358 1459 16360
rect 0 16328 800 16358
rect 1393 16355 1459 16358
rect 58157 16418 58223 16421
rect 59200 16418 60000 16448
rect 58157 16416 60000 16418
rect 58157 16360 58162 16416
rect 58218 16360 60000 16416
rect 58157 16358 60000 16360
rect 58157 16355 58223 16358
rect 10576 16352 10896 16353
rect 10576 16288 10584 16352
rect 10648 16288 10664 16352
rect 10728 16288 10744 16352
rect 10808 16288 10824 16352
rect 10888 16288 10896 16352
rect 10576 16287 10896 16288
rect 29840 16352 30160 16353
rect 29840 16288 29848 16352
rect 29912 16288 29928 16352
rect 29992 16288 30008 16352
rect 30072 16288 30088 16352
rect 30152 16288 30160 16352
rect 29840 16287 30160 16288
rect 49104 16352 49424 16353
rect 49104 16288 49112 16352
rect 49176 16288 49192 16352
rect 49256 16288 49272 16352
rect 49336 16288 49352 16352
rect 49416 16288 49424 16352
rect 59200 16328 60000 16358
rect 49104 16287 49424 16288
rect 20208 15808 20528 15809
rect 0 15738 800 15768
rect 20208 15744 20216 15808
rect 20280 15744 20296 15808
rect 20360 15744 20376 15808
rect 20440 15744 20456 15808
rect 20520 15744 20528 15808
rect 20208 15743 20528 15744
rect 39472 15808 39792 15809
rect 39472 15744 39480 15808
rect 39544 15744 39560 15808
rect 39624 15744 39640 15808
rect 39704 15744 39720 15808
rect 39784 15744 39792 15808
rect 39472 15743 39792 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 1577 15602 1643 15605
rect 47209 15602 47275 15605
rect 1577 15600 47275 15602
rect 1577 15544 1582 15600
rect 1638 15544 47214 15600
rect 47270 15544 47275 15600
rect 1577 15542 47275 15544
rect 1577 15539 1643 15542
rect 47209 15539 47275 15542
rect 10576 15264 10896 15265
rect 10576 15200 10584 15264
rect 10648 15200 10664 15264
rect 10728 15200 10744 15264
rect 10808 15200 10824 15264
rect 10888 15200 10896 15264
rect 10576 15199 10896 15200
rect 29840 15264 30160 15265
rect 29840 15200 29848 15264
rect 29912 15200 29928 15264
rect 29992 15200 30008 15264
rect 30072 15200 30088 15264
rect 30152 15200 30160 15264
rect 29840 15199 30160 15200
rect 49104 15264 49424 15265
rect 49104 15200 49112 15264
rect 49176 15200 49192 15264
rect 49256 15200 49272 15264
rect 49336 15200 49352 15264
rect 49416 15200 49424 15264
rect 49104 15199 49424 15200
rect 58157 15058 58223 15061
rect 59200 15058 60000 15088
rect 58157 15056 60000 15058
rect 58157 15000 58162 15056
rect 58218 15000 60000 15056
rect 58157 14998 60000 15000
rect 58157 14995 58223 14998
rect 59200 14968 60000 14998
rect 20208 14720 20528 14721
rect 20208 14656 20216 14720
rect 20280 14656 20296 14720
rect 20360 14656 20376 14720
rect 20440 14656 20456 14720
rect 20520 14656 20528 14720
rect 20208 14655 20528 14656
rect 39472 14720 39792 14721
rect 39472 14656 39480 14720
rect 39544 14656 39560 14720
rect 39624 14656 39640 14720
rect 39704 14656 39720 14720
rect 39784 14656 39792 14720
rect 39472 14655 39792 14656
rect 0 14378 800 14408
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14288 800 14318
rect 1393 14315 1459 14318
rect 58157 14378 58223 14381
rect 59200 14378 60000 14408
rect 58157 14376 60000 14378
rect 58157 14320 58162 14376
rect 58218 14320 60000 14376
rect 58157 14318 60000 14320
rect 58157 14315 58223 14318
rect 59200 14288 60000 14318
rect 10576 14176 10896 14177
rect 10576 14112 10584 14176
rect 10648 14112 10664 14176
rect 10728 14112 10744 14176
rect 10808 14112 10824 14176
rect 10888 14112 10896 14176
rect 10576 14111 10896 14112
rect 29840 14176 30160 14177
rect 29840 14112 29848 14176
rect 29912 14112 29928 14176
rect 29992 14112 30008 14176
rect 30072 14112 30088 14176
rect 30152 14112 30160 14176
rect 29840 14111 30160 14112
rect 49104 14176 49424 14177
rect 49104 14112 49112 14176
rect 49176 14112 49192 14176
rect 49256 14112 49272 14176
rect 49336 14112 49352 14176
rect 49416 14112 49424 14176
rect 49104 14111 49424 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 20208 13632 20528 13633
rect 20208 13568 20216 13632
rect 20280 13568 20296 13632
rect 20360 13568 20376 13632
rect 20440 13568 20456 13632
rect 20520 13568 20528 13632
rect 20208 13567 20528 13568
rect 39472 13632 39792 13633
rect 39472 13568 39480 13632
rect 39544 13568 39560 13632
rect 39624 13568 39640 13632
rect 39704 13568 39720 13632
rect 39784 13568 39792 13632
rect 39472 13567 39792 13568
rect 10576 13088 10896 13089
rect 0 13018 800 13048
rect 10576 13024 10584 13088
rect 10648 13024 10664 13088
rect 10728 13024 10744 13088
rect 10808 13024 10824 13088
rect 10888 13024 10896 13088
rect 10576 13023 10896 13024
rect 29840 13088 30160 13089
rect 29840 13024 29848 13088
rect 29912 13024 29928 13088
rect 29992 13024 30008 13088
rect 30072 13024 30088 13088
rect 30152 13024 30160 13088
rect 29840 13023 30160 13024
rect 49104 13088 49424 13089
rect 49104 13024 49112 13088
rect 49176 13024 49192 13088
rect 49256 13024 49272 13088
rect 49336 13024 49352 13088
rect 49416 13024 49424 13088
rect 49104 13023 49424 13024
rect 1393 13018 1459 13021
rect 0 13016 1459 13018
rect 0 12960 1398 13016
rect 1454 12960 1459 13016
rect 0 12958 1459 12960
rect 0 12928 800 12958
rect 1393 12955 1459 12958
rect 57881 13018 57947 13021
rect 59200 13018 60000 13048
rect 57881 13016 60000 13018
rect 57881 12960 57886 13016
rect 57942 12960 60000 13016
rect 57881 12958 60000 12960
rect 57881 12955 57947 12958
rect 59200 12928 60000 12958
rect 20208 12544 20528 12545
rect 20208 12480 20216 12544
rect 20280 12480 20296 12544
rect 20360 12480 20376 12544
rect 20440 12480 20456 12544
rect 20520 12480 20528 12544
rect 20208 12479 20528 12480
rect 39472 12544 39792 12545
rect 39472 12480 39480 12544
rect 39544 12480 39560 12544
rect 39624 12480 39640 12544
rect 39704 12480 39720 12544
rect 39784 12480 39792 12544
rect 39472 12479 39792 12480
rect 58157 12338 58223 12341
rect 59200 12338 60000 12368
rect 58157 12336 60000 12338
rect 58157 12280 58162 12336
rect 58218 12280 60000 12336
rect 58157 12278 60000 12280
rect 58157 12275 58223 12278
rect 59200 12248 60000 12278
rect 10576 12000 10896 12001
rect 10576 11936 10584 12000
rect 10648 11936 10664 12000
rect 10728 11936 10744 12000
rect 10808 11936 10824 12000
rect 10888 11936 10896 12000
rect 10576 11935 10896 11936
rect 29840 12000 30160 12001
rect 29840 11936 29848 12000
rect 29912 11936 29928 12000
rect 29992 11936 30008 12000
rect 30072 11936 30088 12000
rect 30152 11936 30160 12000
rect 29840 11935 30160 11936
rect 49104 12000 49424 12001
rect 49104 11936 49112 12000
rect 49176 11936 49192 12000
rect 49256 11936 49272 12000
rect 49336 11936 49352 12000
rect 49416 11936 49424 12000
rect 49104 11935 49424 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 58157 11658 58223 11661
rect 59200 11658 60000 11688
rect 58157 11656 60000 11658
rect 58157 11600 58162 11656
rect 58218 11600 60000 11656
rect 58157 11598 60000 11600
rect 58157 11595 58223 11598
rect 59200 11568 60000 11598
rect 20208 11456 20528 11457
rect 20208 11392 20216 11456
rect 20280 11392 20296 11456
rect 20360 11392 20376 11456
rect 20440 11392 20456 11456
rect 20520 11392 20528 11456
rect 20208 11391 20528 11392
rect 39472 11456 39792 11457
rect 39472 11392 39480 11456
rect 39544 11392 39560 11456
rect 39624 11392 39640 11456
rect 39704 11392 39720 11456
rect 39784 11392 39792 11456
rect 39472 11391 39792 11392
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 10576 10912 10896 10913
rect 10576 10848 10584 10912
rect 10648 10848 10664 10912
rect 10728 10848 10744 10912
rect 10808 10848 10824 10912
rect 10888 10848 10896 10912
rect 10576 10847 10896 10848
rect 29840 10912 30160 10913
rect 29840 10848 29848 10912
rect 29912 10848 29928 10912
rect 29992 10848 30008 10912
rect 30072 10848 30088 10912
rect 30152 10848 30160 10912
rect 29840 10847 30160 10848
rect 49104 10912 49424 10913
rect 49104 10848 49112 10912
rect 49176 10848 49192 10912
rect 49256 10848 49272 10912
rect 49336 10848 49352 10912
rect 49416 10848 49424 10912
rect 49104 10847 49424 10848
rect 20208 10368 20528 10369
rect 20208 10304 20216 10368
rect 20280 10304 20296 10368
rect 20360 10304 20376 10368
rect 20440 10304 20456 10368
rect 20520 10304 20528 10368
rect 20208 10303 20528 10304
rect 39472 10368 39792 10369
rect 39472 10304 39480 10368
rect 39544 10304 39560 10368
rect 39624 10304 39640 10368
rect 39704 10304 39720 10368
rect 39784 10304 39792 10368
rect 39472 10303 39792 10304
rect 58157 10298 58223 10301
rect 59200 10298 60000 10328
rect 58157 10296 60000 10298
rect 58157 10240 58162 10296
rect 58218 10240 60000 10296
rect 58157 10238 60000 10240
rect 58157 10235 58223 10238
rect 59200 10208 60000 10238
rect 10576 9824 10896 9825
rect 10576 9760 10584 9824
rect 10648 9760 10664 9824
rect 10728 9760 10744 9824
rect 10808 9760 10824 9824
rect 10888 9760 10896 9824
rect 10576 9759 10896 9760
rect 29840 9824 30160 9825
rect 29840 9760 29848 9824
rect 29912 9760 29928 9824
rect 29992 9760 30008 9824
rect 30072 9760 30088 9824
rect 30152 9760 30160 9824
rect 29840 9759 30160 9760
rect 49104 9824 49424 9825
rect 49104 9760 49112 9824
rect 49176 9760 49192 9824
rect 49256 9760 49272 9824
rect 49336 9760 49352 9824
rect 49416 9760 49424 9824
rect 49104 9759 49424 9760
rect 0 9618 800 9648
rect 1485 9618 1551 9621
rect 0 9616 1551 9618
rect 0 9560 1490 9616
rect 1546 9560 1551 9616
rect 0 9558 1551 9560
rect 0 9528 800 9558
rect 1485 9555 1551 9558
rect 58157 9618 58223 9621
rect 59200 9618 60000 9648
rect 58157 9616 60000 9618
rect 58157 9560 58162 9616
rect 58218 9560 60000 9616
rect 58157 9558 60000 9560
rect 58157 9555 58223 9558
rect 59200 9528 60000 9558
rect 20208 9280 20528 9281
rect 20208 9216 20216 9280
rect 20280 9216 20296 9280
rect 20360 9216 20376 9280
rect 20440 9216 20456 9280
rect 20520 9216 20528 9280
rect 20208 9215 20528 9216
rect 39472 9280 39792 9281
rect 39472 9216 39480 9280
rect 39544 9216 39560 9280
rect 39624 9216 39640 9280
rect 39704 9216 39720 9280
rect 39784 9216 39792 9280
rect 39472 9215 39792 9216
rect 0 8938 800 8968
rect 1393 8938 1459 8941
rect 0 8936 1459 8938
rect 0 8880 1398 8936
rect 1454 8880 1459 8936
rect 0 8878 1459 8880
rect 0 8848 800 8878
rect 1393 8875 1459 8878
rect 10576 8736 10896 8737
rect 10576 8672 10584 8736
rect 10648 8672 10664 8736
rect 10728 8672 10744 8736
rect 10808 8672 10824 8736
rect 10888 8672 10896 8736
rect 10576 8671 10896 8672
rect 29840 8736 30160 8737
rect 29840 8672 29848 8736
rect 29912 8672 29928 8736
rect 29992 8672 30008 8736
rect 30072 8672 30088 8736
rect 30152 8672 30160 8736
rect 29840 8671 30160 8672
rect 49104 8736 49424 8737
rect 49104 8672 49112 8736
rect 49176 8672 49192 8736
rect 49256 8672 49272 8736
rect 49336 8672 49352 8736
rect 49416 8672 49424 8736
rect 49104 8671 49424 8672
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 58157 8258 58223 8261
rect 59200 8258 60000 8288
rect 58157 8256 60000 8258
rect 58157 8200 58162 8256
rect 58218 8200 60000 8256
rect 58157 8198 60000 8200
rect 58157 8195 58223 8198
rect 20208 8192 20528 8193
rect 20208 8128 20216 8192
rect 20280 8128 20296 8192
rect 20360 8128 20376 8192
rect 20440 8128 20456 8192
rect 20520 8128 20528 8192
rect 20208 8127 20528 8128
rect 39472 8192 39792 8193
rect 39472 8128 39480 8192
rect 39544 8128 39560 8192
rect 39624 8128 39640 8192
rect 39704 8128 39720 8192
rect 39784 8128 39792 8192
rect 59200 8168 60000 8198
rect 39472 8127 39792 8128
rect 10576 7648 10896 7649
rect 10576 7584 10584 7648
rect 10648 7584 10664 7648
rect 10728 7584 10744 7648
rect 10808 7584 10824 7648
rect 10888 7584 10896 7648
rect 10576 7583 10896 7584
rect 29840 7648 30160 7649
rect 29840 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30160 7648
rect 29840 7583 30160 7584
rect 49104 7648 49424 7649
rect 49104 7584 49112 7648
rect 49176 7584 49192 7648
rect 49256 7584 49272 7648
rect 49336 7584 49352 7648
rect 49416 7584 49424 7648
rect 49104 7583 49424 7584
rect 58157 7578 58223 7581
rect 59200 7578 60000 7608
rect 58157 7576 60000 7578
rect 58157 7520 58162 7576
rect 58218 7520 60000 7576
rect 58157 7518 60000 7520
rect 58157 7515 58223 7518
rect 59200 7488 60000 7518
rect 20208 7104 20528 7105
rect 20208 7040 20216 7104
rect 20280 7040 20296 7104
rect 20360 7040 20376 7104
rect 20440 7040 20456 7104
rect 20520 7040 20528 7104
rect 20208 7039 20528 7040
rect 39472 7104 39792 7105
rect 39472 7040 39480 7104
rect 39544 7040 39560 7104
rect 39624 7040 39640 7104
rect 39704 7040 39720 7104
rect 39784 7040 39792 7104
rect 39472 7039 39792 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 58065 6898 58131 6901
rect 59200 6898 60000 6928
rect 58065 6896 60000 6898
rect 58065 6840 58070 6896
rect 58126 6840 60000 6896
rect 58065 6838 60000 6840
rect 58065 6835 58131 6838
rect 59200 6808 60000 6838
rect 10576 6560 10896 6561
rect 10576 6496 10584 6560
rect 10648 6496 10664 6560
rect 10728 6496 10744 6560
rect 10808 6496 10824 6560
rect 10888 6496 10896 6560
rect 10576 6495 10896 6496
rect 29840 6560 30160 6561
rect 29840 6496 29848 6560
rect 29912 6496 29928 6560
rect 29992 6496 30008 6560
rect 30072 6496 30088 6560
rect 30152 6496 30160 6560
rect 29840 6495 30160 6496
rect 49104 6560 49424 6561
rect 49104 6496 49112 6560
rect 49176 6496 49192 6560
rect 49256 6496 49272 6560
rect 49336 6496 49352 6560
rect 49416 6496 49424 6560
rect 49104 6495 49424 6496
rect 0 6218 800 6248
rect 1393 6218 1459 6221
rect 0 6216 1459 6218
rect 0 6160 1398 6216
rect 1454 6160 1459 6216
rect 0 6158 1459 6160
rect 0 6128 800 6158
rect 1393 6155 1459 6158
rect 20208 6016 20528 6017
rect 20208 5952 20216 6016
rect 20280 5952 20296 6016
rect 20360 5952 20376 6016
rect 20440 5952 20456 6016
rect 20520 5952 20528 6016
rect 20208 5951 20528 5952
rect 39472 6016 39792 6017
rect 39472 5952 39480 6016
rect 39544 5952 39560 6016
rect 39624 5952 39640 6016
rect 39704 5952 39720 6016
rect 39784 5952 39792 6016
rect 39472 5951 39792 5952
rect 58157 5538 58223 5541
rect 59200 5538 60000 5568
rect 58157 5536 60000 5538
rect 58157 5480 58162 5536
rect 58218 5480 60000 5536
rect 58157 5478 60000 5480
rect 58157 5475 58223 5478
rect 10576 5472 10896 5473
rect 10576 5408 10584 5472
rect 10648 5408 10664 5472
rect 10728 5408 10744 5472
rect 10808 5408 10824 5472
rect 10888 5408 10896 5472
rect 10576 5407 10896 5408
rect 29840 5472 30160 5473
rect 29840 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30160 5472
rect 29840 5407 30160 5408
rect 49104 5472 49424 5473
rect 49104 5408 49112 5472
rect 49176 5408 49192 5472
rect 49256 5408 49272 5472
rect 49336 5408 49352 5472
rect 49416 5408 49424 5472
rect 59200 5448 60000 5478
rect 49104 5407 49424 5408
rect 20208 4928 20528 4929
rect 0 4858 800 4888
rect 20208 4864 20216 4928
rect 20280 4864 20296 4928
rect 20360 4864 20376 4928
rect 20440 4864 20456 4928
rect 20520 4864 20528 4928
rect 20208 4863 20528 4864
rect 39472 4928 39792 4929
rect 39472 4864 39480 4928
rect 39544 4864 39560 4928
rect 39624 4864 39640 4928
rect 39704 4864 39720 4928
rect 39784 4864 39792 4928
rect 39472 4863 39792 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4768 800 4798
rect 1393 4795 1459 4798
rect 58065 4858 58131 4861
rect 59200 4858 60000 4888
rect 58065 4856 60000 4858
rect 58065 4800 58070 4856
rect 58126 4800 60000 4856
rect 58065 4798 60000 4800
rect 58065 4795 58131 4798
rect 59200 4768 60000 4798
rect 10576 4384 10896 4385
rect 10576 4320 10584 4384
rect 10648 4320 10664 4384
rect 10728 4320 10744 4384
rect 10808 4320 10824 4384
rect 10888 4320 10896 4384
rect 10576 4319 10896 4320
rect 29840 4384 30160 4385
rect 29840 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30160 4384
rect 29840 4319 30160 4320
rect 49104 4384 49424 4385
rect 49104 4320 49112 4384
rect 49176 4320 49192 4384
rect 49256 4320 49272 4384
rect 49336 4320 49352 4384
rect 49416 4320 49424 4384
rect 49104 4319 49424 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 57789 4178 57855 4181
rect 59200 4178 60000 4208
rect 57789 4176 60000 4178
rect 57789 4120 57794 4176
rect 57850 4120 60000 4176
rect 57789 4118 60000 4120
rect 57789 4115 57855 4118
rect 59200 4088 60000 4118
rect 20208 3840 20528 3841
rect 20208 3776 20216 3840
rect 20280 3776 20296 3840
rect 20360 3776 20376 3840
rect 20440 3776 20456 3840
rect 20520 3776 20528 3840
rect 20208 3775 20528 3776
rect 39472 3840 39792 3841
rect 39472 3776 39480 3840
rect 39544 3776 39560 3840
rect 39624 3776 39640 3840
rect 39704 3776 39720 3840
rect 39784 3776 39792 3840
rect 39472 3775 39792 3776
rect 0 3498 800 3528
rect 1393 3498 1459 3501
rect 0 3496 1459 3498
rect 0 3440 1398 3496
rect 1454 3440 1459 3496
rect 0 3438 1459 3440
rect 0 3408 800 3438
rect 1393 3435 1459 3438
rect 10576 3296 10896 3297
rect 10576 3232 10584 3296
rect 10648 3232 10664 3296
rect 10728 3232 10744 3296
rect 10808 3232 10824 3296
rect 10888 3232 10896 3296
rect 10576 3231 10896 3232
rect 29840 3296 30160 3297
rect 29840 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30160 3296
rect 29840 3231 30160 3232
rect 49104 3296 49424 3297
rect 49104 3232 49112 3296
rect 49176 3232 49192 3296
rect 49256 3232 49272 3296
rect 49336 3232 49352 3296
rect 49416 3232 49424 3296
rect 49104 3231 49424 3232
rect 16021 3090 16087 3093
rect 49693 3090 49759 3093
rect 16021 3088 49759 3090
rect 16021 3032 16026 3088
rect 16082 3032 49698 3088
rect 49754 3032 49759 3088
rect 16021 3030 49759 3032
rect 16021 3027 16087 3030
rect 49693 3027 49759 3030
rect 5717 2954 5783 2957
rect 43621 2954 43687 2957
rect 5717 2952 43687 2954
rect 5717 2896 5722 2952
rect 5778 2896 43626 2952
rect 43682 2896 43687 2952
rect 5717 2894 43687 2896
rect 5717 2891 5783 2894
rect 43621 2891 43687 2894
rect 57881 2818 57947 2821
rect 59200 2818 60000 2848
rect 57881 2816 60000 2818
rect 57881 2760 57886 2816
rect 57942 2760 60000 2816
rect 57881 2758 60000 2760
rect 57881 2755 57947 2758
rect 20208 2752 20528 2753
rect 20208 2688 20216 2752
rect 20280 2688 20296 2752
rect 20360 2688 20376 2752
rect 20440 2688 20456 2752
rect 20520 2688 20528 2752
rect 20208 2687 20528 2688
rect 39472 2752 39792 2753
rect 39472 2688 39480 2752
rect 39544 2688 39560 2752
rect 39624 2688 39640 2752
rect 39704 2688 39720 2752
rect 39784 2688 39792 2752
rect 59200 2728 60000 2758
rect 39472 2687 39792 2688
rect 12157 2682 12223 2685
rect 15285 2682 15351 2685
rect 12157 2680 15351 2682
rect 12157 2624 12162 2680
rect 12218 2624 15290 2680
rect 15346 2624 15351 2680
rect 12157 2622 15351 2624
rect 12157 2619 12223 2622
rect 15285 2619 15351 2622
rect 5165 2410 5231 2413
rect 57697 2410 57763 2413
rect 5165 2408 57763 2410
rect 5165 2352 5170 2408
rect 5226 2352 57702 2408
rect 57758 2352 57763 2408
rect 5165 2350 57763 2352
rect 5165 2347 5231 2350
rect 57697 2347 57763 2350
rect 10576 2208 10896 2209
rect 0 2138 800 2168
rect 10576 2144 10584 2208
rect 10648 2144 10664 2208
rect 10728 2144 10744 2208
rect 10808 2144 10824 2208
rect 10888 2144 10896 2208
rect 10576 2143 10896 2144
rect 29840 2208 30160 2209
rect 29840 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30160 2208
rect 29840 2143 30160 2144
rect 49104 2208 49424 2209
rect 49104 2144 49112 2208
rect 49176 2144 49192 2208
rect 49256 2144 49272 2208
rect 49336 2144 49352 2208
rect 49416 2144 49424 2208
rect 49104 2143 49424 2144
rect 2589 2138 2655 2141
rect 0 2136 2655 2138
rect 0 2080 2594 2136
rect 2650 2080 2655 2136
rect 0 2078 2655 2080
rect 0 2048 800 2078
rect 2589 2075 2655 2078
rect 56409 2138 56475 2141
rect 59200 2138 60000 2168
rect 56409 2136 60000 2138
rect 56409 2080 56414 2136
rect 56470 2080 60000 2136
rect 56409 2078 60000 2080
rect 56409 2075 56475 2078
rect 59200 2048 60000 2078
rect 0 1458 800 1488
rect 1485 1458 1551 1461
rect 0 1456 1551 1458
rect 0 1400 1490 1456
rect 1546 1400 1551 1456
rect 0 1398 1551 1400
rect 0 1368 800 1398
rect 1485 1395 1551 1398
rect 57605 778 57671 781
rect 59200 778 60000 808
rect 57605 776 60000 778
rect 57605 720 57610 776
rect 57666 720 60000 776
rect 57605 718 60000 720
rect 57605 715 57671 718
rect 59200 688 60000 718
<< via3 >>
rect 20216 27772 20280 27776
rect 20216 27716 20220 27772
rect 20220 27716 20276 27772
rect 20276 27716 20280 27772
rect 20216 27712 20280 27716
rect 20296 27772 20360 27776
rect 20296 27716 20300 27772
rect 20300 27716 20356 27772
rect 20356 27716 20360 27772
rect 20296 27712 20360 27716
rect 20376 27772 20440 27776
rect 20376 27716 20380 27772
rect 20380 27716 20436 27772
rect 20436 27716 20440 27772
rect 20376 27712 20440 27716
rect 20456 27772 20520 27776
rect 20456 27716 20460 27772
rect 20460 27716 20516 27772
rect 20516 27716 20520 27772
rect 20456 27712 20520 27716
rect 39480 27772 39544 27776
rect 39480 27716 39484 27772
rect 39484 27716 39540 27772
rect 39540 27716 39544 27772
rect 39480 27712 39544 27716
rect 39560 27772 39624 27776
rect 39560 27716 39564 27772
rect 39564 27716 39620 27772
rect 39620 27716 39624 27772
rect 39560 27712 39624 27716
rect 39640 27772 39704 27776
rect 39640 27716 39644 27772
rect 39644 27716 39700 27772
rect 39700 27716 39704 27772
rect 39640 27712 39704 27716
rect 39720 27772 39784 27776
rect 39720 27716 39724 27772
rect 39724 27716 39780 27772
rect 39780 27716 39784 27772
rect 39720 27712 39784 27716
rect 10584 27228 10648 27232
rect 10584 27172 10588 27228
rect 10588 27172 10644 27228
rect 10644 27172 10648 27228
rect 10584 27168 10648 27172
rect 10664 27228 10728 27232
rect 10664 27172 10668 27228
rect 10668 27172 10724 27228
rect 10724 27172 10728 27228
rect 10664 27168 10728 27172
rect 10744 27228 10808 27232
rect 10744 27172 10748 27228
rect 10748 27172 10804 27228
rect 10804 27172 10808 27228
rect 10744 27168 10808 27172
rect 10824 27228 10888 27232
rect 10824 27172 10828 27228
rect 10828 27172 10884 27228
rect 10884 27172 10888 27228
rect 10824 27168 10888 27172
rect 29848 27228 29912 27232
rect 29848 27172 29852 27228
rect 29852 27172 29908 27228
rect 29908 27172 29912 27228
rect 29848 27168 29912 27172
rect 29928 27228 29992 27232
rect 29928 27172 29932 27228
rect 29932 27172 29988 27228
rect 29988 27172 29992 27228
rect 29928 27168 29992 27172
rect 30008 27228 30072 27232
rect 30008 27172 30012 27228
rect 30012 27172 30068 27228
rect 30068 27172 30072 27228
rect 30008 27168 30072 27172
rect 30088 27228 30152 27232
rect 30088 27172 30092 27228
rect 30092 27172 30148 27228
rect 30148 27172 30152 27228
rect 30088 27168 30152 27172
rect 49112 27228 49176 27232
rect 49112 27172 49116 27228
rect 49116 27172 49172 27228
rect 49172 27172 49176 27228
rect 49112 27168 49176 27172
rect 49192 27228 49256 27232
rect 49192 27172 49196 27228
rect 49196 27172 49252 27228
rect 49252 27172 49256 27228
rect 49192 27168 49256 27172
rect 49272 27228 49336 27232
rect 49272 27172 49276 27228
rect 49276 27172 49332 27228
rect 49332 27172 49336 27228
rect 49272 27168 49336 27172
rect 49352 27228 49416 27232
rect 49352 27172 49356 27228
rect 49356 27172 49412 27228
rect 49412 27172 49416 27228
rect 49352 27168 49416 27172
rect 20216 26684 20280 26688
rect 20216 26628 20220 26684
rect 20220 26628 20276 26684
rect 20276 26628 20280 26684
rect 20216 26624 20280 26628
rect 20296 26684 20360 26688
rect 20296 26628 20300 26684
rect 20300 26628 20356 26684
rect 20356 26628 20360 26684
rect 20296 26624 20360 26628
rect 20376 26684 20440 26688
rect 20376 26628 20380 26684
rect 20380 26628 20436 26684
rect 20436 26628 20440 26684
rect 20376 26624 20440 26628
rect 20456 26684 20520 26688
rect 20456 26628 20460 26684
rect 20460 26628 20516 26684
rect 20516 26628 20520 26684
rect 20456 26624 20520 26628
rect 39480 26684 39544 26688
rect 39480 26628 39484 26684
rect 39484 26628 39540 26684
rect 39540 26628 39544 26684
rect 39480 26624 39544 26628
rect 39560 26684 39624 26688
rect 39560 26628 39564 26684
rect 39564 26628 39620 26684
rect 39620 26628 39624 26684
rect 39560 26624 39624 26628
rect 39640 26684 39704 26688
rect 39640 26628 39644 26684
rect 39644 26628 39700 26684
rect 39700 26628 39704 26684
rect 39640 26624 39704 26628
rect 39720 26684 39784 26688
rect 39720 26628 39724 26684
rect 39724 26628 39780 26684
rect 39780 26628 39784 26684
rect 39720 26624 39784 26628
rect 10584 26140 10648 26144
rect 10584 26084 10588 26140
rect 10588 26084 10644 26140
rect 10644 26084 10648 26140
rect 10584 26080 10648 26084
rect 10664 26140 10728 26144
rect 10664 26084 10668 26140
rect 10668 26084 10724 26140
rect 10724 26084 10728 26140
rect 10664 26080 10728 26084
rect 10744 26140 10808 26144
rect 10744 26084 10748 26140
rect 10748 26084 10804 26140
rect 10804 26084 10808 26140
rect 10744 26080 10808 26084
rect 10824 26140 10888 26144
rect 10824 26084 10828 26140
rect 10828 26084 10884 26140
rect 10884 26084 10888 26140
rect 10824 26080 10888 26084
rect 29848 26140 29912 26144
rect 29848 26084 29852 26140
rect 29852 26084 29908 26140
rect 29908 26084 29912 26140
rect 29848 26080 29912 26084
rect 29928 26140 29992 26144
rect 29928 26084 29932 26140
rect 29932 26084 29988 26140
rect 29988 26084 29992 26140
rect 29928 26080 29992 26084
rect 30008 26140 30072 26144
rect 30008 26084 30012 26140
rect 30012 26084 30068 26140
rect 30068 26084 30072 26140
rect 30008 26080 30072 26084
rect 30088 26140 30152 26144
rect 30088 26084 30092 26140
rect 30092 26084 30148 26140
rect 30148 26084 30152 26140
rect 30088 26080 30152 26084
rect 49112 26140 49176 26144
rect 49112 26084 49116 26140
rect 49116 26084 49172 26140
rect 49172 26084 49176 26140
rect 49112 26080 49176 26084
rect 49192 26140 49256 26144
rect 49192 26084 49196 26140
rect 49196 26084 49252 26140
rect 49252 26084 49256 26140
rect 49192 26080 49256 26084
rect 49272 26140 49336 26144
rect 49272 26084 49276 26140
rect 49276 26084 49332 26140
rect 49332 26084 49336 26140
rect 49272 26080 49336 26084
rect 49352 26140 49416 26144
rect 49352 26084 49356 26140
rect 49356 26084 49412 26140
rect 49412 26084 49416 26140
rect 49352 26080 49416 26084
rect 20216 25596 20280 25600
rect 20216 25540 20220 25596
rect 20220 25540 20276 25596
rect 20276 25540 20280 25596
rect 20216 25536 20280 25540
rect 20296 25596 20360 25600
rect 20296 25540 20300 25596
rect 20300 25540 20356 25596
rect 20356 25540 20360 25596
rect 20296 25536 20360 25540
rect 20376 25596 20440 25600
rect 20376 25540 20380 25596
rect 20380 25540 20436 25596
rect 20436 25540 20440 25596
rect 20376 25536 20440 25540
rect 20456 25596 20520 25600
rect 20456 25540 20460 25596
rect 20460 25540 20516 25596
rect 20516 25540 20520 25596
rect 20456 25536 20520 25540
rect 39480 25596 39544 25600
rect 39480 25540 39484 25596
rect 39484 25540 39540 25596
rect 39540 25540 39544 25596
rect 39480 25536 39544 25540
rect 39560 25596 39624 25600
rect 39560 25540 39564 25596
rect 39564 25540 39620 25596
rect 39620 25540 39624 25596
rect 39560 25536 39624 25540
rect 39640 25596 39704 25600
rect 39640 25540 39644 25596
rect 39644 25540 39700 25596
rect 39700 25540 39704 25596
rect 39640 25536 39704 25540
rect 39720 25596 39784 25600
rect 39720 25540 39724 25596
rect 39724 25540 39780 25596
rect 39780 25540 39784 25596
rect 39720 25536 39784 25540
rect 10584 25052 10648 25056
rect 10584 24996 10588 25052
rect 10588 24996 10644 25052
rect 10644 24996 10648 25052
rect 10584 24992 10648 24996
rect 10664 25052 10728 25056
rect 10664 24996 10668 25052
rect 10668 24996 10724 25052
rect 10724 24996 10728 25052
rect 10664 24992 10728 24996
rect 10744 25052 10808 25056
rect 10744 24996 10748 25052
rect 10748 24996 10804 25052
rect 10804 24996 10808 25052
rect 10744 24992 10808 24996
rect 10824 25052 10888 25056
rect 10824 24996 10828 25052
rect 10828 24996 10884 25052
rect 10884 24996 10888 25052
rect 10824 24992 10888 24996
rect 29848 25052 29912 25056
rect 29848 24996 29852 25052
rect 29852 24996 29908 25052
rect 29908 24996 29912 25052
rect 29848 24992 29912 24996
rect 29928 25052 29992 25056
rect 29928 24996 29932 25052
rect 29932 24996 29988 25052
rect 29988 24996 29992 25052
rect 29928 24992 29992 24996
rect 30008 25052 30072 25056
rect 30008 24996 30012 25052
rect 30012 24996 30068 25052
rect 30068 24996 30072 25052
rect 30008 24992 30072 24996
rect 30088 25052 30152 25056
rect 30088 24996 30092 25052
rect 30092 24996 30148 25052
rect 30148 24996 30152 25052
rect 30088 24992 30152 24996
rect 49112 25052 49176 25056
rect 49112 24996 49116 25052
rect 49116 24996 49172 25052
rect 49172 24996 49176 25052
rect 49112 24992 49176 24996
rect 49192 25052 49256 25056
rect 49192 24996 49196 25052
rect 49196 24996 49252 25052
rect 49252 24996 49256 25052
rect 49192 24992 49256 24996
rect 49272 25052 49336 25056
rect 49272 24996 49276 25052
rect 49276 24996 49332 25052
rect 49332 24996 49336 25052
rect 49272 24992 49336 24996
rect 49352 25052 49416 25056
rect 49352 24996 49356 25052
rect 49356 24996 49412 25052
rect 49412 24996 49416 25052
rect 49352 24992 49416 24996
rect 20216 24508 20280 24512
rect 20216 24452 20220 24508
rect 20220 24452 20276 24508
rect 20276 24452 20280 24508
rect 20216 24448 20280 24452
rect 20296 24508 20360 24512
rect 20296 24452 20300 24508
rect 20300 24452 20356 24508
rect 20356 24452 20360 24508
rect 20296 24448 20360 24452
rect 20376 24508 20440 24512
rect 20376 24452 20380 24508
rect 20380 24452 20436 24508
rect 20436 24452 20440 24508
rect 20376 24448 20440 24452
rect 20456 24508 20520 24512
rect 20456 24452 20460 24508
rect 20460 24452 20516 24508
rect 20516 24452 20520 24508
rect 20456 24448 20520 24452
rect 39480 24508 39544 24512
rect 39480 24452 39484 24508
rect 39484 24452 39540 24508
rect 39540 24452 39544 24508
rect 39480 24448 39544 24452
rect 39560 24508 39624 24512
rect 39560 24452 39564 24508
rect 39564 24452 39620 24508
rect 39620 24452 39624 24508
rect 39560 24448 39624 24452
rect 39640 24508 39704 24512
rect 39640 24452 39644 24508
rect 39644 24452 39700 24508
rect 39700 24452 39704 24508
rect 39640 24448 39704 24452
rect 39720 24508 39784 24512
rect 39720 24452 39724 24508
rect 39724 24452 39780 24508
rect 39780 24452 39784 24508
rect 39720 24448 39784 24452
rect 10584 23964 10648 23968
rect 10584 23908 10588 23964
rect 10588 23908 10644 23964
rect 10644 23908 10648 23964
rect 10584 23904 10648 23908
rect 10664 23964 10728 23968
rect 10664 23908 10668 23964
rect 10668 23908 10724 23964
rect 10724 23908 10728 23964
rect 10664 23904 10728 23908
rect 10744 23964 10808 23968
rect 10744 23908 10748 23964
rect 10748 23908 10804 23964
rect 10804 23908 10808 23964
rect 10744 23904 10808 23908
rect 10824 23964 10888 23968
rect 10824 23908 10828 23964
rect 10828 23908 10884 23964
rect 10884 23908 10888 23964
rect 10824 23904 10888 23908
rect 29848 23964 29912 23968
rect 29848 23908 29852 23964
rect 29852 23908 29908 23964
rect 29908 23908 29912 23964
rect 29848 23904 29912 23908
rect 29928 23964 29992 23968
rect 29928 23908 29932 23964
rect 29932 23908 29988 23964
rect 29988 23908 29992 23964
rect 29928 23904 29992 23908
rect 30008 23964 30072 23968
rect 30008 23908 30012 23964
rect 30012 23908 30068 23964
rect 30068 23908 30072 23964
rect 30008 23904 30072 23908
rect 30088 23964 30152 23968
rect 30088 23908 30092 23964
rect 30092 23908 30148 23964
rect 30148 23908 30152 23964
rect 30088 23904 30152 23908
rect 49112 23964 49176 23968
rect 49112 23908 49116 23964
rect 49116 23908 49172 23964
rect 49172 23908 49176 23964
rect 49112 23904 49176 23908
rect 49192 23964 49256 23968
rect 49192 23908 49196 23964
rect 49196 23908 49252 23964
rect 49252 23908 49256 23964
rect 49192 23904 49256 23908
rect 49272 23964 49336 23968
rect 49272 23908 49276 23964
rect 49276 23908 49332 23964
rect 49332 23908 49336 23964
rect 49272 23904 49336 23908
rect 49352 23964 49416 23968
rect 49352 23908 49356 23964
rect 49356 23908 49412 23964
rect 49412 23908 49416 23964
rect 49352 23904 49416 23908
rect 20216 23420 20280 23424
rect 20216 23364 20220 23420
rect 20220 23364 20276 23420
rect 20276 23364 20280 23420
rect 20216 23360 20280 23364
rect 20296 23420 20360 23424
rect 20296 23364 20300 23420
rect 20300 23364 20356 23420
rect 20356 23364 20360 23420
rect 20296 23360 20360 23364
rect 20376 23420 20440 23424
rect 20376 23364 20380 23420
rect 20380 23364 20436 23420
rect 20436 23364 20440 23420
rect 20376 23360 20440 23364
rect 20456 23420 20520 23424
rect 20456 23364 20460 23420
rect 20460 23364 20516 23420
rect 20516 23364 20520 23420
rect 20456 23360 20520 23364
rect 39480 23420 39544 23424
rect 39480 23364 39484 23420
rect 39484 23364 39540 23420
rect 39540 23364 39544 23420
rect 39480 23360 39544 23364
rect 39560 23420 39624 23424
rect 39560 23364 39564 23420
rect 39564 23364 39620 23420
rect 39620 23364 39624 23420
rect 39560 23360 39624 23364
rect 39640 23420 39704 23424
rect 39640 23364 39644 23420
rect 39644 23364 39700 23420
rect 39700 23364 39704 23420
rect 39640 23360 39704 23364
rect 39720 23420 39784 23424
rect 39720 23364 39724 23420
rect 39724 23364 39780 23420
rect 39780 23364 39784 23420
rect 39720 23360 39784 23364
rect 10584 22876 10648 22880
rect 10584 22820 10588 22876
rect 10588 22820 10644 22876
rect 10644 22820 10648 22876
rect 10584 22816 10648 22820
rect 10664 22876 10728 22880
rect 10664 22820 10668 22876
rect 10668 22820 10724 22876
rect 10724 22820 10728 22876
rect 10664 22816 10728 22820
rect 10744 22876 10808 22880
rect 10744 22820 10748 22876
rect 10748 22820 10804 22876
rect 10804 22820 10808 22876
rect 10744 22816 10808 22820
rect 10824 22876 10888 22880
rect 10824 22820 10828 22876
rect 10828 22820 10884 22876
rect 10884 22820 10888 22876
rect 10824 22816 10888 22820
rect 29848 22876 29912 22880
rect 29848 22820 29852 22876
rect 29852 22820 29908 22876
rect 29908 22820 29912 22876
rect 29848 22816 29912 22820
rect 29928 22876 29992 22880
rect 29928 22820 29932 22876
rect 29932 22820 29988 22876
rect 29988 22820 29992 22876
rect 29928 22816 29992 22820
rect 30008 22876 30072 22880
rect 30008 22820 30012 22876
rect 30012 22820 30068 22876
rect 30068 22820 30072 22876
rect 30008 22816 30072 22820
rect 30088 22876 30152 22880
rect 30088 22820 30092 22876
rect 30092 22820 30148 22876
rect 30148 22820 30152 22876
rect 30088 22816 30152 22820
rect 49112 22876 49176 22880
rect 49112 22820 49116 22876
rect 49116 22820 49172 22876
rect 49172 22820 49176 22876
rect 49112 22816 49176 22820
rect 49192 22876 49256 22880
rect 49192 22820 49196 22876
rect 49196 22820 49252 22876
rect 49252 22820 49256 22876
rect 49192 22816 49256 22820
rect 49272 22876 49336 22880
rect 49272 22820 49276 22876
rect 49276 22820 49332 22876
rect 49332 22820 49336 22876
rect 49272 22816 49336 22820
rect 49352 22876 49416 22880
rect 49352 22820 49356 22876
rect 49356 22820 49412 22876
rect 49412 22820 49416 22876
rect 49352 22816 49416 22820
rect 20216 22332 20280 22336
rect 20216 22276 20220 22332
rect 20220 22276 20276 22332
rect 20276 22276 20280 22332
rect 20216 22272 20280 22276
rect 20296 22332 20360 22336
rect 20296 22276 20300 22332
rect 20300 22276 20356 22332
rect 20356 22276 20360 22332
rect 20296 22272 20360 22276
rect 20376 22332 20440 22336
rect 20376 22276 20380 22332
rect 20380 22276 20436 22332
rect 20436 22276 20440 22332
rect 20376 22272 20440 22276
rect 20456 22332 20520 22336
rect 20456 22276 20460 22332
rect 20460 22276 20516 22332
rect 20516 22276 20520 22332
rect 20456 22272 20520 22276
rect 39480 22332 39544 22336
rect 39480 22276 39484 22332
rect 39484 22276 39540 22332
rect 39540 22276 39544 22332
rect 39480 22272 39544 22276
rect 39560 22332 39624 22336
rect 39560 22276 39564 22332
rect 39564 22276 39620 22332
rect 39620 22276 39624 22332
rect 39560 22272 39624 22276
rect 39640 22332 39704 22336
rect 39640 22276 39644 22332
rect 39644 22276 39700 22332
rect 39700 22276 39704 22332
rect 39640 22272 39704 22276
rect 39720 22332 39784 22336
rect 39720 22276 39724 22332
rect 39724 22276 39780 22332
rect 39780 22276 39784 22332
rect 39720 22272 39784 22276
rect 10584 21788 10648 21792
rect 10584 21732 10588 21788
rect 10588 21732 10644 21788
rect 10644 21732 10648 21788
rect 10584 21728 10648 21732
rect 10664 21788 10728 21792
rect 10664 21732 10668 21788
rect 10668 21732 10724 21788
rect 10724 21732 10728 21788
rect 10664 21728 10728 21732
rect 10744 21788 10808 21792
rect 10744 21732 10748 21788
rect 10748 21732 10804 21788
rect 10804 21732 10808 21788
rect 10744 21728 10808 21732
rect 10824 21788 10888 21792
rect 10824 21732 10828 21788
rect 10828 21732 10884 21788
rect 10884 21732 10888 21788
rect 10824 21728 10888 21732
rect 29848 21788 29912 21792
rect 29848 21732 29852 21788
rect 29852 21732 29908 21788
rect 29908 21732 29912 21788
rect 29848 21728 29912 21732
rect 29928 21788 29992 21792
rect 29928 21732 29932 21788
rect 29932 21732 29988 21788
rect 29988 21732 29992 21788
rect 29928 21728 29992 21732
rect 30008 21788 30072 21792
rect 30008 21732 30012 21788
rect 30012 21732 30068 21788
rect 30068 21732 30072 21788
rect 30008 21728 30072 21732
rect 30088 21788 30152 21792
rect 30088 21732 30092 21788
rect 30092 21732 30148 21788
rect 30148 21732 30152 21788
rect 30088 21728 30152 21732
rect 49112 21788 49176 21792
rect 49112 21732 49116 21788
rect 49116 21732 49172 21788
rect 49172 21732 49176 21788
rect 49112 21728 49176 21732
rect 49192 21788 49256 21792
rect 49192 21732 49196 21788
rect 49196 21732 49252 21788
rect 49252 21732 49256 21788
rect 49192 21728 49256 21732
rect 49272 21788 49336 21792
rect 49272 21732 49276 21788
rect 49276 21732 49332 21788
rect 49332 21732 49336 21788
rect 49272 21728 49336 21732
rect 49352 21788 49416 21792
rect 49352 21732 49356 21788
rect 49356 21732 49412 21788
rect 49412 21732 49416 21788
rect 49352 21728 49416 21732
rect 20216 21244 20280 21248
rect 20216 21188 20220 21244
rect 20220 21188 20276 21244
rect 20276 21188 20280 21244
rect 20216 21184 20280 21188
rect 20296 21244 20360 21248
rect 20296 21188 20300 21244
rect 20300 21188 20356 21244
rect 20356 21188 20360 21244
rect 20296 21184 20360 21188
rect 20376 21244 20440 21248
rect 20376 21188 20380 21244
rect 20380 21188 20436 21244
rect 20436 21188 20440 21244
rect 20376 21184 20440 21188
rect 20456 21244 20520 21248
rect 20456 21188 20460 21244
rect 20460 21188 20516 21244
rect 20516 21188 20520 21244
rect 20456 21184 20520 21188
rect 39480 21244 39544 21248
rect 39480 21188 39484 21244
rect 39484 21188 39540 21244
rect 39540 21188 39544 21244
rect 39480 21184 39544 21188
rect 39560 21244 39624 21248
rect 39560 21188 39564 21244
rect 39564 21188 39620 21244
rect 39620 21188 39624 21244
rect 39560 21184 39624 21188
rect 39640 21244 39704 21248
rect 39640 21188 39644 21244
rect 39644 21188 39700 21244
rect 39700 21188 39704 21244
rect 39640 21184 39704 21188
rect 39720 21244 39784 21248
rect 39720 21188 39724 21244
rect 39724 21188 39780 21244
rect 39780 21188 39784 21244
rect 39720 21184 39784 21188
rect 10584 20700 10648 20704
rect 10584 20644 10588 20700
rect 10588 20644 10644 20700
rect 10644 20644 10648 20700
rect 10584 20640 10648 20644
rect 10664 20700 10728 20704
rect 10664 20644 10668 20700
rect 10668 20644 10724 20700
rect 10724 20644 10728 20700
rect 10664 20640 10728 20644
rect 10744 20700 10808 20704
rect 10744 20644 10748 20700
rect 10748 20644 10804 20700
rect 10804 20644 10808 20700
rect 10744 20640 10808 20644
rect 10824 20700 10888 20704
rect 10824 20644 10828 20700
rect 10828 20644 10884 20700
rect 10884 20644 10888 20700
rect 10824 20640 10888 20644
rect 29848 20700 29912 20704
rect 29848 20644 29852 20700
rect 29852 20644 29908 20700
rect 29908 20644 29912 20700
rect 29848 20640 29912 20644
rect 29928 20700 29992 20704
rect 29928 20644 29932 20700
rect 29932 20644 29988 20700
rect 29988 20644 29992 20700
rect 29928 20640 29992 20644
rect 30008 20700 30072 20704
rect 30008 20644 30012 20700
rect 30012 20644 30068 20700
rect 30068 20644 30072 20700
rect 30008 20640 30072 20644
rect 30088 20700 30152 20704
rect 30088 20644 30092 20700
rect 30092 20644 30148 20700
rect 30148 20644 30152 20700
rect 30088 20640 30152 20644
rect 49112 20700 49176 20704
rect 49112 20644 49116 20700
rect 49116 20644 49172 20700
rect 49172 20644 49176 20700
rect 49112 20640 49176 20644
rect 49192 20700 49256 20704
rect 49192 20644 49196 20700
rect 49196 20644 49252 20700
rect 49252 20644 49256 20700
rect 49192 20640 49256 20644
rect 49272 20700 49336 20704
rect 49272 20644 49276 20700
rect 49276 20644 49332 20700
rect 49332 20644 49336 20700
rect 49272 20640 49336 20644
rect 49352 20700 49416 20704
rect 49352 20644 49356 20700
rect 49356 20644 49412 20700
rect 49412 20644 49416 20700
rect 49352 20640 49416 20644
rect 20216 20156 20280 20160
rect 20216 20100 20220 20156
rect 20220 20100 20276 20156
rect 20276 20100 20280 20156
rect 20216 20096 20280 20100
rect 20296 20156 20360 20160
rect 20296 20100 20300 20156
rect 20300 20100 20356 20156
rect 20356 20100 20360 20156
rect 20296 20096 20360 20100
rect 20376 20156 20440 20160
rect 20376 20100 20380 20156
rect 20380 20100 20436 20156
rect 20436 20100 20440 20156
rect 20376 20096 20440 20100
rect 20456 20156 20520 20160
rect 20456 20100 20460 20156
rect 20460 20100 20516 20156
rect 20516 20100 20520 20156
rect 20456 20096 20520 20100
rect 39480 20156 39544 20160
rect 39480 20100 39484 20156
rect 39484 20100 39540 20156
rect 39540 20100 39544 20156
rect 39480 20096 39544 20100
rect 39560 20156 39624 20160
rect 39560 20100 39564 20156
rect 39564 20100 39620 20156
rect 39620 20100 39624 20156
rect 39560 20096 39624 20100
rect 39640 20156 39704 20160
rect 39640 20100 39644 20156
rect 39644 20100 39700 20156
rect 39700 20100 39704 20156
rect 39640 20096 39704 20100
rect 39720 20156 39784 20160
rect 39720 20100 39724 20156
rect 39724 20100 39780 20156
rect 39780 20100 39784 20156
rect 39720 20096 39784 20100
rect 10584 19612 10648 19616
rect 10584 19556 10588 19612
rect 10588 19556 10644 19612
rect 10644 19556 10648 19612
rect 10584 19552 10648 19556
rect 10664 19612 10728 19616
rect 10664 19556 10668 19612
rect 10668 19556 10724 19612
rect 10724 19556 10728 19612
rect 10664 19552 10728 19556
rect 10744 19612 10808 19616
rect 10744 19556 10748 19612
rect 10748 19556 10804 19612
rect 10804 19556 10808 19612
rect 10744 19552 10808 19556
rect 10824 19612 10888 19616
rect 10824 19556 10828 19612
rect 10828 19556 10884 19612
rect 10884 19556 10888 19612
rect 10824 19552 10888 19556
rect 29848 19612 29912 19616
rect 29848 19556 29852 19612
rect 29852 19556 29908 19612
rect 29908 19556 29912 19612
rect 29848 19552 29912 19556
rect 29928 19612 29992 19616
rect 29928 19556 29932 19612
rect 29932 19556 29988 19612
rect 29988 19556 29992 19612
rect 29928 19552 29992 19556
rect 30008 19612 30072 19616
rect 30008 19556 30012 19612
rect 30012 19556 30068 19612
rect 30068 19556 30072 19612
rect 30008 19552 30072 19556
rect 30088 19612 30152 19616
rect 30088 19556 30092 19612
rect 30092 19556 30148 19612
rect 30148 19556 30152 19612
rect 30088 19552 30152 19556
rect 49112 19612 49176 19616
rect 49112 19556 49116 19612
rect 49116 19556 49172 19612
rect 49172 19556 49176 19612
rect 49112 19552 49176 19556
rect 49192 19612 49256 19616
rect 49192 19556 49196 19612
rect 49196 19556 49252 19612
rect 49252 19556 49256 19612
rect 49192 19552 49256 19556
rect 49272 19612 49336 19616
rect 49272 19556 49276 19612
rect 49276 19556 49332 19612
rect 49332 19556 49336 19612
rect 49272 19552 49336 19556
rect 49352 19612 49416 19616
rect 49352 19556 49356 19612
rect 49356 19556 49412 19612
rect 49412 19556 49416 19612
rect 49352 19552 49416 19556
rect 20216 19068 20280 19072
rect 20216 19012 20220 19068
rect 20220 19012 20276 19068
rect 20276 19012 20280 19068
rect 20216 19008 20280 19012
rect 20296 19068 20360 19072
rect 20296 19012 20300 19068
rect 20300 19012 20356 19068
rect 20356 19012 20360 19068
rect 20296 19008 20360 19012
rect 20376 19068 20440 19072
rect 20376 19012 20380 19068
rect 20380 19012 20436 19068
rect 20436 19012 20440 19068
rect 20376 19008 20440 19012
rect 20456 19068 20520 19072
rect 20456 19012 20460 19068
rect 20460 19012 20516 19068
rect 20516 19012 20520 19068
rect 20456 19008 20520 19012
rect 39480 19068 39544 19072
rect 39480 19012 39484 19068
rect 39484 19012 39540 19068
rect 39540 19012 39544 19068
rect 39480 19008 39544 19012
rect 39560 19068 39624 19072
rect 39560 19012 39564 19068
rect 39564 19012 39620 19068
rect 39620 19012 39624 19068
rect 39560 19008 39624 19012
rect 39640 19068 39704 19072
rect 39640 19012 39644 19068
rect 39644 19012 39700 19068
rect 39700 19012 39704 19068
rect 39640 19008 39704 19012
rect 39720 19068 39784 19072
rect 39720 19012 39724 19068
rect 39724 19012 39780 19068
rect 39780 19012 39784 19068
rect 39720 19008 39784 19012
rect 10584 18524 10648 18528
rect 10584 18468 10588 18524
rect 10588 18468 10644 18524
rect 10644 18468 10648 18524
rect 10584 18464 10648 18468
rect 10664 18524 10728 18528
rect 10664 18468 10668 18524
rect 10668 18468 10724 18524
rect 10724 18468 10728 18524
rect 10664 18464 10728 18468
rect 10744 18524 10808 18528
rect 10744 18468 10748 18524
rect 10748 18468 10804 18524
rect 10804 18468 10808 18524
rect 10744 18464 10808 18468
rect 10824 18524 10888 18528
rect 10824 18468 10828 18524
rect 10828 18468 10884 18524
rect 10884 18468 10888 18524
rect 10824 18464 10888 18468
rect 29848 18524 29912 18528
rect 29848 18468 29852 18524
rect 29852 18468 29908 18524
rect 29908 18468 29912 18524
rect 29848 18464 29912 18468
rect 29928 18524 29992 18528
rect 29928 18468 29932 18524
rect 29932 18468 29988 18524
rect 29988 18468 29992 18524
rect 29928 18464 29992 18468
rect 30008 18524 30072 18528
rect 30008 18468 30012 18524
rect 30012 18468 30068 18524
rect 30068 18468 30072 18524
rect 30008 18464 30072 18468
rect 30088 18524 30152 18528
rect 30088 18468 30092 18524
rect 30092 18468 30148 18524
rect 30148 18468 30152 18524
rect 30088 18464 30152 18468
rect 49112 18524 49176 18528
rect 49112 18468 49116 18524
rect 49116 18468 49172 18524
rect 49172 18468 49176 18524
rect 49112 18464 49176 18468
rect 49192 18524 49256 18528
rect 49192 18468 49196 18524
rect 49196 18468 49252 18524
rect 49252 18468 49256 18524
rect 49192 18464 49256 18468
rect 49272 18524 49336 18528
rect 49272 18468 49276 18524
rect 49276 18468 49332 18524
rect 49332 18468 49336 18524
rect 49272 18464 49336 18468
rect 49352 18524 49416 18528
rect 49352 18468 49356 18524
rect 49356 18468 49412 18524
rect 49412 18468 49416 18524
rect 49352 18464 49416 18468
rect 20216 17980 20280 17984
rect 20216 17924 20220 17980
rect 20220 17924 20276 17980
rect 20276 17924 20280 17980
rect 20216 17920 20280 17924
rect 20296 17980 20360 17984
rect 20296 17924 20300 17980
rect 20300 17924 20356 17980
rect 20356 17924 20360 17980
rect 20296 17920 20360 17924
rect 20376 17980 20440 17984
rect 20376 17924 20380 17980
rect 20380 17924 20436 17980
rect 20436 17924 20440 17980
rect 20376 17920 20440 17924
rect 20456 17980 20520 17984
rect 20456 17924 20460 17980
rect 20460 17924 20516 17980
rect 20516 17924 20520 17980
rect 20456 17920 20520 17924
rect 39480 17980 39544 17984
rect 39480 17924 39484 17980
rect 39484 17924 39540 17980
rect 39540 17924 39544 17980
rect 39480 17920 39544 17924
rect 39560 17980 39624 17984
rect 39560 17924 39564 17980
rect 39564 17924 39620 17980
rect 39620 17924 39624 17980
rect 39560 17920 39624 17924
rect 39640 17980 39704 17984
rect 39640 17924 39644 17980
rect 39644 17924 39700 17980
rect 39700 17924 39704 17980
rect 39640 17920 39704 17924
rect 39720 17980 39784 17984
rect 39720 17924 39724 17980
rect 39724 17924 39780 17980
rect 39780 17924 39784 17980
rect 39720 17920 39784 17924
rect 10584 17436 10648 17440
rect 10584 17380 10588 17436
rect 10588 17380 10644 17436
rect 10644 17380 10648 17436
rect 10584 17376 10648 17380
rect 10664 17436 10728 17440
rect 10664 17380 10668 17436
rect 10668 17380 10724 17436
rect 10724 17380 10728 17436
rect 10664 17376 10728 17380
rect 10744 17436 10808 17440
rect 10744 17380 10748 17436
rect 10748 17380 10804 17436
rect 10804 17380 10808 17436
rect 10744 17376 10808 17380
rect 10824 17436 10888 17440
rect 10824 17380 10828 17436
rect 10828 17380 10884 17436
rect 10884 17380 10888 17436
rect 10824 17376 10888 17380
rect 29848 17436 29912 17440
rect 29848 17380 29852 17436
rect 29852 17380 29908 17436
rect 29908 17380 29912 17436
rect 29848 17376 29912 17380
rect 29928 17436 29992 17440
rect 29928 17380 29932 17436
rect 29932 17380 29988 17436
rect 29988 17380 29992 17436
rect 29928 17376 29992 17380
rect 30008 17436 30072 17440
rect 30008 17380 30012 17436
rect 30012 17380 30068 17436
rect 30068 17380 30072 17436
rect 30008 17376 30072 17380
rect 30088 17436 30152 17440
rect 30088 17380 30092 17436
rect 30092 17380 30148 17436
rect 30148 17380 30152 17436
rect 30088 17376 30152 17380
rect 49112 17436 49176 17440
rect 49112 17380 49116 17436
rect 49116 17380 49172 17436
rect 49172 17380 49176 17436
rect 49112 17376 49176 17380
rect 49192 17436 49256 17440
rect 49192 17380 49196 17436
rect 49196 17380 49252 17436
rect 49252 17380 49256 17436
rect 49192 17376 49256 17380
rect 49272 17436 49336 17440
rect 49272 17380 49276 17436
rect 49276 17380 49332 17436
rect 49332 17380 49336 17436
rect 49272 17376 49336 17380
rect 49352 17436 49416 17440
rect 49352 17380 49356 17436
rect 49356 17380 49412 17436
rect 49412 17380 49416 17436
rect 49352 17376 49416 17380
rect 20216 16892 20280 16896
rect 20216 16836 20220 16892
rect 20220 16836 20276 16892
rect 20276 16836 20280 16892
rect 20216 16832 20280 16836
rect 20296 16892 20360 16896
rect 20296 16836 20300 16892
rect 20300 16836 20356 16892
rect 20356 16836 20360 16892
rect 20296 16832 20360 16836
rect 20376 16892 20440 16896
rect 20376 16836 20380 16892
rect 20380 16836 20436 16892
rect 20436 16836 20440 16892
rect 20376 16832 20440 16836
rect 20456 16892 20520 16896
rect 20456 16836 20460 16892
rect 20460 16836 20516 16892
rect 20516 16836 20520 16892
rect 20456 16832 20520 16836
rect 39480 16892 39544 16896
rect 39480 16836 39484 16892
rect 39484 16836 39540 16892
rect 39540 16836 39544 16892
rect 39480 16832 39544 16836
rect 39560 16892 39624 16896
rect 39560 16836 39564 16892
rect 39564 16836 39620 16892
rect 39620 16836 39624 16892
rect 39560 16832 39624 16836
rect 39640 16892 39704 16896
rect 39640 16836 39644 16892
rect 39644 16836 39700 16892
rect 39700 16836 39704 16892
rect 39640 16832 39704 16836
rect 39720 16892 39784 16896
rect 39720 16836 39724 16892
rect 39724 16836 39780 16892
rect 39780 16836 39784 16892
rect 39720 16832 39784 16836
rect 10584 16348 10648 16352
rect 10584 16292 10588 16348
rect 10588 16292 10644 16348
rect 10644 16292 10648 16348
rect 10584 16288 10648 16292
rect 10664 16348 10728 16352
rect 10664 16292 10668 16348
rect 10668 16292 10724 16348
rect 10724 16292 10728 16348
rect 10664 16288 10728 16292
rect 10744 16348 10808 16352
rect 10744 16292 10748 16348
rect 10748 16292 10804 16348
rect 10804 16292 10808 16348
rect 10744 16288 10808 16292
rect 10824 16348 10888 16352
rect 10824 16292 10828 16348
rect 10828 16292 10884 16348
rect 10884 16292 10888 16348
rect 10824 16288 10888 16292
rect 29848 16348 29912 16352
rect 29848 16292 29852 16348
rect 29852 16292 29908 16348
rect 29908 16292 29912 16348
rect 29848 16288 29912 16292
rect 29928 16348 29992 16352
rect 29928 16292 29932 16348
rect 29932 16292 29988 16348
rect 29988 16292 29992 16348
rect 29928 16288 29992 16292
rect 30008 16348 30072 16352
rect 30008 16292 30012 16348
rect 30012 16292 30068 16348
rect 30068 16292 30072 16348
rect 30008 16288 30072 16292
rect 30088 16348 30152 16352
rect 30088 16292 30092 16348
rect 30092 16292 30148 16348
rect 30148 16292 30152 16348
rect 30088 16288 30152 16292
rect 49112 16348 49176 16352
rect 49112 16292 49116 16348
rect 49116 16292 49172 16348
rect 49172 16292 49176 16348
rect 49112 16288 49176 16292
rect 49192 16348 49256 16352
rect 49192 16292 49196 16348
rect 49196 16292 49252 16348
rect 49252 16292 49256 16348
rect 49192 16288 49256 16292
rect 49272 16348 49336 16352
rect 49272 16292 49276 16348
rect 49276 16292 49332 16348
rect 49332 16292 49336 16348
rect 49272 16288 49336 16292
rect 49352 16348 49416 16352
rect 49352 16292 49356 16348
rect 49356 16292 49412 16348
rect 49412 16292 49416 16348
rect 49352 16288 49416 16292
rect 20216 15804 20280 15808
rect 20216 15748 20220 15804
rect 20220 15748 20276 15804
rect 20276 15748 20280 15804
rect 20216 15744 20280 15748
rect 20296 15804 20360 15808
rect 20296 15748 20300 15804
rect 20300 15748 20356 15804
rect 20356 15748 20360 15804
rect 20296 15744 20360 15748
rect 20376 15804 20440 15808
rect 20376 15748 20380 15804
rect 20380 15748 20436 15804
rect 20436 15748 20440 15804
rect 20376 15744 20440 15748
rect 20456 15804 20520 15808
rect 20456 15748 20460 15804
rect 20460 15748 20516 15804
rect 20516 15748 20520 15804
rect 20456 15744 20520 15748
rect 39480 15804 39544 15808
rect 39480 15748 39484 15804
rect 39484 15748 39540 15804
rect 39540 15748 39544 15804
rect 39480 15744 39544 15748
rect 39560 15804 39624 15808
rect 39560 15748 39564 15804
rect 39564 15748 39620 15804
rect 39620 15748 39624 15804
rect 39560 15744 39624 15748
rect 39640 15804 39704 15808
rect 39640 15748 39644 15804
rect 39644 15748 39700 15804
rect 39700 15748 39704 15804
rect 39640 15744 39704 15748
rect 39720 15804 39784 15808
rect 39720 15748 39724 15804
rect 39724 15748 39780 15804
rect 39780 15748 39784 15804
rect 39720 15744 39784 15748
rect 10584 15260 10648 15264
rect 10584 15204 10588 15260
rect 10588 15204 10644 15260
rect 10644 15204 10648 15260
rect 10584 15200 10648 15204
rect 10664 15260 10728 15264
rect 10664 15204 10668 15260
rect 10668 15204 10724 15260
rect 10724 15204 10728 15260
rect 10664 15200 10728 15204
rect 10744 15260 10808 15264
rect 10744 15204 10748 15260
rect 10748 15204 10804 15260
rect 10804 15204 10808 15260
rect 10744 15200 10808 15204
rect 10824 15260 10888 15264
rect 10824 15204 10828 15260
rect 10828 15204 10884 15260
rect 10884 15204 10888 15260
rect 10824 15200 10888 15204
rect 29848 15260 29912 15264
rect 29848 15204 29852 15260
rect 29852 15204 29908 15260
rect 29908 15204 29912 15260
rect 29848 15200 29912 15204
rect 29928 15260 29992 15264
rect 29928 15204 29932 15260
rect 29932 15204 29988 15260
rect 29988 15204 29992 15260
rect 29928 15200 29992 15204
rect 30008 15260 30072 15264
rect 30008 15204 30012 15260
rect 30012 15204 30068 15260
rect 30068 15204 30072 15260
rect 30008 15200 30072 15204
rect 30088 15260 30152 15264
rect 30088 15204 30092 15260
rect 30092 15204 30148 15260
rect 30148 15204 30152 15260
rect 30088 15200 30152 15204
rect 49112 15260 49176 15264
rect 49112 15204 49116 15260
rect 49116 15204 49172 15260
rect 49172 15204 49176 15260
rect 49112 15200 49176 15204
rect 49192 15260 49256 15264
rect 49192 15204 49196 15260
rect 49196 15204 49252 15260
rect 49252 15204 49256 15260
rect 49192 15200 49256 15204
rect 49272 15260 49336 15264
rect 49272 15204 49276 15260
rect 49276 15204 49332 15260
rect 49332 15204 49336 15260
rect 49272 15200 49336 15204
rect 49352 15260 49416 15264
rect 49352 15204 49356 15260
rect 49356 15204 49412 15260
rect 49412 15204 49416 15260
rect 49352 15200 49416 15204
rect 20216 14716 20280 14720
rect 20216 14660 20220 14716
rect 20220 14660 20276 14716
rect 20276 14660 20280 14716
rect 20216 14656 20280 14660
rect 20296 14716 20360 14720
rect 20296 14660 20300 14716
rect 20300 14660 20356 14716
rect 20356 14660 20360 14716
rect 20296 14656 20360 14660
rect 20376 14716 20440 14720
rect 20376 14660 20380 14716
rect 20380 14660 20436 14716
rect 20436 14660 20440 14716
rect 20376 14656 20440 14660
rect 20456 14716 20520 14720
rect 20456 14660 20460 14716
rect 20460 14660 20516 14716
rect 20516 14660 20520 14716
rect 20456 14656 20520 14660
rect 39480 14716 39544 14720
rect 39480 14660 39484 14716
rect 39484 14660 39540 14716
rect 39540 14660 39544 14716
rect 39480 14656 39544 14660
rect 39560 14716 39624 14720
rect 39560 14660 39564 14716
rect 39564 14660 39620 14716
rect 39620 14660 39624 14716
rect 39560 14656 39624 14660
rect 39640 14716 39704 14720
rect 39640 14660 39644 14716
rect 39644 14660 39700 14716
rect 39700 14660 39704 14716
rect 39640 14656 39704 14660
rect 39720 14716 39784 14720
rect 39720 14660 39724 14716
rect 39724 14660 39780 14716
rect 39780 14660 39784 14716
rect 39720 14656 39784 14660
rect 10584 14172 10648 14176
rect 10584 14116 10588 14172
rect 10588 14116 10644 14172
rect 10644 14116 10648 14172
rect 10584 14112 10648 14116
rect 10664 14172 10728 14176
rect 10664 14116 10668 14172
rect 10668 14116 10724 14172
rect 10724 14116 10728 14172
rect 10664 14112 10728 14116
rect 10744 14172 10808 14176
rect 10744 14116 10748 14172
rect 10748 14116 10804 14172
rect 10804 14116 10808 14172
rect 10744 14112 10808 14116
rect 10824 14172 10888 14176
rect 10824 14116 10828 14172
rect 10828 14116 10884 14172
rect 10884 14116 10888 14172
rect 10824 14112 10888 14116
rect 29848 14172 29912 14176
rect 29848 14116 29852 14172
rect 29852 14116 29908 14172
rect 29908 14116 29912 14172
rect 29848 14112 29912 14116
rect 29928 14172 29992 14176
rect 29928 14116 29932 14172
rect 29932 14116 29988 14172
rect 29988 14116 29992 14172
rect 29928 14112 29992 14116
rect 30008 14172 30072 14176
rect 30008 14116 30012 14172
rect 30012 14116 30068 14172
rect 30068 14116 30072 14172
rect 30008 14112 30072 14116
rect 30088 14172 30152 14176
rect 30088 14116 30092 14172
rect 30092 14116 30148 14172
rect 30148 14116 30152 14172
rect 30088 14112 30152 14116
rect 49112 14172 49176 14176
rect 49112 14116 49116 14172
rect 49116 14116 49172 14172
rect 49172 14116 49176 14172
rect 49112 14112 49176 14116
rect 49192 14172 49256 14176
rect 49192 14116 49196 14172
rect 49196 14116 49252 14172
rect 49252 14116 49256 14172
rect 49192 14112 49256 14116
rect 49272 14172 49336 14176
rect 49272 14116 49276 14172
rect 49276 14116 49332 14172
rect 49332 14116 49336 14172
rect 49272 14112 49336 14116
rect 49352 14172 49416 14176
rect 49352 14116 49356 14172
rect 49356 14116 49412 14172
rect 49412 14116 49416 14172
rect 49352 14112 49416 14116
rect 20216 13628 20280 13632
rect 20216 13572 20220 13628
rect 20220 13572 20276 13628
rect 20276 13572 20280 13628
rect 20216 13568 20280 13572
rect 20296 13628 20360 13632
rect 20296 13572 20300 13628
rect 20300 13572 20356 13628
rect 20356 13572 20360 13628
rect 20296 13568 20360 13572
rect 20376 13628 20440 13632
rect 20376 13572 20380 13628
rect 20380 13572 20436 13628
rect 20436 13572 20440 13628
rect 20376 13568 20440 13572
rect 20456 13628 20520 13632
rect 20456 13572 20460 13628
rect 20460 13572 20516 13628
rect 20516 13572 20520 13628
rect 20456 13568 20520 13572
rect 39480 13628 39544 13632
rect 39480 13572 39484 13628
rect 39484 13572 39540 13628
rect 39540 13572 39544 13628
rect 39480 13568 39544 13572
rect 39560 13628 39624 13632
rect 39560 13572 39564 13628
rect 39564 13572 39620 13628
rect 39620 13572 39624 13628
rect 39560 13568 39624 13572
rect 39640 13628 39704 13632
rect 39640 13572 39644 13628
rect 39644 13572 39700 13628
rect 39700 13572 39704 13628
rect 39640 13568 39704 13572
rect 39720 13628 39784 13632
rect 39720 13572 39724 13628
rect 39724 13572 39780 13628
rect 39780 13572 39784 13628
rect 39720 13568 39784 13572
rect 10584 13084 10648 13088
rect 10584 13028 10588 13084
rect 10588 13028 10644 13084
rect 10644 13028 10648 13084
rect 10584 13024 10648 13028
rect 10664 13084 10728 13088
rect 10664 13028 10668 13084
rect 10668 13028 10724 13084
rect 10724 13028 10728 13084
rect 10664 13024 10728 13028
rect 10744 13084 10808 13088
rect 10744 13028 10748 13084
rect 10748 13028 10804 13084
rect 10804 13028 10808 13084
rect 10744 13024 10808 13028
rect 10824 13084 10888 13088
rect 10824 13028 10828 13084
rect 10828 13028 10884 13084
rect 10884 13028 10888 13084
rect 10824 13024 10888 13028
rect 29848 13084 29912 13088
rect 29848 13028 29852 13084
rect 29852 13028 29908 13084
rect 29908 13028 29912 13084
rect 29848 13024 29912 13028
rect 29928 13084 29992 13088
rect 29928 13028 29932 13084
rect 29932 13028 29988 13084
rect 29988 13028 29992 13084
rect 29928 13024 29992 13028
rect 30008 13084 30072 13088
rect 30008 13028 30012 13084
rect 30012 13028 30068 13084
rect 30068 13028 30072 13084
rect 30008 13024 30072 13028
rect 30088 13084 30152 13088
rect 30088 13028 30092 13084
rect 30092 13028 30148 13084
rect 30148 13028 30152 13084
rect 30088 13024 30152 13028
rect 49112 13084 49176 13088
rect 49112 13028 49116 13084
rect 49116 13028 49172 13084
rect 49172 13028 49176 13084
rect 49112 13024 49176 13028
rect 49192 13084 49256 13088
rect 49192 13028 49196 13084
rect 49196 13028 49252 13084
rect 49252 13028 49256 13084
rect 49192 13024 49256 13028
rect 49272 13084 49336 13088
rect 49272 13028 49276 13084
rect 49276 13028 49332 13084
rect 49332 13028 49336 13084
rect 49272 13024 49336 13028
rect 49352 13084 49416 13088
rect 49352 13028 49356 13084
rect 49356 13028 49412 13084
rect 49412 13028 49416 13084
rect 49352 13024 49416 13028
rect 20216 12540 20280 12544
rect 20216 12484 20220 12540
rect 20220 12484 20276 12540
rect 20276 12484 20280 12540
rect 20216 12480 20280 12484
rect 20296 12540 20360 12544
rect 20296 12484 20300 12540
rect 20300 12484 20356 12540
rect 20356 12484 20360 12540
rect 20296 12480 20360 12484
rect 20376 12540 20440 12544
rect 20376 12484 20380 12540
rect 20380 12484 20436 12540
rect 20436 12484 20440 12540
rect 20376 12480 20440 12484
rect 20456 12540 20520 12544
rect 20456 12484 20460 12540
rect 20460 12484 20516 12540
rect 20516 12484 20520 12540
rect 20456 12480 20520 12484
rect 39480 12540 39544 12544
rect 39480 12484 39484 12540
rect 39484 12484 39540 12540
rect 39540 12484 39544 12540
rect 39480 12480 39544 12484
rect 39560 12540 39624 12544
rect 39560 12484 39564 12540
rect 39564 12484 39620 12540
rect 39620 12484 39624 12540
rect 39560 12480 39624 12484
rect 39640 12540 39704 12544
rect 39640 12484 39644 12540
rect 39644 12484 39700 12540
rect 39700 12484 39704 12540
rect 39640 12480 39704 12484
rect 39720 12540 39784 12544
rect 39720 12484 39724 12540
rect 39724 12484 39780 12540
rect 39780 12484 39784 12540
rect 39720 12480 39784 12484
rect 10584 11996 10648 12000
rect 10584 11940 10588 11996
rect 10588 11940 10644 11996
rect 10644 11940 10648 11996
rect 10584 11936 10648 11940
rect 10664 11996 10728 12000
rect 10664 11940 10668 11996
rect 10668 11940 10724 11996
rect 10724 11940 10728 11996
rect 10664 11936 10728 11940
rect 10744 11996 10808 12000
rect 10744 11940 10748 11996
rect 10748 11940 10804 11996
rect 10804 11940 10808 11996
rect 10744 11936 10808 11940
rect 10824 11996 10888 12000
rect 10824 11940 10828 11996
rect 10828 11940 10884 11996
rect 10884 11940 10888 11996
rect 10824 11936 10888 11940
rect 29848 11996 29912 12000
rect 29848 11940 29852 11996
rect 29852 11940 29908 11996
rect 29908 11940 29912 11996
rect 29848 11936 29912 11940
rect 29928 11996 29992 12000
rect 29928 11940 29932 11996
rect 29932 11940 29988 11996
rect 29988 11940 29992 11996
rect 29928 11936 29992 11940
rect 30008 11996 30072 12000
rect 30008 11940 30012 11996
rect 30012 11940 30068 11996
rect 30068 11940 30072 11996
rect 30008 11936 30072 11940
rect 30088 11996 30152 12000
rect 30088 11940 30092 11996
rect 30092 11940 30148 11996
rect 30148 11940 30152 11996
rect 30088 11936 30152 11940
rect 49112 11996 49176 12000
rect 49112 11940 49116 11996
rect 49116 11940 49172 11996
rect 49172 11940 49176 11996
rect 49112 11936 49176 11940
rect 49192 11996 49256 12000
rect 49192 11940 49196 11996
rect 49196 11940 49252 11996
rect 49252 11940 49256 11996
rect 49192 11936 49256 11940
rect 49272 11996 49336 12000
rect 49272 11940 49276 11996
rect 49276 11940 49332 11996
rect 49332 11940 49336 11996
rect 49272 11936 49336 11940
rect 49352 11996 49416 12000
rect 49352 11940 49356 11996
rect 49356 11940 49412 11996
rect 49412 11940 49416 11996
rect 49352 11936 49416 11940
rect 20216 11452 20280 11456
rect 20216 11396 20220 11452
rect 20220 11396 20276 11452
rect 20276 11396 20280 11452
rect 20216 11392 20280 11396
rect 20296 11452 20360 11456
rect 20296 11396 20300 11452
rect 20300 11396 20356 11452
rect 20356 11396 20360 11452
rect 20296 11392 20360 11396
rect 20376 11452 20440 11456
rect 20376 11396 20380 11452
rect 20380 11396 20436 11452
rect 20436 11396 20440 11452
rect 20376 11392 20440 11396
rect 20456 11452 20520 11456
rect 20456 11396 20460 11452
rect 20460 11396 20516 11452
rect 20516 11396 20520 11452
rect 20456 11392 20520 11396
rect 39480 11452 39544 11456
rect 39480 11396 39484 11452
rect 39484 11396 39540 11452
rect 39540 11396 39544 11452
rect 39480 11392 39544 11396
rect 39560 11452 39624 11456
rect 39560 11396 39564 11452
rect 39564 11396 39620 11452
rect 39620 11396 39624 11452
rect 39560 11392 39624 11396
rect 39640 11452 39704 11456
rect 39640 11396 39644 11452
rect 39644 11396 39700 11452
rect 39700 11396 39704 11452
rect 39640 11392 39704 11396
rect 39720 11452 39784 11456
rect 39720 11396 39724 11452
rect 39724 11396 39780 11452
rect 39780 11396 39784 11452
rect 39720 11392 39784 11396
rect 10584 10908 10648 10912
rect 10584 10852 10588 10908
rect 10588 10852 10644 10908
rect 10644 10852 10648 10908
rect 10584 10848 10648 10852
rect 10664 10908 10728 10912
rect 10664 10852 10668 10908
rect 10668 10852 10724 10908
rect 10724 10852 10728 10908
rect 10664 10848 10728 10852
rect 10744 10908 10808 10912
rect 10744 10852 10748 10908
rect 10748 10852 10804 10908
rect 10804 10852 10808 10908
rect 10744 10848 10808 10852
rect 10824 10908 10888 10912
rect 10824 10852 10828 10908
rect 10828 10852 10884 10908
rect 10884 10852 10888 10908
rect 10824 10848 10888 10852
rect 29848 10908 29912 10912
rect 29848 10852 29852 10908
rect 29852 10852 29908 10908
rect 29908 10852 29912 10908
rect 29848 10848 29912 10852
rect 29928 10908 29992 10912
rect 29928 10852 29932 10908
rect 29932 10852 29988 10908
rect 29988 10852 29992 10908
rect 29928 10848 29992 10852
rect 30008 10908 30072 10912
rect 30008 10852 30012 10908
rect 30012 10852 30068 10908
rect 30068 10852 30072 10908
rect 30008 10848 30072 10852
rect 30088 10908 30152 10912
rect 30088 10852 30092 10908
rect 30092 10852 30148 10908
rect 30148 10852 30152 10908
rect 30088 10848 30152 10852
rect 49112 10908 49176 10912
rect 49112 10852 49116 10908
rect 49116 10852 49172 10908
rect 49172 10852 49176 10908
rect 49112 10848 49176 10852
rect 49192 10908 49256 10912
rect 49192 10852 49196 10908
rect 49196 10852 49252 10908
rect 49252 10852 49256 10908
rect 49192 10848 49256 10852
rect 49272 10908 49336 10912
rect 49272 10852 49276 10908
rect 49276 10852 49332 10908
rect 49332 10852 49336 10908
rect 49272 10848 49336 10852
rect 49352 10908 49416 10912
rect 49352 10852 49356 10908
rect 49356 10852 49412 10908
rect 49412 10852 49416 10908
rect 49352 10848 49416 10852
rect 20216 10364 20280 10368
rect 20216 10308 20220 10364
rect 20220 10308 20276 10364
rect 20276 10308 20280 10364
rect 20216 10304 20280 10308
rect 20296 10364 20360 10368
rect 20296 10308 20300 10364
rect 20300 10308 20356 10364
rect 20356 10308 20360 10364
rect 20296 10304 20360 10308
rect 20376 10364 20440 10368
rect 20376 10308 20380 10364
rect 20380 10308 20436 10364
rect 20436 10308 20440 10364
rect 20376 10304 20440 10308
rect 20456 10364 20520 10368
rect 20456 10308 20460 10364
rect 20460 10308 20516 10364
rect 20516 10308 20520 10364
rect 20456 10304 20520 10308
rect 39480 10364 39544 10368
rect 39480 10308 39484 10364
rect 39484 10308 39540 10364
rect 39540 10308 39544 10364
rect 39480 10304 39544 10308
rect 39560 10364 39624 10368
rect 39560 10308 39564 10364
rect 39564 10308 39620 10364
rect 39620 10308 39624 10364
rect 39560 10304 39624 10308
rect 39640 10364 39704 10368
rect 39640 10308 39644 10364
rect 39644 10308 39700 10364
rect 39700 10308 39704 10364
rect 39640 10304 39704 10308
rect 39720 10364 39784 10368
rect 39720 10308 39724 10364
rect 39724 10308 39780 10364
rect 39780 10308 39784 10364
rect 39720 10304 39784 10308
rect 10584 9820 10648 9824
rect 10584 9764 10588 9820
rect 10588 9764 10644 9820
rect 10644 9764 10648 9820
rect 10584 9760 10648 9764
rect 10664 9820 10728 9824
rect 10664 9764 10668 9820
rect 10668 9764 10724 9820
rect 10724 9764 10728 9820
rect 10664 9760 10728 9764
rect 10744 9820 10808 9824
rect 10744 9764 10748 9820
rect 10748 9764 10804 9820
rect 10804 9764 10808 9820
rect 10744 9760 10808 9764
rect 10824 9820 10888 9824
rect 10824 9764 10828 9820
rect 10828 9764 10884 9820
rect 10884 9764 10888 9820
rect 10824 9760 10888 9764
rect 29848 9820 29912 9824
rect 29848 9764 29852 9820
rect 29852 9764 29908 9820
rect 29908 9764 29912 9820
rect 29848 9760 29912 9764
rect 29928 9820 29992 9824
rect 29928 9764 29932 9820
rect 29932 9764 29988 9820
rect 29988 9764 29992 9820
rect 29928 9760 29992 9764
rect 30008 9820 30072 9824
rect 30008 9764 30012 9820
rect 30012 9764 30068 9820
rect 30068 9764 30072 9820
rect 30008 9760 30072 9764
rect 30088 9820 30152 9824
rect 30088 9764 30092 9820
rect 30092 9764 30148 9820
rect 30148 9764 30152 9820
rect 30088 9760 30152 9764
rect 49112 9820 49176 9824
rect 49112 9764 49116 9820
rect 49116 9764 49172 9820
rect 49172 9764 49176 9820
rect 49112 9760 49176 9764
rect 49192 9820 49256 9824
rect 49192 9764 49196 9820
rect 49196 9764 49252 9820
rect 49252 9764 49256 9820
rect 49192 9760 49256 9764
rect 49272 9820 49336 9824
rect 49272 9764 49276 9820
rect 49276 9764 49332 9820
rect 49332 9764 49336 9820
rect 49272 9760 49336 9764
rect 49352 9820 49416 9824
rect 49352 9764 49356 9820
rect 49356 9764 49412 9820
rect 49412 9764 49416 9820
rect 49352 9760 49416 9764
rect 20216 9276 20280 9280
rect 20216 9220 20220 9276
rect 20220 9220 20276 9276
rect 20276 9220 20280 9276
rect 20216 9216 20280 9220
rect 20296 9276 20360 9280
rect 20296 9220 20300 9276
rect 20300 9220 20356 9276
rect 20356 9220 20360 9276
rect 20296 9216 20360 9220
rect 20376 9276 20440 9280
rect 20376 9220 20380 9276
rect 20380 9220 20436 9276
rect 20436 9220 20440 9276
rect 20376 9216 20440 9220
rect 20456 9276 20520 9280
rect 20456 9220 20460 9276
rect 20460 9220 20516 9276
rect 20516 9220 20520 9276
rect 20456 9216 20520 9220
rect 39480 9276 39544 9280
rect 39480 9220 39484 9276
rect 39484 9220 39540 9276
rect 39540 9220 39544 9276
rect 39480 9216 39544 9220
rect 39560 9276 39624 9280
rect 39560 9220 39564 9276
rect 39564 9220 39620 9276
rect 39620 9220 39624 9276
rect 39560 9216 39624 9220
rect 39640 9276 39704 9280
rect 39640 9220 39644 9276
rect 39644 9220 39700 9276
rect 39700 9220 39704 9276
rect 39640 9216 39704 9220
rect 39720 9276 39784 9280
rect 39720 9220 39724 9276
rect 39724 9220 39780 9276
rect 39780 9220 39784 9276
rect 39720 9216 39784 9220
rect 10584 8732 10648 8736
rect 10584 8676 10588 8732
rect 10588 8676 10644 8732
rect 10644 8676 10648 8732
rect 10584 8672 10648 8676
rect 10664 8732 10728 8736
rect 10664 8676 10668 8732
rect 10668 8676 10724 8732
rect 10724 8676 10728 8732
rect 10664 8672 10728 8676
rect 10744 8732 10808 8736
rect 10744 8676 10748 8732
rect 10748 8676 10804 8732
rect 10804 8676 10808 8732
rect 10744 8672 10808 8676
rect 10824 8732 10888 8736
rect 10824 8676 10828 8732
rect 10828 8676 10884 8732
rect 10884 8676 10888 8732
rect 10824 8672 10888 8676
rect 29848 8732 29912 8736
rect 29848 8676 29852 8732
rect 29852 8676 29908 8732
rect 29908 8676 29912 8732
rect 29848 8672 29912 8676
rect 29928 8732 29992 8736
rect 29928 8676 29932 8732
rect 29932 8676 29988 8732
rect 29988 8676 29992 8732
rect 29928 8672 29992 8676
rect 30008 8732 30072 8736
rect 30008 8676 30012 8732
rect 30012 8676 30068 8732
rect 30068 8676 30072 8732
rect 30008 8672 30072 8676
rect 30088 8732 30152 8736
rect 30088 8676 30092 8732
rect 30092 8676 30148 8732
rect 30148 8676 30152 8732
rect 30088 8672 30152 8676
rect 49112 8732 49176 8736
rect 49112 8676 49116 8732
rect 49116 8676 49172 8732
rect 49172 8676 49176 8732
rect 49112 8672 49176 8676
rect 49192 8732 49256 8736
rect 49192 8676 49196 8732
rect 49196 8676 49252 8732
rect 49252 8676 49256 8732
rect 49192 8672 49256 8676
rect 49272 8732 49336 8736
rect 49272 8676 49276 8732
rect 49276 8676 49332 8732
rect 49332 8676 49336 8732
rect 49272 8672 49336 8676
rect 49352 8732 49416 8736
rect 49352 8676 49356 8732
rect 49356 8676 49412 8732
rect 49412 8676 49416 8732
rect 49352 8672 49416 8676
rect 20216 8188 20280 8192
rect 20216 8132 20220 8188
rect 20220 8132 20276 8188
rect 20276 8132 20280 8188
rect 20216 8128 20280 8132
rect 20296 8188 20360 8192
rect 20296 8132 20300 8188
rect 20300 8132 20356 8188
rect 20356 8132 20360 8188
rect 20296 8128 20360 8132
rect 20376 8188 20440 8192
rect 20376 8132 20380 8188
rect 20380 8132 20436 8188
rect 20436 8132 20440 8188
rect 20376 8128 20440 8132
rect 20456 8188 20520 8192
rect 20456 8132 20460 8188
rect 20460 8132 20516 8188
rect 20516 8132 20520 8188
rect 20456 8128 20520 8132
rect 39480 8188 39544 8192
rect 39480 8132 39484 8188
rect 39484 8132 39540 8188
rect 39540 8132 39544 8188
rect 39480 8128 39544 8132
rect 39560 8188 39624 8192
rect 39560 8132 39564 8188
rect 39564 8132 39620 8188
rect 39620 8132 39624 8188
rect 39560 8128 39624 8132
rect 39640 8188 39704 8192
rect 39640 8132 39644 8188
rect 39644 8132 39700 8188
rect 39700 8132 39704 8188
rect 39640 8128 39704 8132
rect 39720 8188 39784 8192
rect 39720 8132 39724 8188
rect 39724 8132 39780 8188
rect 39780 8132 39784 8188
rect 39720 8128 39784 8132
rect 10584 7644 10648 7648
rect 10584 7588 10588 7644
rect 10588 7588 10644 7644
rect 10644 7588 10648 7644
rect 10584 7584 10648 7588
rect 10664 7644 10728 7648
rect 10664 7588 10668 7644
rect 10668 7588 10724 7644
rect 10724 7588 10728 7644
rect 10664 7584 10728 7588
rect 10744 7644 10808 7648
rect 10744 7588 10748 7644
rect 10748 7588 10804 7644
rect 10804 7588 10808 7644
rect 10744 7584 10808 7588
rect 10824 7644 10888 7648
rect 10824 7588 10828 7644
rect 10828 7588 10884 7644
rect 10884 7588 10888 7644
rect 10824 7584 10888 7588
rect 29848 7644 29912 7648
rect 29848 7588 29852 7644
rect 29852 7588 29908 7644
rect 29908 7588 29912 7644
rect 29848 7584 29912 7588
rect 29928 7644 29992 7648
rect 29928 7588 29932 7644
rect 29932 7588 29988 7644
rect 29988 7588 29992 7644
rect 29928 7584 29992 7588
rect 30008 7644 30072 7648
rect 30008 7588 30012 7644
rect 30012 7588 30068 7644
rect 30068 7588 30072 7644
rect 30008 7584 30072 7588
rect 30088 7644 30152 7648
rect 30088 7588 30092 7644
rect 30092 7588 30148 7644
rect 30148 7588 30152 7644
rect 30088 7584 30152 7588
rect 49112 7644 49176 7648
rect 49112 7588 49116 7644
rect 49116 7588 49172 7644
rect 49172 7588 49176 7644
rect 49112 7584 49176 7588
rect 49192 7644 49256 7648
rect 49192 7588 49196 7644
rect 49196 7588 49252 7644
rect 49252 7588 49256 7644
rect 49192 7584 49256 7588
rect 49272 7644 49336 7648
rect 49272 7588 49276 7644
rect 49276 7588 49332 7644
rect 49332 7588 49336 7644
rect 49272 7584 49336 7588
rect 49352 7644 49416 7648
rect 49352 7588 49356 7644
rect 49356 7588 49412 7644
rect 49412 7588 49416 7644
rect 49352 7584 49416 7588
rect 20216 7100 20280 7104
rect 20216 7044 20220 7100
rect 20220 7044 20276 7100
rect 20276 7044 20280 7100
rect 20216 7040 20280 7044
rect 20296 7100 20360 7104
rect 20296 7044 20300 7100
rect 20300 7044 20356 7100
rect 20356 7044 20360 7100
rect 20296 7040 20360 7044
rect 20376 7100 20440 7104
rect 20376 7044 20380 7100
rect 20380 7044 20436 7100
rect 20436 7044 20440 7100
rect 20376 7040 20440 7044
rect 20456 7100 20520 7104
rect 20456 7044 20460 7100
rect 20460 7044 20516 7100
rect 20516 7044 20520 7100
rect 20456 7040 20520 7044
rect 39480 7100 39544 7104
rect 39480 7044 39484 7100
rect 39484 7044 39540 7100
rect 39540 7044 39544 7100
rect 39480 7040 39544 7044
rect 39560 7100 39624 7104
rect 39560 7044 39564 7100
rect 39564 7044 39620 7100
rect 39620 7044 39624 7100
rect 39560 7040 39624 7044
rect 39640 7100 39704 7104
rect 39640 7044 39644 7100
rect 39644 7044 39700 7100
rect 39700 7044 39704 7100
rect 39640 7040 39704 7044
rect 39720 7100 39784 7104
rect 39720 7044 39724 7100
rect 39724 7044 39780 7100
rect 39780 7044 39784 7100
rect 39720 7040 39784 7044
rect 10584 6556 10648 6560
rect 10584 6500 10588 6556
rect 10588 6500 10644 6556
rect 10644 6500 10648 6556
rect 10584 6496 10648 6500
rect 10664 6556 10728 6560
rect 10664 6500 10668 6556
rect 10668 6500 10724 6556
rect 10724 6500 10728 6556
rect 10664 6496 10728 6500
rect 10744 6556 10808 6560
rect 10744 6500 10748 6556
rect 10748 6500 10804 6556
rect 10804 6500 10808 6556
rect 10744 6496 10808 6500
rect 10824 6556 10888 6560
rect 10824 6500 10828 6556
rect 10828 6500 10884 6556
rect 10884 6500 10888 6556
rect 10824 6496 10888 6500
rect 29848 6556 29912 6560
rect 29848 6500 29852 6556
rect 29852 6500 29908 6556
rect 29908 6500 29912 6556
rect 29848 6496 29912 6500
rect 29928 6556 29992 6560
rect 29928 6500 29932 6556
rect 29932 6500 29988 6556
rect 29988 6500 29992 6556
rect 29928 6496 29992 6500
rect 30008 6556 30072 6560
rect 30008 6500 30012 6556
rect 30012 6500 30068 6556
rect 30068 6500 30072 6556
rect 30008 6496 30072 6500
rect 30088 6556 30152 6560
rect 30088 6500 30092 6556
rect 30092 6500 30148 6556
rect 30148 6500 30152 6556
rect 30088 6496 30152 6500
rect 49112 6556 49176 6560
rect 49112 6500 49116 6556
rect 49116 6500 49172 6556
rect 49172 6500 49176 6556
rect 49112 6496 49176 6500
rect 49192 6556 49256 6560
rect 49192 6500 49196 6556
rect 49196 6500 49252 6556
rect 49252 6500 49256 6556
rect 49192 6496 49256 6500
rect 49272 6556 49336 6560
rect 49272 6500 49276 6556
rect 49276 6500 49332 6556
rect 49332 6500 49336 6556
rect 49272 6496 49336 6500
rect 49352 6556 49416 6560
rect 49352 6500 49356 6556
rect 49356 6500 49412 6556
rect 49412 6500 49416 6556
rect 49352 6496 49416 6500
rect 20216 6012 20280 6016
rect 20216 5956 20220 6012
rect 20220 5956 20276 6012
rect 20276 5956 20280 6012
rect 20216 5952 20280 5956
rect 20296 6012 20360 6016
rect 20296 5956 20300 6012
rect 20300 5956 20356 6012
rect 20356 5956 20360 6012
rect 20296 5952 20360 5956
rect 20376 6012 20440 6016
rect 20376 5956 20380 6012
rect 20380 5956 20436 6012
rect 20436 5956 20440 6012
rect 20376 5952 20440 5956
rect 20456 6012 20520 6016
rect 20456 5956 20460 6012
rect 20460 5956 20516 6012
rect 20516 5956 20520 6012
rect 20456 5952 20520 5956
rect 39480 6012 39544 6016
rect 39480 5956 39484 6012
rect 39484 5956 39540 6012
rect 39540 5956 39544 6012
rect 39480 5952 39544 5956
rect 39560 6012 39624 6016
rect 39560 5956 39564 6012
rect 39564 5956 39620 6012
rect 39620 5956 39624 6012
rect 39560 5952 39624 5956
rect 39640 6012 39704 6016
rect 39640 5956 39644 6012
rect 39644 5956 39700 6012
rect 39700 5956 39704 6012
rect 39640 5952 39704 5956
rect 39720 6012 39784 6016
rect 39720 5956 39724 6012
rect 39724 5956 39780 6012
rect 39780 5956 39784 6012
rect 39720 5952 39784 5956
rect 10584 5468 10648 5472
rect 10584 5412 10588 5468
rect 10588 5412 10644 5468
rect 10644 5412 10648 5468
rect 10584 5408 10648 5412
rect 10664 5468 10728 5472
rect 10664 5412 10668 5468
rect 10668 5412 10724 5468
rect 10724 5412 10728 5468
rect 10664 5408 10728 5412
rect 10744 5468 10808 5472
rect 10744 5412 10748 5468
rect 10748 5412 10804 5468
rect 10804 5412 10808 5468
rect 10744 5408 10808 5412
rect 10824 5468 10888 5472
rect 10824 5412 10828 5468
rect 10828 5412 10884 5468
rect 10884 5412 10888 5468
rect 10824 5408 10888 5412
rect 29848 5468 29912 5472
rect 29848 5412 29852 5468
rect 29852 5412 29908 5468
rect 29908 5412 29912 5468
rect 29848 5408 29912 5412
rect 29928 5468 29992 5472
rect 29928 5412 29932 5468
rect 29932 5412 29988 5468
rect 29988 5412 29992 5468
rect 29928 5408 29992 5412
rect 30008 5468 30072 5472
rect 30008 5412 30012 5468
rect 30012 5412 30068 5468
rect 30068 5412 30072 5468
rect 30008 5408 30072 5412
rect 30088 5468 30152 5472
rect 30088 5412 30092 5468
rect 30092 5412 30148 5468
rect 30148 5412 30152 5468
rect 30088 5408 30152 5412
rect 49112 5468 49176 5472
rect 49112 5412 49116 5468
rect 49116 5412 49172 5468
rect 49172 5412 49176 5468
rect 49112 5408 49176 5412
rect 49192 5468 49256 5472
rect 49192 5412 49196 5468
rect 49196 5412 49252 5468
rect 49252 5412 49256 5468
rect 49192 5408 49256 5412
rect 49272 5468 49336 5472
rect 49272 5412 49276 5468
rect 49276 5412 49332 5468
rect 49332 5412 49336 5468
rect 49272 5408 49336 5412
rect 49352 5468 49416 5472
rect 49352 5412 49356 5468
rect 49356 5412 49412 5468
rect 49412 5412 49416 5468
rect 49352 5408 49416 5412
rect 20216 4924 20280 4928
rect 20216 4868 20220 4924
rect 20220 4868 20276 4924
rect 20276 4868 20280 4924
rect 20216 4864 20280 4868
rect 20296 4924 20360 4928
rect 20296 4868 20300 4924
rect 20300 4868 20356 4924
rect 20356 4868 20360 4924
rect 20296 4864 20360 4868
rect 20376 4924 20440 4928
rect 20376 4868 20380 4924
rect 20380 4868 20436 4924
rect 20436 4868 20440 4924
rect 20376 4864 20440 4868
rect 20456 4924 20520 4928
rect 20456 4868 20460 4924
rect 20460 4868 20516 4924
rect 20516 4868 20520 4924
rect 20456 4864 20520 4868
rect 39480 4924 39544 4928
rect 39480 4868 39484 4924
rect 39484 4868 39540 4924
rect 39540 4868 39544 4924
rect 39480 4864 39544 4868
rect 39560 4924 39624 4928
rect 39560 4868 39564 4924
rect 39564 4868 39620 4924
rect 39620 4868 39624 4924
rect 39560 4864 39624 4868
rect 39640 4924 39704 4928
rect 39640 4868 39644 4924
rect 39644 4868 39700 4924
rect 39700 4868 39704 4924
rect 39640 4864 39704 4868
rect 39720 4924 39784 4928
rect 39720 4868 39724 4924
rect 39724 4868 39780 4924
rect 39780 4868 39784 4924
rect 39720 4864 39784 4868
rect 10584 4380 10648 4384
rect 10584 4324 10588 4380
rect 10588 4324 10644 4380
rect 10644 4324 10648 4380
rect 10584 4320 10648 4324
rect 10664 4380 10728 4384
rect 10664 4324 10668 4380
rect 10668 4324 10724 4380
rect 10724 4324 10728 4380
rect 10664 4320 10728 4324
rect 10744 4380 10808 4384
rect 10744 4324 10748 4380
rect 10748 4324 10804 4380
rect 10804 4324 10808 4380
rect 10744 4320 10808 4324
rect 10824 4380 10888 4384
rect 10824 4324 10828 4380
rect 10828 4324 10884 4380
rect 10884 4324 10888 4380
rect 10824 4320 10888 4324
rect 29848 4380 29912 4384
rect 29848 4324 29852 4380
rect 29852 4324 29908 4380
rect 29908 4324 29912 4380
rect 29848 4320 29912 4324
rect 29928 4380 29992 4384
rect 29928 4324 29932 4380
rect 29932 4324 29988 4380
rect 29988 4324 29992 4380
rect 29928 4320 29992 4324
rect 30008 4380 30072 4384
rect 30008 4324 30012 4380
rect 30012 4324 30068 4380
rect 30068 4324 30072 4380
rect 30008 4320 30072 4324
rect 30088 4380 30152 4384
rect 30088 4324 30092 4380
rect 30092 4324 30148 4380
rect 30148 4324 30152 4380
rect 30088 4320 30152 4324
rect 49112 4380 49176 4384
rect 49112 4324 49116 4380
rect 49116 4324 49172 4380
rect 49172 4324 49176 4380
rect 49112 4320 49176 4324
rect 49192 4380 49256 4384
rect 49192 4324 49196 4380
rect 49196 4324 49252 4380
rect 49252 4324 49256 4380
rect 49192 4320 49256 4324
rect 49272 4380 49336 4384
rect 49272 4324 49276 4380
rect 49276 4324 49332 4380
rect 49332 4324 49336 4380
rect 49272 4320 49336 4324
rect 49352 4380 49416 4384
rect 49352 4324 49356 4380
rect 49356 4324 49412 4380
rect 49412 4324 49416 4380
rect 49352 4320 49416 4324
rect 20216 3836 20280 3840
rect 20216 3780 20220 3836
rect 20220 3780 20276 3836
rect 20276 3780 20280 3836
rect 20216 3776 20280 3780
rect 20296 3836 20360 3840
rect 20296 3780 20300 3836
rect 20300 3780 20356 3836
rect 20356 3780 20360 3836
rect 20296 3776 20360 3780
rect 20376 3836 20440 3840
rect 20376 3780 20380 3836
rect 20380 3780 20436 3836
rect 20436 3780 20440 3836
rect 20376 3776 20440 3780
rect 20456 3836 20520 3840
rect 20456 3780 20460 3836
rect 20460 3780 20516 3836
rect 20516 3780 20520 3836
rect 20456 3776 20520 3780
rect 39480 3836 39544 3840
rect 39480 3780 39484 3836
rect 39484 3780 39540 3836
rect 39540 3780 39544 3836
rect 39480 3776 39544 3780
rect 39560 3836 39624 3840
rect 39560 3780 39564 3836
rect 39564 3780 39620 3836
rect 39620 3780 39624 3836
rect 39560 3776 39624 3780
rect 39640 3836 39704 3840
rect 39640 3780 39644 3836
rect 39644 3780 39700 3836
rect 39700 3780 39704 3836
rect 39640 3776 39704 3780
rect 39720 3836 39784 3840
rect 39720 3780 39724 3836
rect 39724 3780 39780 3836
rect 39780 3780 39784 3836
rect 39720 3776 39784 3780
rect 10584 3292 10648 3296
rect 10584 3236 10588 3292
rect 10588 3236 10644 3292
rect 10644 3236 10648 3292
rect 10584 3232 10648 3236
rect 10664 3292 10728 3296
rect 10664 3236 10668 3292
rect 10668 3236 10724 3292
rect 10724 3236 10728 3292
rect 10664 3232 10728 3236
rect 10744 3292 10808 3296
rect 10744 3236 10748 3292
rect 10748 3236 10804 3292
rect 10804 3236 10808 3292
rect 10744 3232 10808 3236
rect 10824 3292 10888 3296
rect 10824 3236 10828 3292
rect 10828 3236 10884 3292
rect 10884 3236 10888 3292
rect 10824 3232 10888 3236
rect 29848 3292 29912 3296
rect 29848 3236 29852 3292
rect 29852 3236 29908 3292
rect 29908 3236 29912 3292
rect 29848 3232 29912 3236
rect 29928 3292 29992 3296
rect 29928 3236 29932 3292
rect 29932 3236 29988 3292
rect 29988 3236 29992 3292
rect 29928 3232 29992 3236
rect 30008 3292 30072 3296
rect 30008 3236 30012 3292
rect 30012 3236 30068 3292
rect 30068 3236 30072 3292
rect 30008 3232 30072 3236
rect 30088 3292 30152 3296
rect 30088 3236 30092 3292
rect 30092 3236 30148 3292
rect 30148 3236 30152 3292
rect 30088 3232 30152 3236
rect 49112 3292 49176 3296
rect 49112 3236 49116 3292
rect 49116 3236 49172 3292
rect 49172 3236 49176 3292
rect 49112 3232 49176 3236
rect 49192 3292 49256 3296
rect 49192 3236 49196 3292
rect 49196 3236 49252 3292
rect 49252 3236 49256 3292
rect 49192 3232 49256 3236
rect 49272 3292 49336 3296
rect 49272 3236 49276 3292
rect 49276 3236 49332 3292
rect 49332 3236 49336 3292
rect 49272 3232 49336 3236
rect 49352 3292 49416 3296
rect 49352 3236 49356 3292
rect 49356 3236 49412 3292
rect 49412 3236 49416 3292
rect 49352 3232 49416 3236
rect 20216 2748 20280 2752
rect 20216 2692 20220 2748
rect 20220 2692 20276 2748
rect 20276 2692 20280 2748
rect 20216 2688 20280 2692
rect 20296 2748 20360 2752
rect 20296 2692 20300 2748
rect 20300 2692 20356 2748
rect 20356 2692 20360 2748
rect 20296 2688 20360 2692
rect 20376 2748 20440 2752
rect 20376 2692 20380 2748
rect 20380 2692 20436 2748
rect 20436 2692 20440 2748
rect 20376 2688 20440 2692
rect 20456 2748 20520 2752
rect 20456 2692 20460 2748
rect 20460 2692 20516 2748
rect 20516 2692 20520 2748
rect 20456 2688 20520 2692
rect 39480 2748 39544 2752
rect 39480 2692 39484 2748
rect 39484 2692 39540 2748
rect 39540 2692 39544 2748
rect 39480 2688 39544 2692
rect 39560 2748 39624 2752
rect 39560 2692 39564 2748
rect 39564 2692 39620 2748
rect 39620 2692 39624 2748
rect 39560 2688 39624 2692
rect 39640 2748 39704 2752
rect 39640 2692 39644 2748
rect 39644 2692 39700 2748
rect 39700 2692 39704 2748
rect 39640 2688 39704 2692
rect 39720 2748 39784 2752
rect 39720 2692 39724 2748
rect 39724 2692 39780 2748
rect 39780 2692 39784 2748
rect 39720 2688 39784 2692
rect 10584 2204 10648 2208
rect 10584 2148 10588 2204
rect 10588 2148 10644 2204
rect 10644 2148 10648 2204
rect 10584 2144 10648 2148
rect 10664 2204 10728 2208
rect 10664 2148 10668 2204
rect 10668 2148 10724 2204
rect 10724 2148 10728 2204
rect 10664 2144 10728 2148
rect 10744 2204 10808 2208
rect 10744 2148 10748 2204
rect 10748 2148 10804 2204
rect 10804 2148 10808 2204
rect 10744 2144 10808 2148
rect 10824 2204 10888 2208
rect 10824 2148 10828 2204
rect 10828 2148 10884 2204
rect 10884 2148 10888 2204
rect 10824 2144 10888 2148
rect 29848 2204 29912 2208
rect 29848 2148 29852 2204
rect 29852 2148 29908 2204
rect 29908 2148 29912 2204
rect 29848 2144 29912 2148
rect 29928 2204 29992 2208
rect 29928 2148 29932 2204
rect 29932 2148 29988 2204
rect 29988 2148 29992 2204
rect 29928 2144 29992 2148
rect 30008 2204 30072 2208
rect 30008 2148 30012 2204
rect 30012 2148 30068 2204
rect 30068 2148 30072 2204
rect 30008 2144 30072 2148
rect 30088 2204 30152 2208
rect 30088 2148 30092 2204
rect 30092 2148 30148 2204
rect 30148 2148 30152 2204
rect 30088 2144 30152 2148
rect 49112 2204 49176 2208
rect 49112 2148 49116 2204
rect 49116 2148 49172 2204
rect 49172 2148 49176 2204
rect 49112 2144 49176 2148
rect 49192 2204 49256 2208
rect 49192 2148 49196 2204
rect 49196 2148 49252 2204
rect 49252 2148 49256 2204
rect 49192 2144 49256 2148
rect 49272 2204 49336 2208
rect 49272 2148 49276 2204
rect 49276 2148 49332 2204
rect 49332 2148 49336 2204
rect 49272 2144 49336 2148
rect 49352 2204 49416 2208
rect 49352 2148 49356 2204
rect 49356 2148 49412 2204
rect 49412 2148 49416 2204
rect 49352 2144 49416 2148
<< metal4 >>
rect 10576 27232 10896 27792
rect 10576 27168 10584 27232
rect 10648 27168 10664 27232
rect 10728 27168 10744 27232
rect 10808 27168 10824 27232
rect 10888 27168 10896 27232
rect 10576 26144 10896 27168
rect 10576 26080 10584 26144
rect 10648 26080 10664 26144
rect 10728 26080 10744 26144
rect 10808 26080 10824 26144
rect 10888 26080 10896 26144
rect 10576 25056 10896 26080
rect 10576 24992 10584 25056
rect 10648 24992 10664 25056
rect 10728 24992 10744 25056
rect 10808 24992 10824 25056
rect 10888 24992 10896 25056
rect 10576 23968 10896 24992
rect 10576 23904 10584 23968
rect 10648 23904 10664 23968
rect 10728 23904 10744 23968
rect 10808 23904 10824 23968
rect 10888 23904 10896 23968
rect 10576 23619 10896 23904
rect 10576 23383 10618 23619
rect 10854 23383 10896 23619
rect 10576 22880 10896 23383
rect 10576 22816 10584 22880
rect 10648 22816 10664 22880
rect 10728 22816 10744 22880
rect 10808 22816 10824 22880
rect 10888 22816 10896 22880
rect 10576 21792 10896 22816
rect 10576 21728 10584 21792
rect 10648 21728 10664 21792
rect 10728 21728 10744 21792
rect 10808 21728 10824 21792
rect 10888 21728 10896 21792
rect 10576 20704 10896 21728
rect 10576 20640 10584 20704
rect 10648 20640 10664 20704
rect 10728 20640 10744 20704
rect 10808 20640 10824 20704
rect 10888 20640 10896 20704
rect 10576 19616 10896 20640
rect 10576 19552 10584 19616
rect 10648 19552 10664 19616
rect 10728 19552 10744 19616
rect 10808 19552 10824 19616
rect 10888 19552 10896 19616
rect 10576 18528 10896 19552
rect 10576 18464 10584 18528
rect 10648 18464 10664 18528
rect 10728 18464 10744 18528
rect 10808 18464 10824 18528
rect 10888 18464 10896 18528
rect 10576 17440 10896 18464
rect 10576 17376 10584 17440
rect 10648 17376 10664 17440
rect 10728 17376 10744 17440
rect 10808 17376 10824 17440
rect 10888 17376 10896 17440
rect 10576 16352 10896 17376
rect 10576 16288 10584 16352
rect 10648 16288 10664 16352
rect 10728 16288 10744 16352
rect 10808 16288 10824 16352
rect 10888 16288 10896 16352
rect 10576 15264 10896 16288
rect 10576 15200 10584 15264
rect 10648 15200 10664 15264
rect 10728 15200 10744 15264
rect 10808 15200 10824 15264
rect 10888 15200 10896 15264
rect 10576 15070 10896 15200
rect 10576 14834 10618 15070
rect 10854 14834 10896 15070
rect 10576 14176 10896 14834
rect 10576 14112 10584 14176
rect 10648 14112 10664 14176
rect 10728 14112 10744 14176
rect 10808 14112 10824 14176
rect 10888 14112 10896 14176
rect 10576 13088 10896 14112
rect 10576 13024 10584 13088
rect 10648 13024 10664 13088
rect 10728 13024 10744 13088
rect 10808 13024 10824 13088
rect 10888 13024 10896 13088
rect 10576 12000 10896 13024
rect 10576 11936 10584 12000
rect 10648 11936 10664 12000
rect 10728 11936 10744 12000
rect 10808 11936 10824 12000
rect 10888 11936 10896 12000
rect 10576 10912 10896 11936
rect 10576 10848 10584 10912
rect 10648 10848 10664 10912
rect 10728 10848 10744 10912
rect 10808 10848 10824 10912
rect 10888 10848 10896 10912
rect 10576 9824 10896 10848
rect 10576 9760 10584 9824
rect 10648 9760 10664 9824
rect 10728 9760 10744 9824
rect 10808 9760 10824 9824
rect 10888 9760 10896 9824
rect 10576 8736 10896 9760
rect 10576 8672 10584 8736
rect 10648 8672 10664 8736
rect 10728 8672 10744 8736
rect 10808 8672 10824 8736
rect 10888 8672 10896 8736
rect 10576 7648 10896 8672
rect 10576 7584 10584 7648
rect 10648 7584 10664 7648
rect 10728 7584 10744 7648
rect 10808 7584 10824 7648
rect 10888 7584 10896 7648
rect 10576 6560 10896 7584
rect 10576 6496 10584 6560
rect 10648 6520 10664 6560
rect 10728 6520 10744 6560
rect 10808 6520 10824 6560
rect 10888 6496 10896 6560
rect 10576 6284 10618 6496
rect 10854 6284 10896 6496
rect 10576 5472 10896 6284
rect 10576 5408 10584 5472
rect 10648 5408 10664 5472
rect 10728 5408 10744 5472
rect 10808 5408 10824 5472
rect 10888 5408 10896 5472
rect 10576 4384 10896 5408
rect 10576 4320 10584 4384
rect 10648 4320 10664 4384
rect 10728 4320 10744 4384
rect 10808 4320 10824 4384
rect 10888 4320 10896 4384
rect 10576 3296 10896 4320
rect 10576 3232 10584 3296
rect 10648 3232 10664 3296
rect 10728 3232 10744 3296
rect 10808 3232 10824 3296
rect 10888 3232 10896 3296
rect 10576 2208 10896 3232
rect 10576 2144 10584 2208
rect 10648 2144 10664 2208
rect 10728 2144 10744 2208
rect 10808 2144 10824 2208
rect 10888 2144 10896 2208
rect 10576 2128 10896 2144
rect 20208 27776 20528 27792
rect 20208 27712 20216 27776
rect 20280 27712 20296 27776
rect 20360 27712 20376 27776
rect 20440 27712 20456 27776
rect 20520 27712 20528 27776
rect 20208 26688 20528 27712
rect 20208 26624 20216 26688
rect 20280 26624 20296 26688
rect 20360 26624 20376 26688
rect 20440 26624 20456 26688
rect 20520 26624 20528 26688
rect 20208 25600 20528 26624
rect 20208 25536 20216 25600
rect 20280 25536 20296 25600
rect 20360 25536 20376 25600
rect 20440 25536 20456 25600
rect 20520 25536 20528 25600
rect 20208 24512 20528 25536
rect 20208 24448 20216 24512
rect 20280 24448 20296 24512
rect 20360 24448 20376 24512
rect 20440 24448 20456 24512
rect 20520 24448 20528 24512
rect 20208 23424 20528 24448
rect 20208 23360 20216 23424
rect 20280 23360 20296 23424
rect 20360 23360 20376 23424
rect 20440 23360 20456 23424
rect 20520 23360 20528 23424
rect 20208 22336 20528 23360
rect 20208 22272 20216 22336
rect 20280 22272 20296 22336
rect 20360 22272 20376 22336
rect 20440 22272 20456 22336
rect 20520 22272 20528 22336
rect 20208 21248 20528 22272
rect 20208 21184 20216 21248
rect 20280 21184 20296 21248
rect 20360 21184 20376 21248
rect 20440 21184 20456 21248
rect 20520 21184 20528 21248
rect 20208 20160 20528 21184
rect 20208 20096 20216 20160
rect 20280 20096 20296 20160
rect 20360 20096 20376 20160
rect 20440 20096 20456 20160
rect 20520 20096 20528 20160
rect 20208 19344 20528 20096
rect 20208 19108 20250 19344
rect 20486 19108 20528 19344
rect 20208 19072 20528 19108
rect 20208 19008 20216 19072
rect 20280 19008 20296 19072
rect 20360 19008 20376 19072
rect 20440 19008 20456 19072
rect 20520 19008 20528 19072
rect 20208 17984 20528 19008
rect 20208 17920 20216 17984
rect 20280 17920 20296 17984
rect 20360 17920 20376 17984
rect 20440 17920 20456 17984
rect 20520 17920 20528 17984
rect 20208 16896 20528 17920
rect 20208 16832 20216 16896
rect 20280 16832 20296 16896
rect 20360 16832 20376 16896
rect 20440 16832 20456 16896
rect 20520 16832 20528 16896
rect 20208 15808 20528 16832
rect 20208 15744 20216 15808
rect 20280 15744 20296 15808
rect 20360 15744 20376 15808
rect 20440 15744 20456 15808
rect 20520 15744 20528 15808
rect 20208 14720 20528 15744
rect 20208 14656 20216 14720
rect 20280 14656 20296 14720
rect 20360 14656 20376 14720
rect 20440 14656 20456 14720
rect 20520 14656 20528 14720
rect 20208 13632 20528 14656
rect 20208 13568 20216 13632
rect 20280 13568 20296 13632
rect 20360 13568 20376 13632
rect 20440 13568 20456 13632
rect 20520 13568 20528 13632
rect 20208 12544 20528 13568
rect 20208 12480 20216 12544
rect 20280 12480 20296 12544
rect 20360 12480 20376 12544
rect 20440 12480 20456 12544
rect 20520 12480 20528 12544
rect 20208 11456 20528 12480
rect 20208 11392 20216 11456
rect 20280 11392 20296 11456
rect 20360 11392 20376 11456
rect 20440 11392 20456 11456
rect 20520 11392 20528 11456
rect 20208 10795 20528 11392
rect 20208 10559 20250 10795
rect 20486 10559 20528 10795
rect 20208 10368 20528 10559
rect 20208 10304 20216 10368
rect 20280 10304 20296 10368
rect 20360 10304 20376 10368
rect 20440 10304 20456 10368
rect 20520 10304 20528 10368
rect 20208 9280 20528 10304
rect 20208 9216 20216 9280
rect 20280 9216 20296 9280
rect 20360 9216 20376 9280
rect 20440 9216 20456 9280
rect 20520 9216 20528 9280
rect 20208 8192 20528 9216
rect 20208 8128 20216 8192
rect 20280 8128 20296 8192
rect 20360 8128 20376 8192
rect 20440 8128 20456 8192
rect 20520 8128 20528 8192
rect 20208 7104 20528 8128
rect 20208 7040 20216 7104
rect 20280 7040 20296 7104
rect 20360 7040 20376 7104
rect 20440 7040 20456 7104
rect 20520 7040 20528 7104
rect 20208 6016 20528 7040
rect 20208 5952 20216 6016
rect 20280 5952 20296 6016
rect 20360 5952 20376 6016
rect 20440 5952 20456 6016
rect 20520 5952 20528 6016
rect 20208 4928 20528 5952
rect 20208 4864 20216 4928
rect 20280 4864 20296 4928
rect 20360 4864 20376 4928
rect 20440 4864 20456 4928
rect 20520 4864 20528 4928
rect 20208 3840 20528 4864
rect 20208 3776 20216 3840
rect 20280 3776 20296 3840
rect 20360 3776 20376 3840
rect 20440 3776 20456 3840
rect 20520 3776 20528 3840
rect 20208 2752 20528 3776
rect 20208 2688 20216 2752
rect 20280 2688 20296 2752
rect 20360 2688 20376 2752
rect 20440 2688 20456 2752
rect 20520 2688 20528 2752
rect 20208 2128 20528 2688
rect 29840 27232 30160 27792
rect 29840 27168 29848 27232
rect 29912 27168 29928 27232
rect 29992 27168 30008 27232
rect 30072 27168 30088 27232
rect 30152 27168 30160 27232
rect 29840 26144 30160 27168
rect 29840 26080 29848 26144
rect 29912 26080 29928 26144
rect 29992 26080 30008 26144
rect 30072 26080 30088 26144
rect 30152 26080 30160 26144
rect 29840 25056 30160 26080
rect 29840 24992 29848 25056
rect 29912 24992 29928 25056
rect 29992 24992 30008 25056
rect 30072 24992 30088 25056
rect 30152 24992 30160 25056
rect 29840 23968 30160 24992
rect 29840 23904 29848 23968
rect 29912 23904 29928 23968
rect 29992 23904 30008 23968
rect 30072 23904 30088 23968
rect 30152 23904 30160 23968
rect 29840 23619 30160 23904
rect 29840 23383 29882 23619
rect 30118 23383 30160 23619
rect 29840 22880 30160 23383
rect 29840 22816 29848 22880
rect 29912 22816 29928 22880
rect 29992 22816 30008 22880
rect 30072 22816 30088 22880
rect 30152 22816 30160 22880
rect 29840 21792 30160 22816
rect 29840 21728 29848 21792
rect 29912 21728 29928 21792
rect 29992 21728 30008 21792
rect 30072 21728 30088 21792
rect 30152 21728 30160 21792
rect 29840 20704 30160 21728
rect 29840 20640 29848 20704
rect 29912 20640 29928 20704
rect 29992 20640 30008 20704
rect 30072 20640 30088 20704
rect 30152 20640 30160 20704
rect 29840 19616 30160 20640
rect 29840 19552 29848 19616
rect 29912 19552 29928 19616
rect 29992 19552 30008 19616
rect 30072 19552 30088 19616
rect 30152 19552 30160 19616
rect 29840 18528 30160 19552
rect 29840 18464 29848 18528
rect 29912 18464 29928 18528
rect 29992 18464 30008 18528
rect 30072 18464 30088 18528
rect 30152 18464 30160 18528
rect 29840 17440 30160 18464
rect 29840 17376 29848 17440
rect 29912 17376 29928 17440
rect 29992 17376 30008 17440
rect 30072 17376 30088 17440
rect 30152 17376 30160 17440
rect 29840 16352 30160 17376
rect 29840 16288 29848 16352
rect 29912 16288 29928 16352
rect 29992 16288 30008 16352
rect 30072 16288 30088 16352
rect 30152 16288 30160 16352
rect 29840 15264 30160 16288
rect 29840 15200 29848 15264
rect 29912 15200 29928 15264
rect 29992 15200 30008 15264
rect 30072 15200 30088 15264
rect 30152 15200 30160 15264
rect 29840 15070 30160 15200
rect 29840 14834 29882 15070
rect 30118 14834 30160 15070
rect 29840 14176 30160 14834
rect 29840 14112 29848 14176
rect 29912 14112 29928 14176
rect 29992 14112 30008 14176
rect 30072 14112 30088 14176
rect 30152 14112 30160 14176
rect 29840 13088 30160 14112
rect 29840 13024 29848 13088
rect 29912 13024 29928 13088
rect 29992 13024 30008 13088
rect 30072 13024 30088 13088
rect 30152 13024 30160 13088
rect 29840 12000 30160 13024
rect 29840 11936 29848 12000
rect 29912 11936 29928 12000
rect 29992 11936 30008 12000
rect 30072 11936 30088 12000
rect 30152 11936 30160 12000
rect 29840 10912 30160 11936
rect 29840 10848 29848 10912
rect 29912 10848 29928 10912
rect 29992 10848 30008 10912
rect 30072 10848 30088 10912
rect 30152 10848 30160 10912
rect 29840 9824 30160 10848
rect 29840 9760 29848 9824
rect 29912 9760 29928 9824
rect 29992 9760 30008 9824
rect 30072 9760 30088 9824
rect 30152 9760 30160 9824
rect 29840 8736 30160 9760
rect 29840 8672 29848 8736
rect 29912 8672 29928 8736
rect 29992 8672 30008 8736
rect 30072 8672 30088 8736
rect 30152 8672 30160 8736
rect 29840 7648 30160 8672
rect 29840 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30160 7648
rect 29840 6560 30160 7584
rect 29840 6496 29848 6560
rect 29912 6520 29928 6560
rect 29992 6520 30008 6560
rect 30072 6520 30088 6560
rect 30152 6496 30160 6560
rect 29840 6284 29882 6496
rect 30118 6284 30160 6496
rect 29840 5472 30160 6284
rect 29840 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30160 5472
rect 29840 4384 30160 5408
rect 29840 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30160 4384
rect 29840 3296 30160 4320
rect 29840 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30160 3296
rect 29840 2208 30160 3232
rect 29840 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30160 2208
rect 29840 2128 30160 2144
rect 39472 27776 39792 27792
rect 39472 27712 39480 27776
rect 39544 27712 39560 27776
rect 39624 27712 39640 27776
rect 39704 27712 39720 27776
rect 39784 27712 39792 27776
rect 39472 26688 39792 27712
rect 39472 26624 39480 26688
rect 39544 26624 39560 26688
rect 39624 26624 39640 26688
rect 39704 26624 39720 26688
rect 39784 26624 39792 26688
rect 39472 25600 39792 26624
rect 39472 25536 39480 25600
rect 39544 25536 39560 25600
rect 39624 25536 39640 25600
rect 39704 25536 39720 25600
rect 39784 25536 39792 25600
rect 39472 24512 39792 25536
rect 39472 24448 39480 24512
rect 39544 24448 39560 24512
rect 39624 24448 39640 24512
rect 39704 24448 39720 24512
rect 39784 24448 39792 24512
rect 39472 23424 39792 24448
rect 39472 23360 39480 23424
rect 39544 23360 39560 23424
rect 39624 23360 39640 23424
rect 39704 23360 39720 23424
rect 39784 23360 39792 23424
rect 39472 22336 39792 23360
rect 39472 22272 39480 22336
rect 39544 22272 39560 22336
rect 39624 22272 39640 22336
rect 39704 22272 39720 22336
rect 39784 22272 39792 22336
rect 39472 21248 39792 22272
rect 39472 21184 39480 21248
rect 39544 21184 39560 21248
rect 39624 21184 39640 21248
rect 39704 21184 39720 21248
rect 39784 21184 39792 21248
rect 39472 20160 39792 21184
rect 39472 20096 39480 20160
rect 39544 20096 39560 20160
rect 39624 20096 39640 20160
rect 39704 20096 39720 20160
rect 39784 20096 39792 20160
rect 39472 19344 39792 20096
rect 39472 19108 39514 19344
rect 39750 19108 39792 19344
rect 39472 19072 39792 19108
rect 39472 19008 39480 19072
rect 39544 19008 39560 19072
rect 39624 19008 39640 19072
rect 39704 19008 39720 19072
rect 39784 19008 39792 19072
rect 39472 17984 39792 19008
rect 39472 17920 39480 17984
rect 39544 17920 39560 17984
rect 39624 17920 39640 17984
rect 39704 17920 39720 17984
rect 39784 17920 39792 17984
rect 39472 16896 39792 17920
rect 39472 16832 39480 16896
rect 39544 16832 39560 16896
rect 39624 16832 39640 16896
rect 39704 16832 39720 16896
rect 39784 16832 39792 16896
rect 39472 15808 39792 16832
rect 39472 15744 39480 15808
rect 39544 15744 39560 15808
rect 39624 15744 39640 15808
rect 39704 15744 39720 15808
rect 39784 15744 39792 15808
rect 39472 14720 39792 15744
rect 39472 14656 39480 14720
rect 39544 14656 39560 14720
rect 39624 14656 39640 14720
rect 39704 14656 39720 14720
rect 39784 14656 39792 14720
rect 39472 13632 39792 14656
rect 39472 13568 39480 13632
rect 39544 13568 39560 13632
rect 39624 13568 39640 13632
rect 39704 13568 39720 13632
rect 39784 13568 39792 13632
rect 39472 12544 39792 13568
rect 39472 12480 39480 12544
rect 39544 12480 39560 12544
rect 39624 12480 39640 12544
rect 39704 12480 39720 12544
rect 39784 12480 39792 12544
rect 39472 11456 39792 12480
rect 39472 11392 39480 11456
rect 39544 11392 39560 11456
rect 39624 11392 39640 11456
rect 39704 11392 39720 11456
rect 39784 11392 39792 11456
rect 39472 10795 39792 11392
rect 39472 10559 39514 10795
rect 39750 10559 39792 10795
rect 39472 10368 39792 10559
rect 39472 10304 39480 10368
rect 39544 10304 39560 10368
rect 39624 10304 39640 10368
rect 39704 10304 39720 10368
rect 39784 10304 39792 10368
rect 39472 9280 39792 10304
rect 39472 9216 39480 9280
rect 39544 9216 39560 9280
rect 39624 9216 39640 9280
rect 39704 9216 39720 9280
rect 39784 9216 39792 9280
rect 39472 8192 39792 9216
rect 39472 8128 39480 8192
rect 39544 8128 39560 8192
rect 39624 8128 39640 8192
rect 39704 8128 39720 8192
rect 39784 8128 39792 8192
rect 39472 7104 39792 8128
rect 39472 7040 39480 7104
rect 39544 7040 39560 7104
rect 39624 7040 39640 7104
rect 39704 7040 39720 7104
rect 39784 7040 39792 7104
rect 39472 6016 39792 7040
rect 39472 5952 39480 6016
rect 39544 5952 39560 6016
rect 39624 5952 39640 6016
rect 39704 5952 39720 6016
rect 39784 5952 39792 6016
rect 39472 4928 39792 5952
rect 39472 4864 39480 4928
rect 39544 4864 39560 4928
rect 39624 4864 39640 4928
rect 39704 4864 39720 4928
rect 39784 4864 39792 4928
rect 39472 3840 39792 4864
rect 39472 3776 39480 3840
rect 39544 3776 39560 3840
rect 39624 3776 39640 3840
rect 39704 3776 39720 3840
rect 39784 3776 39792 3840
rect 39472 2752 39792 3776
rect 39472 2688 39480 2752
rect 39544 2688 39560 2752
rect 39624 2688 39640 2752
rect 39704 2688 39720 2752
rect 39784 2688 39792 2752
rect 39472 2128 39792 2688
rect 49104 27232 49424 27792
rect 49104 27168 49112 27232
rect 49176 27168 49192 27232
rect 49256 27168 49272 27232
rect 49336 27168 49352 27232
rect 49416 27168 49424 27232
rect 49104 26144 49424 27168
rect 49104 26080 49112 26144
rect 49176 26080 49192 26144
rect 49256 26080 49272 26144
rect 49336 26080 49352 26144
rect 49416 26080 49424 26144
rect 49104 25056 49424 26080
rect 49104 24992 49112 25056
rect 49176 24992 49192 25056
rect 49256 24992 49272 25056
rect 49336 24992 49352 25056
rect 49416 24992 49424 25056
rect 49104 23968 49424 24992
rect 49104 23904 49112 23968
rect 49176 23904 49192 23968
rect 49256 23904 49272 23968
rect 49336 23904 49352 23968
rect 49416 23904 49424 23968
rect 49104 23619 49424 23904
rect 49104 23383 49146 23619
rect 49382 23383 49424 23619
rect 49104 22880 49424 23383
rect 49104 22816 49112 22880
rect 49176 22816 49192 22880
rect 49256 22816 49272 22880
rect 49336 22816 49352 22880
rect 49416 22816 49424 22880
rect 49104 21792 49424 22816
rect 49104 21728 49112 21792
rect 49176 21728 49192 21792
rect 49256 21728 49272 21792
rect 49336 21728 49352 21792
rect 49416 21728 49424 21792
rect 49104 20704 49424 21728
rect 49104 20640 49112 20704
rect 49176 20640 49192 20704
rect 49256 20640 49272 20704
rect 49336 20640 49352 20704
rect 49416 20640 49424 20704
rect 49104 19616 49424 20640
rect 49104 19552 49112 19616
rect 49176 19552 49192 19616
rect 49256 19552 49272 19616
rect 49336 19552 49352 19616
rect 49416 19552 49424 19616
rect 49104 18528 49424 19552
rect 49104 18464 49112 18528
rect 49176 18464 49192 18528
rect 49256 18464 49272 18528
rect 49336 18464 49352 18528
rect 49416 18464 49424 18528
rect 49104 17440 49424 18464
rect 49104 17376 49112 17440
rect 49176 17376 49192 17440
rect 49256 17376 49272 17440
rect 49336 17376 49352 17440
rect 49416 17376 49424 17440
rect 49104 16352 49424 17376
rect 49104 16288 49112 16352
rect 49176 16288 49192 16352
rect 49256 16288 49272 16352
rect 49336 16288 49352 16352
rect 49416 16288 49424 16352
rect 49104 15264 49424 16288
rect 49104 15200 49112 15264
rect 49176 15200 49192 15264
rect 49256 15200 49272 15264
rect 49336 15200 49352 15264
rect 49416 15200 49424 15264
rect 49104 15070 49424 15200
rect 49104 14834 49146 15070
rect 49382 14834 49424 15070
rect 49104 14176 49424 14834
rect 49104 14112 49112 14176
rect 49176 14112 49192 14176
rect 49256 14112 49272 14176
rect 49336 14112 49352 14176
rect 49416 14112 49424 14176
rect 49104 13088 49424 14112
rect 49104 13024 49112 13088
rect 49176 13024 49192 13088
rect 49256 13024 49272 13088
rect 49336 13024 49352 13088
rect 49416 13024 49424 13088
rect 49104 12000 49424 13024
rect 49104 11936 49112 12000
rect 49176 11936 49192 12000
rect 49256 11936 49272 12000
rect 49336 11936 49352 12000
rect 49416 11936 49424 12000
rect 49104 10912 49424 11936
rect 49104 10848 49112 10912
rect 49176 10848 49192 10912
rect 49256 10848 49272 10912
rect 49336 10848 49352 10912
rect 49416 10848 49424 10912
rect 49104 9824 49424 10848
rect 49104 9760 49112 9824
rect 49176 9760 49192 9824
rect 49256 9760 49272 9824
rect 49336 9760 49352 9824
rect 49416 9760 49424 9824
rect 49104 8736 49424 9760
rect 49104 8672 49112 8736
rect 49176 8672 49192 8736
rect 49256 8672 49272 8736
rect 49336 8672 49352 8736
rect 49416 8672 49424 8736
rect 49104 7648 49424 8672
rect 49104 7584 49112 7648
rect 49176 7584 49192 7648
rect 49256 7584 49272 7648
rect 49336 7584 49352 7648
rect 49416 7584 49424 7648
rect 49104 6560 49424 7584
rect 49104 6496 49112 6560
rect 49176 6520 49192 6560
rect 49256 6520 49272 6560
rect 49336 6520 49352 6560
rect 49416 6496 49424 6560
rect 49104 6284 49146 6496
rect 49382 6284 49424 6496
rect 49104 5472 49424 6284
rect 49104 5408 49112 5472
rect 49176 5408 49192 5472
rect 49256 5408 49272 5472
rect 49336 5408 49352 5472
rect 49416 5408 49424 5472
rect 49104 4384 49424 5408
rect 49104 4320 49112 4384
rect 49176 4320 49192 4384
rect 49256 4320 49272 4384
rect 49336 4320 49352 4384
rect 49416 4320 49424 4384
rect 49104 3296 49424 4320
rect 49104 3232 49112 3296
rect 49176 3232 49192 3296
rect 49256 3232 49272 3296
rect 49336 3232 49352 3296
rect 49416 3232 49424 3296
rect 49104 2208 49424 3232
rect 49104 2144 49112 2208
rect 49176 2144 49192 2208
rect 49256 2144 49272 2208
rect 49336 2144 49352 2208
rect 49416 2144 49424 2208
rect 49104 2128 49424 2144
<< via4 >>
rect 10618 23383 10854 23619
rect 10618 14834 10854 15070
rect 10618 6496 10648 6520
rect 10648 6496 10664 6520
rect 10664 6496 10728 6520
rect 10728 6496 10744 6520
rect 10744 6496 10808 6520
rect 10808 6496 10824 6520
rect 10824 6496 10854 6520
rect 10618 6284 10854 6496
rect 20250 19108 20486 19344
rect 20250 10559 20486 10795
rect 29882 23383 30118 23619
rect 29882 14834 30118 15070
rect 29882 6496 29912 6520
rect 29912 6496 29928 6520
rect 29928 6496 29992 6520
rect 29992 6496 30008 6520
rect 30008 6496 30072 6520
rect 30072 6496 30088 6520
rect 30088 6496 30118 6520
rect 29882 6284 30118 6496
rect 39514 19108 39750 19344
rect 39514 10559 39750 10795
rect 49146 23383 49382 23619
rect 49146 14834 49382 15070
rect 49146 6496 49176 6520
rect 49176 6496 49192 6520
rect 49192 6496 49256 6520
rect 49256 6496 49272 6520
rect 49272 6496 49336 6520
rect 49336 6496 49352 6520
rect 49352 6496 49382 6520
rect 49146 6284 49382 6496
<< metal5 >>
rect 1104 23619 58880 23661
rect 1104 23383 10618 23619
rect 10854 23383 29882 23619
rect 30118 23383 49146 23619
rect 49382 23383 58880 23619
rect 1104 23341 58880 23383
rect 1104 19344 58880 19387
rect 1104 19108 20250 19344
rect 20486 19108 39514 19344
rect 39750 19108 58880 19344
rect 1104 19066 58880 19108
rect 1104 15070 58880 15112
rect 1104 14834 10618 15070
rect 10854 14834 29882 15070
rect 30118 14834 49146 15070
rect 49382 14834 58880 15070
rect 1104 14792 58880 14834
rect 1104 10795 58880 10837
rect 1104 10559 20250 10795
rect 20486 10559 39514 10795
rect 39750 10559 58880 10795
rect 1104 10517 58880 10559
rect 1104 6520 58880 6563
rect 1104 6284 10618 6520
rect 10854 6284 29882 6520
rect 30118 6284 49146 6520
rect 49382 6284 58880 6520
rect 1104 6242 58880 6284
use sky130_fd_sc_hd__decap_3  PHY_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1624047346
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 2208 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output165 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 2208 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 1656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_14
timestamp 1624047346
transform 1 0 2392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1624047346
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25
timestamp 1624047346
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 2944 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output133
timestamp 1624047346
transform -1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1624047346
transform 1 0 3036 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_32
timestamp 1624047346
transform 1 0 4048 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1624047346
transform 1 0 3680 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624047346
transform -1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output154
timestamp 1624047346
transform -1 0 4508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32
timestamp 1624047346
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1624047346
transform 1 0 5520 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1624047346
transform 1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output239
timestamp 1624047346
transform -1 0 5244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output239_A
timestamp 1624047346
transform -1 0 5796 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44
timestamp 1624047346
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_37
timestamp 1624047346
transform 1 0 4508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_45
timestamp 1624047346
transform 1 0 5244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 5796 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52
timestamp 1624047346
transform 1 0 5888 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624047346
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_58
timestamp 1624047346
transform 1 0 6440 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61
timestamp 1624047346
transform 1 0 6716 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624047346
transform -1 0 6716 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  input101 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 6808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624047346
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_66
timestamp 1624047346
transform 1 0 7176 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1624047346
transform 1 0 7268 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1624047346
transform 1 0 7360 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 1624047346
transform -1 0 9016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output171
timestamp 1624047346
transform -1 0 8464 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624047346
transform -1 0 7912 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1624047346
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80
timestamp 1624047346
transform 1 0 8464 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1624047346
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_82
timestamp 1624047346
transform 1 0 8648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_86
timestamp 1624047346
transform 1 0 9016 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1624047346
transform 1 0 9384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86
timestamp 1624047346
transform 1 0 9016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1624047346
transform -1 0 9384 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624047346
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1624047346
transform 1 0 9936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92
timestamp 1624047346
transform 1 0 9568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1624047346
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output180
timestamp 1624047346
transform 1 0 9844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input55 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 9660 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99
timestamp 1624047346
transform 1 0 10212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624047346
transform -1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1624047346
transform 1 0 10488 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output237
timestamp 1624047346
transform -1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1624047346
transform 1 0 10580 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1624047346
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1624047346
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1624047346
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_115
timestamp 1624047346
transform 1 0 11684 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624047346
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624047346
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107
timestamp 1624047346
transform 1 0 10948 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1624047346
transform 1 0 12236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output172
timestamp 1624047346
transform 1 0 12972 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output187
timestamp 1624047346
transform -1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624047346
transform -1 0 12236 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1624047346
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_133
timestamp 1624047346
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_121
timestamp 1624047346
transform 1 0 12236 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1624047346
transform 1 0 12788 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_132
timestamp 1624047346
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_139
timestamp 1624047346
transform 1 0 13892 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_136
timestamp 1624047346
transform 1 0 13616 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1624047346
transform 1 0 14076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__S
timestamp 1624047346
transform 1 0 13708 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output213
timestamp 1624047346
transform -1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1624047346
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_146
timestamp 1624047346
transform 1 0 14536 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624047346
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_147
timestamp 1624047346
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _252_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 14904 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _097_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _210_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 16744 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  output201
timestamp 1624047346
transform -1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_159
timestamp 1624047346
transform 1 0 15732 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1624047346
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_162
timestamp 1624047346
transform 1 0 16008 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_167
timestamp 1624047346
transform 1 0 16468 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_8  _119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 19228 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_2  _277_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 17572 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624047346
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624047346
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624047346
transform -1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_170
timestamp 1624047346
transform 1 0 16744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1624047346
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_172
timestamp 1624047346
transform 1 0 16928 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_175
timestamp 1624047346
transform 1 0 17204 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624047346
transform 1 0 19596 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output176
timestamp 1624047346
transform -1 0 19228 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_188
timestamp 1624047346
transform 1 0 18400 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_192
timestamp 1624047346
transform 1 0 18768 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 1624047346
transform 1 0 19228 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1624047346
transform 1 0 19228 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624047346
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1624047346
transform -1 0 20976 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output160
timestamp 1624047346
transform -1 0 20608 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_204
timestamp 1624047346
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_212
timestamp 1624047346
transform 1 0 20608 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_218
timestamp 1624047346
transform 1 0 21160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_204
timestamp 1624047346
transform 1 0 19872 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_212
timestamp 1624047346
transform 1 0 20608 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_216
timestamp 1624047346
transform 1 0 20976 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _262_
timestamp 1624047346
transform 1 0 21252 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624047346
transform 1 0 22448 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624047346
transform 1 0 22080 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1624047346
transform 1 0 22540 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624047346
transform -1 0 21712 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_228
timestamp 1624047346
transform 1 0 22080 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_233
timestamp 1624047346
transform 1 0 22540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_224
timestamp 1624047346
transform 1 0 21712 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1624047346
transform 1 0 22172 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_244
timestamp 1624047346
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_241
timestamp 1624047346
transform 1 0 23276 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output149
timestamp 1624047346
transform -1 0 23276 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1624047346
transform 1 0 23920 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1624047346
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output219
timestamp 1624047346
transform 1 0 24288 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output147
timestamp 1624047346
transform -1 0 24288 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _124_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 23644 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_236
timestamp 1624047346
transform 1 0 22816 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_252
timestamp 1624047346
transform 1 0 24288 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _125_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 26588 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624047346
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output159
timestamp 1624047346
transform -1 0 26128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output175
timestamp 1624047346
transform 1 0 25024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output147_A
timestamp 1624047346
transform -1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_260
timestamp 1624047346
transform 1 0 25024 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_264
timestamp 1624047346
transform 1 0 25392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_256
timestamp 1624047346
transform 1 0 24656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1624047346
transform 1 0 25392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624047346
transform 1 0 27324 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output150
timestamp 1624047346
transform -1 0 27324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output194
timestamp 1624047346
transform 1 0 26588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_277
timestamp 1624047346
transform 1 0 26588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285
timestamp 1624047346
transform 1 0 27324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_272
timestamp 1624047346
transform 1 0 26128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_276
timestamp 1624047346
transform 1 0 26496 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1624047346
transform 1 0 26956 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1624047346
transform 1 0 27416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1624047346
transform 1 0 27784 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624047346
transform 1 0 27784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1624047346
transform 1 0 28336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 1624047346
transform 1 0 27692 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1624047346
transform 1 0 27876 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_295
timestamp 1624047346
transform 1 0 28244 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_300
timestamp 1624047346
transform 1 0 28704 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_299
timestamp 1624047346
transform 1 0 28612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_303
timestamp 1624047346
transform 1 0 28980 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_8  _091_
timestamp 1624047346
transform 1 0 29072 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _193_
timestamp 1624047346
transform 1 0 29072 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624047346
transform 1 0 30452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_313
timestamp 1624047346
transform 1 0 29900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output142
timestamp 1624047346
transform -1 0 31648 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output193
timestamp 1624047346
transform -1 0 32108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output243
timestamp 1624047346
transform -1 0 31280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624047346
transform -1 0 30728 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_322
timestamp 1624047346
transform 1 0 30728 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_332
timestamp 1624047346
transform 1 0 31648 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_320
timestamp 1624047346
transform 1 0 30544 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_328
timestamp 1624047346
transform 1 0 31280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_332
timestamp 1624047346
transform 1 0 31648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_341
timestamp 1624047346
transform 1 0 32476 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_337
timestamp 1624047346
transform 1 0 32108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output155
timestamp 1624047346
transform 1 0 32384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_343
timestamp 1624047346
transform 1 0 32660 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_344
timestamp 1624047346
transform 1 0 32752 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624047346
transform 1 0 32568 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_349
timestamp 1624047346
transform 1 0 33212 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_349
timestamp 1624047346
transform 1 0 33212 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624047346
transform -1 0 33212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624047346
transform 1 0 33120 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1624047346
transform -1 0 33948 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1624047346
transform 1 0 33580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1624047346
transform 1 0 34592 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _220_
timestamp 1624047346
transform -1 0 35420 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1624047346
transform 1 0 33948 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1624047346
transform 1 0 34500 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_356
timestamp 1624047346
transform 1 0 33856 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_367
timestamp 1624047346
transform 1 0 34868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _102_
timestamp 1624047346
transform 1 0 36248 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_8  _137_
timestamp 1624047346
transform -1 0 37260 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624047346
transform 1 0 35788 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1624047346
transform 1 0 35236 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_373
timestamp 1624047346
transform 1 0 35420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_378
timestamp 1624047346
transform 1 0 35880 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_387
timestamp 1624047346
transform 1 0 36708 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_373
timestamp 1624047346
transform 1 0 35420 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1624047346
transform 1 0 38272 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _150_
timestamp 1624047346
transform 1 0 37260 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624047346
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_402
timestamp 1624047346
transform 1 0 38088 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_393
timestamp 1624047346
transform 1 0 37260 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_400
timestamp 1624047346
transform 1 0 37904 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _222_
timestamp 1624047346
transform 1 0 39744 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624047346
transform 1 0 38456 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output144
timestamp 1624047346
transform -1 0 39284 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output217
timestamp 1624047346
transform 1 0 39008 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_407
timestamp 1624047346
transform 1 0 38548 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_415
timestamp 1624047346
transform 1 0 39284 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_407
timestamp 1624047346
transform 1 0 38548 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_411
timestamp 1624047346
transform 1 0 38916 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_416
timestamp 1624047346
transform 1 0 39376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _265_
timestamp 1624047346
transform 1 0 39928 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _271_
timestamp 1624047346
transform -1 0 41768 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624047346
transform 1 0 41124 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1624047346
transform 1 0 39836 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1624047346
transform 1 0 40756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_436
timestamp 1624047346
transform 1 0 41216 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_429
timestamp 1624047346
transform 1 0 40572 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _141_
timestamp 1624047346
transform 1 0 41584 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _267_
timestamp 1624047346
transform 1 0 42596 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1624047346
transform -1 0 42688 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_445
timestamp 1624047346
transform 1 0 42044 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_442
timestamp 1624047346
transform 1 0 41768 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1624047346
transform 1 0 42688 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _256_
timestamp 1624047346
transform 1 0 43516 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624047346
transform 1 0 43792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624047346
transform 1 0 43056 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1624047346
transform -1 0 44068 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_460
timestamp 1624047346
transform 1 0 43424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_467
timestamp 1624047346
transform 1 0 44068 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_471
timestamp 1624047346
transform 1 0 44436 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_457
timestamp 1624047346
transform 1 0 43148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_470
timestamp 1624047346
transform 1 0 44344 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _284_
timestamp 1624047346
transform 1 0 44528 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1624047346
transform 1 0 45448 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input92
timestamp 1624047346
transform -1 0 46092 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output245
timestamp 1624047346
transform -1 0 45080 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_481
timestamp 1624047346
transform 1 0 45356 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_478
timestamp 1624047346
transform 1 0 45080 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_485
timestamp 1624047346
transform 1 0 45724 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1624047346
transform 1 0 46920 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624047346
transform 1 0 46460 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1624047346
transform -1 0 47288 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output226
timestamp 1624047346
transform 1 0 46184 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1624047346
transform 1 0 46092 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1624047346
transform 1 0 46552 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_489
timestamp 1624047346
transform 1 0 46092 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_494
timestamp 1624047346
transform 1 0 46552 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_502
timestamp 1624047346
transform 1 0 47288 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _139_
timestamp 1624047346
transform -1 0 47932 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624047346
transform 1 0 48300 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1624047346
transform -1 0 48760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output182
timestamp 1624047346
transform -1 0 49128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_507
timestamp 1624047346
transform 1 0 47748 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_513
timestamp 1624047346
transform 1 0 48300 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_518
timestamp 1624047346
transform 1 0 48760 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_509
timestamp 1624047346
transform 1 0 47932 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_514
timestamp 1624047346
transform 1 0 48392 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _258_
timestamp 1624047346
transform 1 0 50140 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624047346
transform 1 0 49128 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1624047346
transform -1 0 50048 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output241
timestamp 1624047346
transform -1 0 50784 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624047346
transform -1 0 49404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_525
timestamp 1624047346
transform 1 0 49404 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_522
timestamp 1624047346
transform 1 0 49128 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_532
timestamp 1624047346
transform 1 0 50048 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624047346
transform 1 0 51796 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output223
timestamp 1624047346
transform -1 0 51888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_542
timestamp 1624047346
transform 1 0 50968 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_550
timestamp 1624047346
transform 1 0 51704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_552
timestamp 1624047346
transform 1 0 51888 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_540
timestamp 1624047346
transform 1 0 50784 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_552
timestamp 1624047346
transform 1 0 51888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_559
timestamp 1624047346
transform 1 0 52532 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output207
timestamp 1624047346
transform -1 0 52624 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1624047346
transform 1 0 52256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1624047346
transform 1 0 52900 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1624047346
transform 1 0 53636 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_566
timestamp 1624047346
transform 1 0 53176 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1624047346
transform -1 0 53728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624047346
transform 1 0 53544 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_572
timestamp 1624047346
transform 1 0 53728 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_560
timestamp 1624047346
transform 1 0 52624 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _221_
timestamp 1624047346
transform 1 0 54004 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624047346
transform 1 0 54464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output134
timestamp 1624047346
transform -1 0 55292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output228
timestamp 1624047346
transform -1 0 55108 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_581
timestamp 1624047346
transform 1 0 54556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_589
timestamp 1624047346
transform 1 0 55292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1624047346
transform 1 0 54280 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_582
timestamp 1624047346
transform 1 0 54648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_587
timestamp 1624047346
transform 1 0 55108 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1624047346
transform -1 0 56028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1624047346
transform -1 0 56028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624047346
transform -1 0 56764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output183
timestamp 1624047346
transform 1 0 56396 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_597
timestamp 1624047346
transform 1 0 56028 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_605
timestamp 1624047346
transform 1 0 56764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_593
timestamp 1624047346
transform 1 0 55660 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_597
timestamp 1624047346
transform 1 0 56028 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_605
timestamp 1624047346
transform 1 0 56764 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _272_
timestamp 1624047346
transform 1 0 57132 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624047346
transform 1 0 57132 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 58236 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_610
timestamp 1624047346
transform 1 0 57224 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_614
timestamp 1624047346
transform 1 0 57592 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1624047346
transform 1 0 58236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_618
timestamp 1624047346
transform 1 0 57960 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624047346
transform -1 0 58880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624047346
transform -1 0 58880 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1624047346
transform 1 0 58512 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624047346
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output168
timestamp 1624047346
transform -1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output218
timestamp 1624047346
transform -1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_7
timestamp 1624047346
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_15
timestamp 1624047346
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624047346
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output232
timestamp 1624047346
transform -1 0 3220 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1624047346
transform -1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_23
timestamp 1624047346
transform 1 0 3220 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1624047346
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output168_A
timestamp 1624047346
transform -1 0 4600 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_38 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 4600 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_50
timestamp 1624047346
transform 1 0 5704 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1624047346
transform -1 0 6808 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 6440 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_62
timestamp 1624047346
transform 1 0 6808 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_74
timestamp 1624047346
transform 1 0 7912 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624047346
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 1624047346
transform 1 0 9476 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1624047346
transform -1 0 10304 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_87
timestamp 1624047346
transform 1 0 9108 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_94
timestamp 1624047346
transform 1 0 9752 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_100
timestamp 1624047346
transform 1 0 10304 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1624047346
transform -1 0 11132 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output237_A
timestamp 1624047346
transform -1 0 11684 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_106
timestamp 1624047346
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1624047346
transform 1 0 11132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_115
timestamp 1624047346
transform 1 0 11684 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output187_A
timestamp 1624047346
transform -1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_127
timestamp 1624047346
transform 1 0 12788 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_131
timestamp 1624047346
transform 1 0 13156 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_134
timestamp 1624047346
transform 1 0 13432 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _196_
timestamp 1624047346
transform -1 0 15180 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624047346
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__A
timestamp 1624047346
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_142
timestamp 1624047346
transform 1 0 14168 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1624047346
transform 1 0 14536 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1624047346
transform -1 0 16376 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1624047346
transform 1 0 15548 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1624047346
transform 1 0 15180 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_159
timestamp 1624047346
transform 1 0 15732 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_166
timestamp 1624047346
transform 1 0 16376 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1624047346
transform 1 0 17388 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1624047346
transform -1 0 17020 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_173
timestamp 1624047346
transform 1 0 17020 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_180
timestamp 1624047346
transform 1 0 17664 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624047346
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624047346
transform 1 0 18400 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624047346
transform -1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_191
timestamp 1624047346
transform 1 0 18676 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1624047346
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1624047346
transform -1 0 21160 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A0
timestamp 1624047346
transform -1 0 20332 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1624047346
transform 1 0 19780 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_209
timestamp 1624047346
transform 1 0 20332 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_215
timestamp 1624047346
transform 1 0 20884 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_218
timestamp 1624047346
transform 1 0 21160 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 1624047346
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__A1
timestamp 1624047346
transform -1 0 22172 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_226
timestamp 1624047346
transform 1 0 21896 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1624047346
transform 1 0 22172 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1624047346
transform -1 0 23368 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output219_A
timestamp 1624047346
transform -1 0 24380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_236
timestamp 1624047346
transform 1 0 22816 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_242
timestamp 1624047346
transform 1 0 23368 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_250
timestamp 1624047346
transform 1 0 24104 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1624047346
transform -1 0 25944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624047346
transform 1 0 24748 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1624047346
transform -1 0 25300 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_253
timestamp 1624047346
transform 1 0 24380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_258
timestamp 1624047346
transform 1 0 24840 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_263
timestamp 1624047346
transform 1 0 25300 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output242
timestamp 1624047346
transform -1 0 27508 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1624047346
transform -1 0 26772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_270
timestamp 1624047346
transform 1 0 25944 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1624047346
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_279
timestamp 1624047346
transform 1 0 26772 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1624047346
transform -1 0 28152 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output204
timestamp 1624047346
transform -1 0 28888 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1624047346
transform 1 0 27508 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_294
timestamp 1624047346
transform 1 0 28152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_302
timestamp 1624047346
transform 1 0 28888 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 1624047346
transform 1 0 29256 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624047346
transform 1 0 29992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624047346
transform -1 0 30728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_309
timestamp 1624047346
transform 1 0 29532 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_313
timestamp 1624047346
transform 1 0 29900 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_315
timestamp 1624047346
transform 1 0 30084 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624047346
transform -1 0 31280 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output243_A
timestamp 1624047346
transform 1 0 31648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_322
timestamp 1624047346
transform 1 0 30728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1624047346
transform 1 0 31280 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_334
timestamp 1624047346
transform 1 0 31832 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 1624047346
transform 1 0 32200 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1624047346
transform -1 0 33028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_341
timestamp 1624047346
transform 1 0 32476 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_347
timestamp 1624047346
transform 1 0 33028 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1624047346
transform -1 0 34316 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1624047346
transform -1 0 34868 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_355
timestamp 1624047346
transform 1 0 33764 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_361
timestamp 1624047346
transform 1 0 34316 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_367
timestamp 1624047346
transform 1 0 34868 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624047346
transform 1 0 35236 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1624047346
transform 1 0 35696 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output198
timestamp 1624047346
transform -1 0 36708 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_372
timestamp 1624047346
transform 1 0 35328 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_379
timestamp 1624047346
transform 1 0 35972 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_387
timestamp 1624047346
transform 1 0 36708 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1624047346
transform -1 0 37352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1624047346
transform -1 0 38272 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_394
timestamp 1624047346
transform 1 0 37352 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_400
timestamp 1624047346
transform 1 0 37904 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_404
timestamp 1624047346
transform 1 0 38272 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1624047346
transform 1 0 38640 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output186
timestamp 1624047346
transform -1 0 39928 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_411
timestamp 1624047346
transform 1 0 38916 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_417
timestamp 1624047346
transform 1 0 39468 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1624047346
transform -1 0 41216 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624047346
transform 1 0 40480 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_422
timestamp 1624047346
transform 1 0 39928 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_429
timestamp 1624047346
transform 1 0 40572 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_436
timestamp 1624047346
transform 1 0 41216 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output185
timestamp 1624047346
transform -1 0 42228 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624047346
transform -1 0 42780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_442
timestamp 1624047346
transform 1 0 41768 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_447
timestamp 1624047346
transform 1 0 42228 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1624047346
transform 1 0 42780 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1624047346
transform -1 0 44068 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1624047346
transform 1 0 44436 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1624047346
transform 1 0 43148 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_460
timestamp 1624047346
transform 1 0 43424 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_467
timestamp 1624047346
transform 1 0 44068 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624047346
transform 1 0 45724 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624047346
transform -1 0 45264 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1624047346
transform -1 0 46000 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_474
timestamp 1624047346
transform 1 0 44712 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1624047346
transform 1 0 45264 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_484
timestamp 1624047346
transform 1 0 45632 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_488
timestamp 1624047346
transform 1 0 46000 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624047346
transform -1 0 47472 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1624047346
transform -1 0 46552 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_494
timestamp 1624047346
transform 1 0 46552 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_504
timestamp 1624047346
transform 1 0 47472 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1624047346
transform -1 0 48208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1624047346
transform -1 0 48760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_512
timestamp 1624047346
transform 1 0 48208 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_518
timestamp 1624047346
transform 1 0 48760 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1624047346
transform -1 0 50232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__S
timestamp 1624047346
transform 1 0 49496 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_528
timestamp 1624047346
transform 1 0 49680 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_534
timestamp 1624047346
transform 1 0 50232 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624047346
transform 1 0 50968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output207_A
timestamp 1624047346
transform -1 0 52164 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_543
timestamp 1624047346
transform 1 0 51060 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_551
timestamp 1624047346
transform 1 0 51796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_555
timestamp 1624047346
transform 1 0 52164 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624047346
transform -1 0 53912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624047346
transform -1 0 53360 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624047346
transform -1 0 52716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_561
timestamp 1624047346
transform 1 0 52716 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_565
timestamp 1624047346
transform 1 0 53084 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_568
timestamp 1624047346
transform 1 0 53360 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1624047346
transform -1 0 55292 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A
timestamp 1624047346
transform -1 0 54464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_574
timestamp 1624047346
transform 1 0 53912 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_580
timestamp 1624047346
transform 1 0 54464 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_586
timestamp 1624047346
transform 1 0 55016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_589
timestamp 1624047346
transform 1 0 55292 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624047346
transform 1 0 56212 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624047346
transform -1 0 56488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624047346
transform -1 0 55844 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_595
timestamp 1624047346
transform 1 0 55844 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_602
timestamp 1624047346
transform 1 0 56488 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output173
timestamp 1624047346
transform 1 0 57868 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output174
timestamp 1624047346
transform 1 0 57132 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_608
timestamp 1624047346
transform 1 0 57040 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 1624047346
transform 1 0 57500 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1624047346
transform 1 0 58236 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624047346
transform -1 0 58880 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624047346
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output178
timestamp 1624047346
transform -1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output220
timestamp 1624047346
transform -1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1624047346
transform 1 0 1748 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15
timestamp 1624047346
transform 1 0 2484 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output133_A
timestamp 1624047346
transform -1 0 3312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output232_A
timestamp 1624047346
transform 1 0 3680 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_21
timestamp 1624047346
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_24
timestamp 1624047346
transform 1 0 3312 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1624047346
transform 1 0 3864 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_42
timestamp 1624047346
transform 1 0 4968 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624047346
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_54
timestamp 1624047346
transform 1 0 6072 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_58
timestamp 1624047346
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_70
timestamp 1624047346
transform 1 0 7544 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_82
timestamp 1624047346
transform 1 0 8648 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output180_A
timestamp 1624047346
transform 1 0 10212 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp 1624047346
transform 1 0 9752 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_98
timestamp 1624047346
transform 1 0 10120 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_101
timestamp 1624047346
transform 1 0 10396 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624047346
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1624047346
transform 1 0 11500 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_115
timestamp 1624047346
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_127
timestamp 1624047346
transform 1 0 12788 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_139
timestamp 1624047346
transform 1 0 13892 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1624047346
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1624047346
transform 1 0 15180 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624047346
transform -1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_156
timestamp 1624047346
transform 1 0 15456 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_162
timestamp 1624047346
transform 1 0 16008 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624047346
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1624047346
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1624047346
transform -1 0 18308 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A
timestamp 1624047346
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_170
timestamp 1624047346
transform 1 0 16744 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_174
timestamp 1624047346
transform 1 0 17112 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1624047346
transform 1 0 17756 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624047346
transform -1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1624047346
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_187
timestamp 1624047346
transform 1 0 18308 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_193
timestamp 1624047346
transform 1 0 18860 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_199
timestamp 1624047346
transform 1 0 19412 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__262__S
timestamp 1624047346
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_211
timestamp 1624047346
transform 1 0 20516 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624047346
transform 1 0 22080 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output149_A
timestamp 1624047346
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_219
timestamp 1624047346
transform 1 0 21252 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_227
timestamp 1624047346
transform 1 0 21988 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_229
timestamp 1624047346
transform 1 0 22172 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1624047346
transform 1 0 22908 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_249
timestamp 1624047346
transform 1 0 24012 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _104_
timestamp 1624047346
transform 1 0 25024 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _213_
timestamp 1624047346
transform -1 0 25944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1624047346
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_253
timestamp 1624047346
transform 1 0 24380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_256
timestamp 1624047346
transform 1 0 24656 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_263
timestamp 1624047346
transform 1 0 25300 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624047346
transform 1 0 27324 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A
timestamp 1624047346
transform -1 0 26496 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_270
timestamp 1624047346
transform 1 0 25944 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_276
timestamp 1624047346
transform 1 0 26496 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_284
timestamp 1624047346
transform 1 0 27232 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_286
timestamp 1624047346
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1624047346
transform -1 0 28336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1624047346
transform 1 0 28888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__S
timestamp 1624047346
transform 1 0 27600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_290
timestamp 1624047346
transform 1 0 27784 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_296
timestamp 1624047346
transform 1 0 28336 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__193__A
timestamp 1624047346
transform -1 0 29624 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_304
timestamp 1624047346
transform 1 0 29072 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_310
timestamp 1624047346
transform 1 0 29624 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_322
timestamp 1624047346
transform 1 0 30728 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_334
timestamp 1624047346
transform 1 0 31832 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624047346
transform 1 0 32568 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_343
timestamp 1624047346
transform 1 0 32660 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_355
timestamp 1624047346
transform 1 0 33764 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_367
timestamp 1624047346
transform 1 0 34868 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624047346
transform -1 0 35696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A
timestamp 1624047346
transform 1 0 36064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_373
timestamp 1624047346
transform 1 0 35420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_376
timestamp 1624047346
transform 1 0 35696 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_382
timestamp 1624047346
transform 1 0 36248 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624047346
transform 1 0 37812 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 1624047346
transform 1 0 36800 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1624047346
transform -1 0 38456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_391
timestamp 1624047346
transform 1 0 37076 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_400
timestamp 1624047346
transform 1 0 37904 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624047346
transform -1 0 39100 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1624047346
transform 1 0 39468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_406
timestamp 1624047346
transform 1 0 38456 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_410
timestamp 1624047346
transform 1 0 38824 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_413
timestamp 1624047346
transform 1 0 39100 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_419
timestamp 1624047346
transform 1 0 39652 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp 1624047346
transform -1 0 41216 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _148_
timestamp 1624047346
transform -1 0 40296 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_426
timestamp 1624047346
transform 1 0 40296 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_432
timestamp 1624047346
transform 1 0 40848 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_436
timestamp 1624047346
transform 1 0 41216 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1624047346
transform -1 0 41860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 1624047346
transform -1 0 42504 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_443
timestamp 1624047346
transform 1 0 41860 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_450
timestamp 1624047346
transform 1 0 42504 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624047346
transform 1 0 43056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624047346
transform -1 0 43608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A0
timestamp 1624047346
transform 1 0 43976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_457
timestamp 1624047346
transform 1 0 43148 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_462
timestamp 1624047346
transform 1 0 43608 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_468
timestamp 1624047346
transform 1 0 44160 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A0
timestamp 1624047346
transform -1 0 44712 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__A1
timestamp 1624047346
transform 1 0 45080 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A1
timestamp 1624047346
transform 1 0 45632 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_474
timestamp 1624047346
transform 1 0 44712 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_480
timestamp 1624047346
transform 1 0 45264 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_486
timestamp 1624047346
transform 1 0 45816 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A
timestamp 1624047346
transform 1 0 47472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__A0
timestamp 1624047346
transform -1 0 46920 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__S
timestamp 1624047346
transform 1 0 46184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_492
timestamp 1624047346
transform 1 0 46368 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_498
timestamp 1624047346
transform 1 0 46920 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624047346
transform 1 0 48300 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_506
timestamp 1624047346
transform 1 0 47656 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_512
timestamp 1624047346
transform 1 0 48208 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_514
timestamp 1624047346
transform 1 0 48392 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_526
timestamp 1624047346
transform 1 0 49496 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_538
timestamp 1624047346
transform 1 0 50600 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_550
timestamp 1624047346
transform 1 0 51704 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624047346
transform 1 0 53544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_562
timestamp 1624047346
transform 1 0 52808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_571
timestamp 1624047346
transform 1 0 53636 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1624047346
transform 1 0 55108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_583
timestamp 1624047346
transform 1 0 54740 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_589
timestamp 1624047346
transform 1 0 55292 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624047346
transform -1 0 56948 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624047346
transform -1 0 56396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1624047346
transform -1 0 55844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_595
timestamp 1624047346
transform 1 0 55844 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_601
timestamp 1624047346
transform 1 0 56396 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1624047346
transform -1 0 58236 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1624047346
transform -1 0 57592 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_607
timestamp 1624047346
transform 1 0 56948 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_614
timestamp 1624047346
transform 1 0 57592 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1624047346
transform 1 0 58236 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624047346
transform -1 0 58880 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624047346
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1624047346
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output165_A
timestamp 1624047346
transform 1 0 2392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_7
timestamp 1624047346
transform 1 0 1748 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_13
timestamp 1624047346
transform 1 0 2300 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_16
timestamp 1624047346
transform 1 0 2576 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624047346
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_28
timestamp 1624047346
transform 1 0 3680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624047346
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624047346
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_54
timestamp 1624047346
transform 1 0 6072 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_66
timestamp 1624047346
transform 1 0 7176 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_78
timestamp 1624047346
transform 1 0 8280 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624047346
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_87
timestamp 1624047346
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_99
timestamp 1624047346
transform 1 0 10212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1624047346
transform 1 0 11316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1624047346
transform 1 0 12420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624047346
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_135
timestamp 1624047346
transform 1 0 13524 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_144
timestamp 1624047346
transform 1 0 14352 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__A1
timestamp 1624047346
transform -1 0 15916 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1624047346
transform -1 0 16560 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_156
timestamp 1624047346
transform 1 0 15456 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1624047346
transform 1 0 15916 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_165
timestamp 1624047346
transform 1 0 16284 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_168
timestamp 1624047346
transform 1 0 16560 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__S
timestamp 1624047346
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_176
timestamp 1624047346
transform 1 0 17296 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_179
timestamp 1624047346
transform 1 0 17572 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624047346
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_191
timestamp 1624047346
transform 1 0 18676 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_199
timestamp 1624047346
transform 1 0 19412 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_201
timestamp 1624047346
transform 1 0 19596 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_213
timestamp 1624047346
transform 1 0 20700 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_225
timestamp 1624047346
transform 1 0 21804 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_237
timestamp 1624047346
transform 1 0 22908 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_249
timestamp 1624047346
transform 1 0 24012 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624047346
transform 1 0 24748 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1624047346
transform 1 0 24840 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output150_A
timestamp 1624047346
transform 1 0 27324 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output194_A
timestamp 1624047346
transform 1 0 26404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_270
timestamp 1624047346
transform 1 0 25944 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1624047346
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_277
timestamp 1624047346
transform 1 0 26588 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A1
timestamp 1624047346
transform 1 0 28612 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_287
timestamp 1624047346
transform 1 0 27508 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_301
timestamp 1624047346
transform 1 0 28796 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624047346
transform 1 0 29992 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output204_A
timestamp 1624047346
transform 1 0 29164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_307
timestamp 1624047346
transform 1 0 29348 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_313
timestamp 1624047346
transform 1 0 29900 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_315
timestamp 1624047346
transform 1 0 30084 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_327
timestamp 1624047346
transform 1 0 31188 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_339
timestamp 1624047346
transform 1 0 32292 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_351
timestamp 1624047346
transform 1 0 33396 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_363
timestamp 1624047346
transform 1 0 34500 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624047346
transform 1 0 35236 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_372
timestamp 1624047346
transform 1 0 35328 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_384
timestamp 1624047346
transform 1 0 36432 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1624047346
transform -1 0 37260 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1624047346
transform 1 0 37628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_390
timestamp 1624047346
transform 1 0 36984 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_393
timestamp 1624047346
transform 1 0 37260 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_399
timestamp 1624047346
transform 1 0 37812 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A0
timestamp 1624047346
transform -1 0 39928 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output144_A
timestamp 1624047346
transform 1 0 38732 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_407
timestamp 1624047346
transform 1 0 38548 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_411
timestamp 1624047346
transform 1 0 38916 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1624047346
transform 1 0 39652 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624047346
transform 1 0 40480 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1624047346
transform -1 0 41216 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_422
timestamp 1624047346
transform 1 0 39928 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_429
timestamp 1624047346
transform 1 0 40572 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_436
timestamp 1624047346
transform 1 0 41216 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1624047346
transform -1 0 42228 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A1
timestamp 1624047346
transform -1 0 42780 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_444
timestamp 1624047346
transform 1 0 41952 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_447
timestamp 1624047346
transform 1 0 42228 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_453
timestamp 1624047346
transform 1 0 42780 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__S
timestamp 1624047346
transform 1 0 43148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__S
timestamp 1624047346
transform 1 0 43700 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__S
timestamp 1624047346
transform 1 0 44252 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_459
timestamp 1624047346
transform 1 0 43332 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_465
timestamp 1624047346
transform 1 0 43884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_471
timestamp 1624047346
transform 1 0 44436 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624047346
transform 1 0 45724 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_483
timestamp 1624047346
transform 1 0 45540 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_486
timestamp 1624047346
transform 1 0 45816 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_498
timestamp 1624047346
transform 1 0 46920 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_510
timestamp 1624047346
transform 1 0 48024 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_522
timestamp 1624047346
transform 1 0 49128 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_534
timestamp 1624047346
transform 1 0 50232 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624047346
transform 1 0 50968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_543
timestamp 1624047346
transform 1 0 51060 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_555
timestamp 1624047346
transform 1 0 52164 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_567
timestamp 1624047346
transform 1 0 53268 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_579
timestamp 1624047346
transform 1 0 54372 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624047346
transform 1 0 56212 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1624047346
transform -1 0 56856 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_591
timestamp 1624047346
transform 1 0 55476 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_600
timestamp 1624047346
transform 1 0 56304 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_606
timestamp 1624047346
transform 1 0 56856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1624047346
transform -1 0 58236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 1624047346
transform -1 0 57500 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_613
timestamp 1624047346
transform 1 0 57500 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_621
timestamp 1624047346
transform 1 0 58236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624047346
transform -1 0 58880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624047346
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1624047346
transform -1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output178_A
timestamp 1624047346
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_5
timestamp 1624047346
transform 1 0 1564 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_11
timestamp 1624047346
transform 1 0 2116 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_23
timestamp 1624047346
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_35
timestamp 1624047346
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1624047346
transform 1 0 5428 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624047346
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1624047346
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_58
timestamp 1624047346
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1624047346
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1624047346
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1624047346
transform 1 0 9752 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624047346
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_106
timestamp 1624047346
transform 1 0 10856 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_115
timestamp 1624047346
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_127
timestamp 1624047346
transform 1 0 12788 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_139
timestamp 1624047346
transform 1 0 13892 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_151
timestamp 1624047346
transform 1 0 14996 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_163
timestamp 1624047346
transform 1 0 16100 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624047346
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output201_A
timestamp 1624047346
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_174
timestamp 1624047346
transform 1 0 17112 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_186
timestamp 1624047346
transform 1 0 18216 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_198
timestamp 1624047346
transform 1 0 19320 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_210
timestamp 1624047346
transform 1 0 20424 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624047346
transform 1 0 22080 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_222
timestamp 1624047346
transform 1 0 21528 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_229
timestamp 1624047346
transform 1 0 22172 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_241
timestamp 1624047346
transform 1 0 23276 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1624047346
transform 1 0 25300 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_253
timestamp 1624047346
transform 1 0 24380 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_261
timestamp 1624047346
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_266
timestamp 1624047346
transform 1 0 25576 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624047346
transform 1 0 27324 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_278
timestamp 1624047346
transform 1 0 26680 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_284
timestamp 1624047346
transform 1 0 27232 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_286
timestamp 1624047346
transform 1 0 27416 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_298
timestamp 1624047346
transform 1 0 28520 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_310
timestamp 1624047346
transform 1 0 29624 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_322
timestamp 1624047346
transform 1 0 30728 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_334
timestamp 1624047346
transform 1 0 31832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624047346
transform 1 0 32568 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_343
timestamp 1624047346
transform 1 0 32660 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_2  _253_
timestamp 1624047346
transform -1 0 35328 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1624047346
transform 1 0 33948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_355
timestamp 1624047346
transform 1 0 33764 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_359
timestamp 1624047346
transform 1 0 34132 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__S
timestamp 1624047346
transform 1 0 35696 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_372
timestamp 1624047346
transform 1 0 35328 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_378
timestamp 1624047346
transform 1 0 35880 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624047346
transform 1 0 37812 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_390
timestamp 1624047346
transform 1 0 36984 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_398
timestamp 1624047346
transform 1 0 37720 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_400
timestamp 1624047346
transform 1 0 37904 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__S
timestamp 1624047346
transform 1 0 39560 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_412
timestamp 1624047346
transform 1 0 39008 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_420
timestamp 1624047346
transform 1 0 39744 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1624047346
transform -1 0 40940 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A0
timestamp 1624047346
transform -1 0 41492 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__S
timestamp 1624047346
transform 1 0 40204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_424
timestamp 1624047346
transform 1 0 40112 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_427
timestamp 1624047346
transform 1 0 40388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_433
timestamp 1624047346
transform 1 0 40940 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_439
timestamp 1624047346
transform 1 0 41492 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_451
timestamp 1624047346
transform 1 0 42596 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624047346
transform 1 0 43056 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_455
timestamp 1624047346
transform 1 0 42964 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_457
timestamp 1624047346
transform 1 0 43148 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_469
timestamp 1624047346
transform 1 0 44252 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_481
timestamp 1624047346
transform 1 0 45356 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_493
timestamp 1624047346
transform 1 0 46460 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_505
timestamp 1624047346
transform 1 0 47564 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624047346
transform 1 0 48300 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_514
timestamp 1624047346
transform 1 0 48392 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_526
timestamp 1624047346
transform 1 0 49496 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_538
timestamp 1624047346
transform 1 0 50600 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_550
timestamp 1624047346
transform 1 0 51704 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624047346
transform 1 0 53544 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_562
timestamp 1624047346
transform 1 0 52808 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_571
timestamp 1624047346
transform 1 0 53636 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_583
timestamp 1624047346
transform 1 0 54740 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1624047346
transform -1 0 57040 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__272__S
timestamp 1624047346
transform 1 0 56304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_595
timestamp 1624047346
transform 1 0 55844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_599
timestamp 1624047346
transform 1 0 56212 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_602
timestamp 1624047346
transform 1 0 56488 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1624047346
transform -1 0 58236 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624047346
transform -1 0 57592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_608
timestamp 1624047346
transform 1 0 57040 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_614
timestamp 1624047346
transform 1 0 57592 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1624047346
transform 1 0 58236 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624047346
transform -1 0 58880 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624047346
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624047346
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output238
timestamp 1624047346
transform -1 0 1748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1624047346
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1624047346
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_7
timestamp 1624047346
transform 1 0 1748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624047346
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1624047346
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624047346
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_19
timestamp 1624047346
transform 1 0 2852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_31
timestamp 1624047346
transform 1 0 3956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_42
timestamp 1624047346
transform 1 0 4968 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1624047346
transform 1 0 5060 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624047346
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_54
timestamp 1624047346
transform 1 0 6072 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_66
timestamp 1624047346
transform 1 0 7176 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1624047346
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_58
timestamp 1624047346
transform 1 0 6440 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_78
timestamp 1624047346
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_70
timestamp 1624047346
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_82
timestamp 1624047346
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624047346
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_87
timestamp 1624047346
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_99
timestamp 1624047346
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_94
timestamp 1624047346
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624047346
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_111
timestamp 1624047346
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_106
timestamp 1624047346
transform 1 0 10856 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_115
timestamp 1624047346
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_123
timestamp 1624047346
transform 1 0 12420 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1624047346
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624047346
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1624047346
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_144
timestamp 1624047346
transform 1 0 14352 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_139
timestamp 1624047346
transform 1 0 13892 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_151
timestamp 1624047346
transform 1 0 14996 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_156
timestamp 1624047346
transform 1 0 15456 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1624047346
transform 1 0 16560 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_163
timestamp 1624047346
transform 1 0 16100 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624047346
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1624047346
transform 1 0 17664 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_172
timestamp 1624047346
transform 1 0 16928 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1624047346
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624047346
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_192
timestamp 1624047346
transform 1 0 18768 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_201
timestamp 1624047346
transform 1 0 19596 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1624047346
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_213
timestamp 1624047346
transform 1 0 20700 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1624047346
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624047346
transform 1 0 22080 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_225
timestamp 1624047346
transform 1 0 21804 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_220
timestamp 1624047346
transform 1 0 21344 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_229
timestamp 1624047346
transform 1 0 22172 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_237
timestamp 1624047346
transform 1 0 22908 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_249
timestamp 1624047346
transform 1 0 24012 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_241
timestamp 1624047346
transform 1 0 23276 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624047346
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1624047346
transform 1 0 24840 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_253
timestamp 1624047346
transform 1 0 24380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_265
timestamp 1624047346
transform 1 0 25484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624047346
transform 1 0 27324 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_270
timestamp 1624047346
transform 1 0 25944 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_282
timestamp 1624047346
transform 1 0 27048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_277
timestamp 1624047346
transform 1 0 26588 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_286
timestamp 1624047346
transform 1 0 27416 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_294
timestamp 1624047346
transform 1 0 28152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_298
timestamp 1624047346
transform 1 0 28520 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624047346
transform 1 0 29992 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_306
timestamp 1624047346
transform 1 0 29256 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_315
timestamp 1624047346
transform 1 0 30084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_310
timestamp 1624047346
transform 1 0 29624 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_327
timestamp 1624047346
transform 1 0 31188 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_322
timestamp 1624047346
transform 1 0 30728 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_334
timestamp 1624047346
transform 1 0 31832 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624047346
transform 1 0 32568 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_339
timestamp 1624047346
transform 1 0 32292 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_351
timestamp 1624047346
transform 1 0 33396 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_343
timestamp 1624047346
transform 1 0 32660 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_363
timestamp 1624047346
transform 1 0 34500 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_355
timestamp 1624047346
transform 1 0 33764 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_367
timestamp 1624047346
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624047346
transform 1 0 35236 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_372
timestamp 1624047346
transform 1 0 35328 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_384
timestamp 1624047346
transform 1 0 36432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_379
timestamp 1624047346
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624047346
transform 1 0 37812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_396
timestamp 1624047346
transform 1 0 37536 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_391
timestamp 1624047346
transform 1 0 37076 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_400
timestamp 1624047346
transform 1 0 37904 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_408
timestamp 1624047346
transform 1 0 38640 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_420
timestamp 1624047346
transform 1 0 39744 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_412
timestamp 1624047346
transform 1 0 39008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624047346
transform 1 0 40480 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A1
timestamp 1624047346
transform 1 0 40756 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_429
timestamp 1624047346
transform 1 0 40572 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1624047346
transform 1 0 40940 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_424
timestamp 1624047346
transform 1 0 40112 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_436
timestamp 1624047346
transform 1 0 41216 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1624047346
transform 1 0 42044 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_448
timestamp 1624047346
transform 1 0 42320 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624047346
transform 1 0 43056 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1624047346
transform 1 0 43148 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_469
timestamp 1624047346
transform 1 0 44252 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_457
timestamp 1624047346
transform 1 0 43148 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_469
timestamp 1624047346
transform 1 0 44252 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624047346
transform 1 0 45724 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_481
timestamp 1624047346
transform 1 0 45356 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_486
timestamp 1624047346
transform 1 0 45816 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_481
timestamp 1624047346
transform 1 0 45356 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_498
timestamp 1624047346
transform 1 0 46920 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_493
timestamp 1624047346
transform 1 0 46460 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1624047346
transform 1 0 47564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624047346
transform 1 0 48300 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_510
timestamp 1624047346
transform 1 0 48024 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_514
timestamp 1624047346
transform 1 0 48392 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_522
timestamp 1624047346
transform 1 0 49128 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_534
timestamp 1624047346
transform 1 0 50232 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_526
timestamp 1624047346
transform 1 0 49496 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_538
timestamp 1624047346
transform 1 0 50600 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624047346
transform 1 0 50968 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_543
timestamp 1624047346
transform 1 0 51060 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_555
timestamp 1624047346
transform 1 0 52164 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_550
timestamp 1624047346
transform 1 0 51704 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624047346
transform 1 0 53544 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_567
timestamp 1624047346
transform 1 0 53268 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_562
timestamp 1624047346
transform 1 0 52808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_571
timestamp 1624047346
transform 1 0 53636 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_579
timestamp 1624047346
transform 1 0 54372 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_583
timestamp 1624047346
transform 1 0 54740 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624047346
transform 1 0 56212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_591
timestamp 1624047346
transform 1 0 55476 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_600
timestamp 1624047346
transform 1 0 56304 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_606
timestamp 1624047346
transform 1 0 56856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_595
timestamp 1624047346
transform 1 0 55844 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output224
timestamp 1624047346
transform 1 0 57868 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1624047346
transform -1 0 57132 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output224_A
timestamp 1624047346
transform -1 0 57868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_609
timestamp 1624047346
transform 1 0 57132 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1624047346
transform 1 0 58236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_607
timestamp 1624047346
transform 1 0 56948 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1624047346
transform 1 0 57868 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624047346
transform -1 0 58880 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624047346
transform -1 0 58880 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _268_
timestamp 1624047346
transform 1 0 1932 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624047346
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__S
timestamp 1624047346
transform -1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_5
timestamp 1624047346
transform 1 0 1564 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624047346
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__268__A0
timestamp 1624047346
transform -1 0 3312 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1624047346
transform 1 0 2760 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1624047346
transform 1 0 3312 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_28
timestamp 1624047346
transform 1 0 3680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1624047346
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1624047346
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_54
timestamp 1624047346
transform 1 0 6072 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_66
timestamp 1624047346
transform 1 0 7176 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_78
timestamp 1624047346
transform 1 0 8280 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624047346
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_87
timestamp 1624047346
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_99
timestamp 1624047346
transform 1 0 10212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_111
timestamp 1624047346
transform 1 0 11316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_123
timestamp 1624047346
transform 1 0 12420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624047346
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_135
timestamp 1624047346
transform 1 0 13524 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_144
timestamp 1624047346
transform 1 0 14352 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_156
timestamp 1624047346
transform 1 0 15456 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1624047346
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1624047346
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624047346
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_192
timestamp 1624047346
transform 1 0 18768 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_201
timestamp 1624047346
transform 1 0 19596 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_213
timestamp 1624047346
transform 1 0 20700 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_225
timestamp 1624047346
transform 1 0 21804 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_237
timestamp 1624047346
transform 1 0 22908 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_249
timestamp 1624047346
transform 1 0 24012 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624047346
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_258
timestamp 1624047346
transform 1 0 24840 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_270
timestamp 1624047346
transform 1 0 25944 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_282
timestamp 1624047346
transform 1 0 27048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_294
timestamp 1624047346
transform 1 0 28152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624047346
transform 1 0 29992 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_306
timestamp 1624047346
transform 1 0 29256 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_315
timestamp 1624047346
transform 1 0 30084 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_327
timestamp 1624047346
transform 1 0 31188 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_339
timestamp 1624047346
transform 1 0 32292 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_351
timestamp 1624047346
transform 1 0 33396 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_363
timestamp 1624047346
transform 1 0 34500 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1624047346
transform 1 0 35236 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_372
timestamp 1624047346
transform 1 0 35328 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_384
timestamp 1624047346
transform 1 0 36432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_396
timestamp 1624047346
transform 1 0 37536 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_408
timestamp 1624047346
transform 1 0 38640 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_420
timestamp 1624047346
transform 1 0 39744 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1624047346
transform 1 0 40480 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_429
timestamp 1624047346
transform 1 0 40572 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_441
timestamp 1624047346
transform 1 0 41676 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_453
timestamp 1624047346
transform 1 0 42780 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_465
timestamp 1624047346
transform 1 0 43884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1624047346
transform 1 0 45724 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_477
timestamp 1624047346
transform 1 0 44988 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_486
timestamp 1624047346
transform 1 0 45816 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_498
timestamp 1624047346
transform 1 0 46920 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_510
timestamp 1624047346
transform 1 0 48024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_522
timestamp 1624047346
transform 1 0 49128 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_534
timestamp 1624047346
transform 1 0 50232 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1624047346
transform 1 0 50968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_543
timestamp 1624047346
transform 1 0 51060 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_555
timestamp 1624047346
transform 1 0 52164 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_567
timestamp 1624047346
transform 1 0 53268 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1624047346
transform -1 0 54188 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_573
timestamp 1624047346
transform 1 0 53820 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_577
timestamp 1624047346
transform 1 0 54188 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_589
timestamp 1624047346
transform 1 0 55292 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1624047346
transform 1 0 56212 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_597
timestamp 1624047346
transform 1 0 56028 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_600
timestamp 1624047346
transform 1 0 56304 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1624047346
transform -1 0 58236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1624047346
transform -1 0 57500 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_608
timestamp 1624047346
transform 1 0 57040 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_613
timestamp 1624047346
transform 1 0 57500 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_621
timestamp 1624047346
transform 1 0 58236 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624047346
transform -1 0 58880 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624047346
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1624047346
transform -1 0 1656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624047346
transform -1 0 2208 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1624047346
transform 1 0 1656 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_12
timestamp 1624047346
transform 1 0 2208 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_24
timestamp 1624047346
transform 1 0 3312 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_36
timestamp 1624047346
transform 1 0 4416 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1624047346
transform 1 0 5520 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1624047346
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_56
timestamp 1624047346
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_58
timestamp 1624047346
transform 1 0 6440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_70
timestamp 1624047346
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_82
timestamp 1624047346
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_94
timestamp 1624047346
transform 1 0 9752 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1624047346
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_106
timestamp 1624047346
transform 1 0 10856 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1624047346
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_127
timestamp 1624047346
transform 1 0 12788 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_139
timestamp 1624047346
transform 1 0 13892 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_151
timestamp 1624047346
transform 1 0 14996 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_163
timestamp 1624047346
transform 1 0 16100 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1624047346
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_172
timestamp 1624047346
transform 1 0 16928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1624047346
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1624047346
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1624047346
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1624047346
transform 1 0 22080 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_220
timestamp 1624047346
transform 1 0 21344 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_229
timestamp 1624047346
transform 1 0 22172 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_241
timestamp 1624047346
transform 1 0 23276 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_253
timestamp 1624047346
transform 1 0 24380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_265
timestamp 1624047346
transform 1 0 25484 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1624047346
transform 1 0 27324 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1624047346
transform -1 0 26312 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_271
timestamp 1624047346
transform 1 0 26036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_274
timestamp 1624047346
transform 1 0 26312 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_282
timestamp 1624047346
transform 1 0 27048 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_286
timestamp 1624047346
transform 1 0 27416 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _127_
timestamp 1624047346
transform -1 0 28244 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1624047346
transform -1 0 28796 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1624047346
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_301
timestamp 1624047346
transform 1 0 28796 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_313
timestamp 1624047346
transform 1 0 29900 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_325
timestamp 1624047346
transform 1 0 31004 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1624047346
transform 1 0 32568 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_337
timestamp 1624047346
transform 1 0 32108 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_341
timestamp 1624047346
transform 1 0 32476 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_343
timestamp 1624047346
transform 1 0 32660 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_355
timestamp 1624047346
transform 1 0 33764 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1624047346
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1624047346
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1624047346
transform 1 0 37812 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_391
timestamp 1624047346
transform 1 0 37076 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_400
timestamp 1624047346
transform 1 0 37904 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_412
timestamp 1624047346
transform 1 0 39008 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_424
timestamp 1624047346
transform 1 0 40112 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_436
timestamp 1624047346
transform 1 0 41216 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_448
timestamp 1624047346
transform 1 0 42320 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1624047346
transform 1 0 43056 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_457
timestamp 1624047346
transform 1 0 43148 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_469
timestamp 1624047346
transform 1 0 44252 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_481
timestamp 1624047346
transform 1 0 45356 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_493
timestamp 1624047346
transform 1 0 46460 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_505
timestamp 1624047346
transform 1 0 47564 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1624047346
transform 1 0 48300 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_514
timestamp 1624047346
transform 1 0 48392 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_526
timestamp 1624047346
transform 1 0 49496 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_538
timestamp 1624047346
transform 1 0 50600 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_550
timestamp 1624047346
transform 1 0 51704 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1624047346
transform 1 0 53544 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_562
timestamp 1624047346
transform 1 0 52808 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_571
timestamp 1624047346
transform 1 0 53636 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_583
timestamp 1624047346
transform 1 0 54740 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_595
timestamp 1624047346
transform 1 0 55844 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 1624047346
transform -1 0 58236 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1624047346
transform -1 0 57592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_607
timestamp 1624047346
transform 1 0 56948 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_611
timestamp 1624047346
transform 1 0 57316 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_614
timestamp 1624047346
transform 1 0 57592 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_621
timestamp 1624047346
transform 1 0 58236 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624047346
transform -1 0 58880 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624047346
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624047346
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624047346
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1624047346
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624047346
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1624047346
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1624047346
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1624047346
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1624047346
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1624047346
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1624047346
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_87
timestamp 1624047346
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_99
timestamp 1624047346
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1624047346
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1624047346
transform 1 0 12420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1624047346
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_135
timestamp 1624047346
transform 1 0 13524 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_144
timestamp 1624047346
transform 1 0 14352 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_156
timestamp 1624047346
transform 1 0 15456 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_168
timestamp 1624047346
transform 1 0 16560 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_180
timestamp 1624047346
transform 1 0 17664 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1624047346
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_192
timestamp 1624047346
transform 1 0 18768 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_201
timestamp 1624047346
transform 1 0 19596 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_213
timestamp 1624047346
transform 1 0 20700 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_225
timestamp 1624047346
transform 1 0 21804 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_237
timestamp 1624047346
transform 1 0 22908 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_249
timestamp 1624047346
transform 1 0 24012 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _216_
timestamp 1624047346
transform -1 0 26128 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1624047346
transform 1 0 24748 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_258
timestamp 1624047346
transform 1 0 24840 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_266
timestamp 1624047346
transform 1 0 25576 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _215_
timestamp 1624047346
transform -1 0 27140 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_10_272
timestamp 1624047346
transform 1 0 26128 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_283
timestamp 1624047346
transform 1 0 27140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_295
timestamp 1624047346
transform 1 0 28244 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1624047346
transform 1 0 29992 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_307
timestamp 1624047346
transform 1 0 29348 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_313
timestamp 1624047346
transform 1 0 29900 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_315
timestamp 1624047346
transform 1 0 30084 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_327
timestamp 1624047346
transform 1 0 31188 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_339
timestamp 1624047346
transform 1 0 32292 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_351
timestamp 1624047346
transform 1 0 33396 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_363
timestamp 1624047346
transform 1 0 34500 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1624047346
transform 1 0 35236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_372
timestamp 1624047346
transform 1 0 35328 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_384
timestamp 1624047346
transform 1 0 36432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_396
timestamp 1624047346
transform 1 0 37536 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_408
timestamp 1624047346
transform 1 0 38640 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_420
timestamp 1624047346
transform 1 0 39744 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1624047346
transform 1 0 40480 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_429
timestamp 1624047346
transform 1 0 40572 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_441
timestamp 1624047346
transform 1 0 41676 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_453
timestamp 1624047346
transform 1 0 42780 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_465
timestamp 1624047346
transform 1 0 43884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1624047346
transform 1 0 45724 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_477
timestamp 1624047346
transform 1 0 44988 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_486
timestamp 1624047346
transform 1 0 45816 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_498
timestamp 1624047346
transform 1 0 46920 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_510
timestamp 1624047346
transform 1 0 48024 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_522
timestamp 1624047346
transform 1 0 49128 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_534
timestamp 1624047346
transform 1 0 50232 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1624047346
transform 1 0 50968 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_543
timestamp 1624047346
transform 1 0 51060 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_555
timestamp 1624047346
transform 1 0 52164 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_567
timestamp 1624047346
transform 1 0 53268 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_579
timestamp 1624047346
transform 1 0 54372 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1624047346
transform 1 0 56212 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_591
timestamp 1624047346
transform 1 0 55476 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_600
timestamp 1624047346
transform 1 0 56304 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_612
timestamp 1624047346
transform 1 0 57408 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624047346
transform -1 0 58880 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_624
timestamp 1624047346
transform 1 0 58512 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624047346
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output161
timestamp 1624047346
transform -1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output161_A
timestamp 1624047346
transform -1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1624047346
transform 1 0 1748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_13
timestamp 1624047346
transform 1 0 2300 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1624047346
transform 1 0 3404 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1624047346
transform 1 0 4508 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_49
timestamp 1624047346
transform 1 0 5612 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1624047346
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_58
timestamp 1624047346
transform 1 0 6440 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__S
timestamp 1624047346
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_70
timestamp 1624047346
transform 1 0 7544 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_84
timestamp 1624047346
transform 1 0 8832 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp 1624047346
transform 1 0 9200 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A0
timestamp 1624047346
transform 1 0 10396 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_97
timestamp 1624047346
transform 1 0 10028 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1624047346
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_103
timestamp 1624047346
transform 1 0 10580 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_111
timestamp 1624047346
transform 1 0 11316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_115
timestamp 1624047346
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_127
timestamp 1624047346
transform 1 0 12788 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_139
timestamp 1624047346
transform 1 0 13892 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_151
timestamp 1624047346
transform 1 0 14996 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_163
timestamp 1624047346
transform 1 0 16100 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1624047346
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_172
timestamp 1624047346
transform 1 0 16928 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1624047346
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1624047346
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1624047346
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1624047346
transform 1 0 22080 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_220
timestamp 1624047346
transform 1 0 21344 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_229
timestamp 1624047346
transform 1 0 22172 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_241
timestamp 1624047346
transform 1 0 23276 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_253
timestamp 1624047346
transform 1 0 24380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_265
timestamp 1624047346
transform 1 0 25484 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1624047346
transform 1 0 27324 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A
timestamp 1624047346
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_273
timestamp 1624047346
transform 1 0 26220 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_278
timestamp 1624047346
transform 1 0 26680 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_284
timestamp 1624047346
transform 1 0 27232 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_286
timestamp 1624047346
transform 1 0 27416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_298
timestamp 1624047346
transform 1 0 28520 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1624047346
transform 1 0 29624 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_322
timestamp 1624047346
transform 1 0 30728 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_334
timestamp 1624047346
transform 1 0 31832 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1624047346
transform 1 0 32568 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_343
timestamp 1624047346
transform 1 0 32660 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_355
timestamp 1624047346
transform 1 0 33764 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1624047346
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1624047346
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1624047346
transform 1 0 37812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_391
timestamp 1624047346
transform 1 0 37076 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_400
timestamp 1624047346
transform 1 0 37904 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_412
timestamp 1624047346
transform 1 0 39008 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_424
timestamp 1624047346
transform 1 0 40112 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_436
timestamp 1624047346
transform 1 0 41216 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_448
timestamp 1624047346
transform 1 0 42320 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1624047346
transform 1 0 43056 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_457
timestamp 1624047346
transform 1 0 43148 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_469
timestamp 1624047346
transform 1 0 44252 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_481
timestamp 1624047346
transform 1 0 45356 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_493
timestamp 1624047346
transform 1 0 46460 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1624047346
transform 1 0 47564 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1624047346
transform 1 0 48300 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_514
timestamp 1624047346
transform 1 0 48392 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_526
timestamp 1624047346
transform 1 0 49496 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_538
timestamp 1624047346
transform 1 0 50600 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_550
timestamp 1624047346
transform 1 0 51704 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1624047346
transform 1 0 53544 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_562
timestamp 1624047346
transform 1 0 52808 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_571
timestamp 1624047346
transform 1 0 53636 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_583
timestamp 1624047346
transform 1 0 54740 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_595
timestamp 1624047346
transform 1 0 55844 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output164
timestamp 1624047346
transform 1 0 57868 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output164_A
timestamp 1624047346
transform 1 0 57316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_607
timestamp 1624047346
transform 1 0 56948 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_613
timestamp 1624047346
transform 1 0 57500 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_621
timestamp 1624047346
transform 1 0 58236 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624047346
transform -1 0 58880 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624047346
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output234
timestamp 1624047346
transform -1 0 1748 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1624047346
transform 1 0 1748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1624047346
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_19
timestamp 1624047346
transform 1 0 2852 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624047346
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1624047346
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1624047346
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1624047346
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_66
timestamp 1624047346
transform 1 0 7176 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_78
timestamp 1624047346
transform 1 0 8280 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1624047346
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_87
timestamp 1624047346
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_99
timestamp 1624047346
transform 1 0 10212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_111
timestamp 1624047346
transform 1 0 11316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_123
timestamp 1624047346
transform 1 0 12420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1624047346
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_135
timestamp 1624047346
transform 1 0 13524 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_144
timestamp 1624047346
transform 1 0 14352 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_156
timestamp 1624047346
transform 1 0 15456 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_168
timestamp 1624047346
transform 1 0 16560 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_180
timestamp 1624047346
transform 1 0 17664 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1624047346
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_192
timestamp 1624047346
transform 1 0 18768 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1624047346
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_213
timestamp 1624047346
transform 1 0 20700 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_225
timestamp 1624047346
transform 1 0 21804 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_237
timestamp 1624047346
transform 1 0 22908 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_249
timestamp 1624047346
transform 1 0 24012 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1624047346
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_258
timestamp 1624047346
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_270
timestamp 1624047346
transform 1 0 25944 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_282
timestamp 1624047346
transform 1 0 27048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_294
timestamp 1624047346
transform 1 0 28152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1624047346
transform 1 0 29992 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_306
timestamp 1624047346
transform 1 0 29256 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_315
timestamp 1624047346
transform 1 0 30084 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_327
timestamp 1624047346
transform 1 0 31188 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_339
timestamp 1624047346
transform 1 0 32292 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_351
timestamp 1624047346
transform 1 0 33396 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_363
timestamp 1624047346
transform 1 0 34500 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1624047346
transform 1 0 35236 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_372
timestamp 1624047346
transform 1 0 35328 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_384
timestamp 1624047346
transform 1 0 36432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_396
timestamp 1624047346
transform 1 0 37536 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_408
timestamp 1624047346
transform 1 0 38640 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_420
timestamp 1624047346
transform 1 0 39744 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1624047346
transform 1 0 40480 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_429
timestamp 1624047346
transform 1 0 40572 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_441
timestamp 1624047346
transform 1 0 41676 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_453
timestamp 1624047346
transform 1 0 42780 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_465
timestamp 1624047346
transform 1 0 43884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1624047346
transform 1 0 45724 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_477
timestamp 1624047346
transform 1 0 44988 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_486
timestamp 1624047346
transform 1 0 45816 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_498
timestamp 1624047346
transform 1 0 46920 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_510
timestamp 1624047346
transform 1 0 48024 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_522
timestamp 1624047346
transform 1 0 49128 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_534
timestamp 1624047346
transform 1 0 50232 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1624047346
transform 1 0 50968 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_543
timestamp 1624047346
transform 1 0 51060 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_555
timestamp 1624047346
transform 1 0 52164 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_567
timestamp 1624047346
transform 1 0 53268 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_579
timestamp 1624047346
transform 1 0 54372 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1624047346
transform 1 0 56212 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_591
timestamp 1624047346
transform 1 0 55476 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_600
timestamp 1624047346
transform 1 0 56304 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_612
timestamp 1624047346
transform 1 0 57408 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624047346
transform -1 0 58880 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_624
timestamp 1624047346
transform 1 0 58512 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624047346
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624047346
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1624047346
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1624047346
transform -1 0 1564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_7
timestamp 1624047346
transform 1 0 1748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_5
timestamp 1624047346
transform 1 0 1564 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1624047346
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_19
timestamp 1624047346
transform 1 0 2852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_31
timestamp 1624047346
transform 1 0 3956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_17
timestamp 1624047346
transform 1 0 2668 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1624047346
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_43
timestamp 1624047346
transform 1 0 5060 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1624047346
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1624047346
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_55
timestamp 1624047346
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1624047346
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1624047346
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1624047346
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1624047346
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_82
timestamp 1624047346
transform 1 0 8648 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_78
timestamp 1624047346
transform 1 0 8280 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1624047346
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1624047346
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_87
timestamp 1624047346
transform 1 0 9108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_99
timestamp 1624047346
transform 1 0 10212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1624047346
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_106
timestamp 1624047346
transform 1 0 10856 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_115
timestamp 1624047346
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_111
timestamp 1624047346
transform 1 0 11316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_127
timestamp 1624047346
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_123
timestamp 1624047346
transform 1 0 12420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1624047346
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_139
timestamp 1624047346
transform 1 0 13892 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_151
timestamp 1624047346
transform 1 0 14996 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_135
timestamp 1624047346
transform 1 0 13524 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_144
timestamp 1624047346
transform 1 0 14352 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_163
timestamp 1624047346
transform 1 0 16100 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_156
timestamp 1624047346
transform 1 0 15456 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_168
timestamp 1624047346
transform 1 0 16560 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1624047346
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_172
timestamp 1624047346
transform 1 0 16928 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1624047346
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_180
timestamp 1624047346
transform 1 0 17664 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1624047346
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1624047346
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_192
timestamp 1624047346
transform 1 0 18768 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_201
timestamp 1624047346
transform 1 0 19596 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1624047346
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_213
timestamp 1624047346
transform 1 0 20700 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1624047346
transform 1 0 22080 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_220
timestamp 1624047346
transform 1 0 21344 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_229
timestamp 1624047346
transform 1 0 22172 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_225
timestamp 1624047346
transform 1 0 21804 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_241
timestamp 1624047346
transform 1 0 23276 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_237
timestamp 1624047346
transform 1 0 22908 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_249
timestamp 1624047346
transform 1 0 24012 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1624047346
transform 1 0 24748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_253
timestamp 1624047346
transform 1 0 24380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_265
timestamp 1624047346
transform 1 0 25484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_258
timestamp 1624047346
transform 1 0 24840 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1624047346
transform 1 0 27324 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_277
timestamp 1624047346
transform 1 0 26588 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_286
timestamp 1624047346
transform 1 0 27416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_270
timestamp 1624047346
transform 1 0 25944 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_282
timestamp 1624047346
transform 1 0 27048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_298
timestamp 1624047346
transform 1 0 28520 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_294
timestamp 1624047346
transform 1 0 28152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1624047346
transform 1 0 29992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_310
timestamp 1624047346
transform 1 0 29624 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_306
timestamp 1624047346
transform 1 0 29256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_315
timestamp 1624047346
transform 1 0 30084 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_322
timestamp 1624047346
transform 1 0 30728 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_334
timestamp 1624047346
transform 1 0 31832 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_327
timestamp 1624047346
transform 1 0 31188 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1624047346
transform 1 0 32568 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_343
timestamp 1624047346
transform 1 0 32660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_339
timestamp 1624047346
transform 1 0 32292 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_351
timestamp 1624047346
transform 1 0 33396 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _199_
timestamp 1624047346
transform 1 0 35144 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A
timestamp 1624047346
transform 1 0 34592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_355
timestamp 1624047346
transform 1 0 33764 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_363
timestamp 1624047346
transform 1 0 34500 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_366
timestamp 1624047346
transform 1 0 34776 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_363
timestamp 1624047346
transform 1 0 34500 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1624047346
transform 1 0 35236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_375
timestamp 1624047346
transform 1 0 35604 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_387
timestamp 1624047346
transform 1 0 36708 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_372
timestamp 1624047346
transform 1 0 35328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_384
timestamp 1624047346
transform 1 0 36432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1624047346
transform 1 0 37812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_400
timestamp 1624047346
transform 1 0 37904 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_396
timestamp 1624047346
transform 1 0 37536 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_412
timestamp 1624047346
transform 1 0 39008 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_408
timestamp 1624047346
transform 1 0 38640 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_420
timestamp 1624047346
transform 1 0 39744 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1624047346
transform 1 0 40480 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_424
timestamp 1624047346
transform 1 0 40112 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_436
timestamp 1624047346
transform 1 0 41216 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_429
timestamp 1624047346
transform 1 0 40572 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_448
timestamp 1624047346
transform 1 0 42320 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_441
timestamp 1624047346
transform 1 0 41676 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_453
timestamp 1624047346
transform 1 0 42780 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1624047346
transform 1 0 43056 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_457
timestamp 1624047346
transform 1 0 43148 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_469
timestamp 1624047346
transform 1 0 44252 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_465
timestamp 1624047346
transform 1 0 43884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1624047346
transform 1 0 45724 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_481
timestamp 1624047346
transform 1 0 45356 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_477
timestamp 1624047346
transform 1 0 44988 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_486
timestamp 1624047346
transform 1 0 45816 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_493
timestamp 1624047346
transform 1 0 46460 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1624047346
transform 1 0 47564 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_498
timestamp 1624047346
transform 1 0 46920 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1624047346
transform 1 0 48300 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_514
timestamp 1624047346
transform 1 0 48392 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_510
timestamp 1624047346
transform 1 0 48024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_526
timestamp 1624047346
transform 1 0 49496 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_538
timestamp 1624047346
transform 1 0 50600 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_522
timestamp 1624047346
transform 1 0 49128 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_534
timestamp 1624047346
transform 1 0 50232 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1624047346
transform 1 0 50968 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_550
timestamp 1624047346
transform 1 0 51704 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_543
timestamp 1624047346
transform 1 0 51060 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_555
timestamp 1624047346
transform 1 0 52164 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1624047346
transform 1 0 53544 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_562
timestamp 1624047346
transform 1 0 52808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_571
timestamp 1624047346
transform 1 0 53636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_567
timestamp 1624047346
transform 1 0 53268 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_583
timestamp 1624047346
transform 1 0 54740 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_579
timestamp 1624047346
transform 1 0 54372 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1624047346
transform 1 0 56212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_595
timestamp 1624047346
transform 1 0 55844 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_591
timestamp 1624047346
transform 1 0 55476 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_600
timestamp 1624047346
transform 1 0 56304 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_608
timestamp 1624047346
transform 1 0 57040 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_607
timestamp 1624047346
transform 1 0 56948 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_613
timestamp 1624047346
transform 1 0 57500 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_613
timestamp 1624047346
transform 1 0 57500 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output148_A
timestamp 1624047346
transform -1 0 57500 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1624047346
transform -1 0 57500 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output148
timestamp 1624047346
transform 1 0 57868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1624047346
transform 1 0 57868 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_621
timestamp 1624047346
transform 1 0 58236 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_621
timestamp 1624047346
transform 1 0 58236 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624047346
transform -1 0 58880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624047346
transform -1 0 58880 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624047346
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624047346
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624047346
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1624047346
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1624047346
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1624047346
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1624047346
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_58
timestamp 1624047346
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_70
timestamp 1624047346
transform 1 0 7544 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1624047346
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1624047346
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1624047346
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_106
timestamp 1624047346
transform 1 0 10856 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_115
timestamp 1624047346
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1624047346
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1624047346
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_151
timestamp 1624047346
transform 1 0 14996 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_163
timestamp 1624047346
transform 1 0 16100 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1624047346
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_172
timestamp 1624047346
transform 1 0 16928 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1624047346
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1624047346
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1624047346
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1624047346
transform 1 0 22080 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_220
timestamp 1624047346
transform 1 0 21344 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_229
timestamp 1624047346
transform 1 0 22172 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A
timestamp 1624047346
transform 1 0 23828 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_241
timestamp 1624047346
transform 1 0 23276 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1624047346
transform 1 0 24012 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _200_
timestamp 1624047346
transform -1 0 24840 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_15_258
timestamp 1624047346
transform 1 0 24840 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1624047346
transform 1 0 27324 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_270
timestamp 1624047346
transform 1 0 25944 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_282
timestamp 1624047346
transform 1 0 27048 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_286
timestamp 1624047346
transform 1 0 27416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_298
timestamp 1624047346
transform 1 0 28520 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_310
timestamp 1624047346
transform 1 0 29624 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_322
timestamp 1624047346
transform 1 0 30728 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_334
timestamp 1624047346
transform 1 0 31832 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1624047346
transform 1 0 32568 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_343
timestamp 1624047346
transform 1 0 32660 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_355
timestamp 1624047346
transform 1 0 33764 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1624047346
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1624047346
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1624047346
transform 1 0 37812 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_391
timestamp 1624047346
transform 1 0 37076 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_400
timestamp 1624047346
transform 1 0 37904 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_412
timestamp 1624047346
transform 1 0 39008 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_424
timestamp 1624047346
transform 1 0 40112 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_436
timestamp 1624047346
transform 1 0 41216 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_448
timestamp 1624047346
transform 1 0 42320 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1624047346
transform 1 0 43056 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_457
timestamp 1624047346
transform 1 0 43148 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_469
timestamp 1624047346
transform 1 0 44252 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_481
timestamp 1624047346
transform 1 0 45356 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_493
timestamp 1624047346
transform 1 0 46460 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_505
timestamp 1624047346
transform 1 0 47564 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1624047346
transform 1 0 48300 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_514
timestamp 1624047346
transform 1 0 48392 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_526
timestamp 1624047346
transform 1 0 49496 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_538
timestamp 1624047346
transform 1 0 50600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_550
timestamp 1624047346
transform 1 0 51704 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1624047346
transform 1 0 53544 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_562
timestamp 1624047346
transform 1 0 52808 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_571
timestamp 1624047346
transform 1 0 53636 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_583
timestamp 1624047346
transform 1 0 54740 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__S
timestamp 1624047346
transform 1 0 56764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_595
timestamp 1624047346
transform 1 0 55844 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_603
timestamp 1624047346
transform 1 0 56580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_607
timestamp 1624047346
transform 1 0 56948 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_619
timestamp 1624047346
transform 1 0 58052 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624047346
transform -1 0 58880 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624047346
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output188
timestamp 1624047346
transform -1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output188_A
timestamp 1624047346
transform -1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_7
timestamp 1624047346
transform 1 0 1748 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_13
timestamp 1624047346
transform 1 0 2300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1624047346
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_25
timestamp 1624047346
transform 1 0 3404 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624047346
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624047346
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_54
timestamp 1624047346
transform 1 0 6072 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_66
timestamp 1624047346
transform 1 0 7176 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_78
timestamp 1624047346
transform 1 0 8280 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1624047346
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_87
timestamp 1624047346
transform 1 0 9108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_99
timestamp 1624047346
transform 1 0 10212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_111
timestamp 1624047346
transform 1 0 11316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1624047346
transform 1 0 12420 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1624047346
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_135
timestamp 1624047346
transform 1 0 13524 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_144
timestamp 1624047346
transform 1 0 14352 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_156
timestamp 1624047346
transform 1 0 15456 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_168
timestamp 1624047346
transform 1 0 16560 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_180
timestamp 1624047346
transform 1 0 17664 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1624047346
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_192
timestamp 1624047346
transform 1 0 18768 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_201
timestamp 1624047346
transform 1 0 19596 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_213
timestamp 1624047346
transform 1 0 20700 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_225
timestamp 1624047346
transform 1 0 21804 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_237
timestamp 1624047346
transform 1 0 22908 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_249
timestamp 1624047346
transform 1 0 24012 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1624047346
transform 1 0 24748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_258
timestamp 1624047346
transform 1 0 24840 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_270
timestamp 1624047346
transform 1 0 25944 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_282
timestamp 1624047346
transform 1 0 27048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_294
timestamp 1624047346
transform 1 0 28152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1624047346
transform 1 0 29992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_306
timestamp 1624047346
transform 1 0 29256 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_315
timestamp 1624047346
transform 1 0 30084 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_327
timestamp 1624047346
transform 1 0 31188 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_339
timestamp 1624047346
transform 1 0 32292 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_351
timestamp 1624047346
transform 1 0 33396 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_363
timestamp 1624047346
transform 1 0 34500 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1624047346
transform 1 0 35236 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_372
timestamp 1624047346
transform 1 0 35328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_384
timestamp 1624047346
transform 1 0 36432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_396
timestamp 1624047346
transform 1 0 37536 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_408
timestamp 1624047346
transform 1 0 38640 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_420
timestamp 1624047346
transform 1 0 39744 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1624047346
transform 1 0 40480 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_429
timestamp 1624047346
transform 1 0 40572 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_441
timestamp 1624047346
transform 1 0 41676 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_453
timestamp 1624047346
transform 1 0 42780 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_465
timestamp 1624047346
transform 1 0 43884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1624047346
transform 1 0 45724 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_477
timestamp 1624047346
transform 1 0 44988 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_486
timestamp 1624047346
transform 1 0 45816 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_498
timestamp 1624047346
transform 1 0 46920 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_510
timestamp 1624047346
transform 1 0 48024 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_522
timestamp 1624047346
transform 1 0 49128 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_534
timestamp 1624047346
transform 1 0 50232 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1624047346
transform 1 0 50968 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_543
timestamp 1624047346
transform 1 0 51060 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_555
timestamp 1624047346
transform 1 0 52164 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_567
timestamp 1624047346
transform 1 0 53268 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_579
timestamp 1624047346
transform 1 0 54372 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1624047346
transform 1 0 56212 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A1
timestamp 1624047346
transform 1 0 56580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_591
timestamp 1624047346
transform 1 0 55476 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_600
timestamp 1624047346
transform 1 0 56304 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_605
timestamp 1624047346
transform 1 0 56764 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _263_
timestamp 1624047346
transform -1 0 57960 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_16_618
timestamp 1624047346
transform 1 0 57960 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624047346
transform -1 0 58880 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_624
timestamp 1624047346
transform 1 0 58512 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624047346
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1624047346
transform -1 0 1748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output127_A
timestamp 1624047346
transform -1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1624047346
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_13
timestamp 1624047346
transform 1 0 2300 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_25
timestamp 1624047346
transform 1 0 3404 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_37
timestamp 1624047346
transform 1 0 4508 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_49
timestamp 1624047346
transform 1 0 5612 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1624047346
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1624047346
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_70
timestamp 1624047346
transform 1 0 7544 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_82
timestamp 1624047346
transform 1 0 8648 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_94
timestamp 1624047346
transform 1 0 9752 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1624047346
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_106
timestamp 1624047346
transform 1 0 10856 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_115
timestamp 1624047346
transform 1 0 11684 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_127
timestamp 1624047346
transform 1 0 12788 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_139
timestamp 1624047346
transform 1 0 13892 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_151
timestamp 1624047346
transform 1 0 14996 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_163
timestamp 1624047346
transform 1 0 16100 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1624047346
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_172
timestamp 1624047346
transform 1 0 16928 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1624047346
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1624047346
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1624047346
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1624047346
transform 1 0 22080 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_220
timestamp 1624047346
transform 1 0 21344 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1624047346
transform 1 0 22172 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_241
timestamp 1624047346
transform 1 0 23276 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_253
timestamp 1624047346
transform 1 0 24380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_265
timestamp 1624047346
transform 1 0 25484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1624047346
transform 1 0 27324 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_277
timestamp 1624047346
transform 1 0 26588 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_286
timestamp 1624047346
transform 1 0 27416 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_298
timestamp 1624047346
transform 1 0 28520 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_310
timestamp 1624047346
transform 1 0 29624 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_322
timestamp 1624047346
transform 1 0 30728 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_334
timestamp 1624047346
transform 1 0 31832 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1624047346
transform 1 0 32568 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_343
timestamp 1624047346
transform 1 0 32660 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_355
timestamp 1624047346
transform 1 0 33764 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1624047346
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1624047346
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1624047346
transform 1 0 37812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_391
timestamp 1624047346
transform 1 0 37076 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_400
timestamp 1624047346
transform 1 0 37904 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_412
timestamp 1624047346
transform 1 0 39008 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_424
timestamp 1624047346
transform 1 0 40112 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_436
timestamp 1624047346
transform 1 0 41216 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_448
timestamp 1624047346
transform 1 0 42320 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1624047346
transform 1 0 43056 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_457
timestamp 1624047346
transform 1 0 43148 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_469
timestamp 1624047346
transform 1 0 44252 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_481
timestamp 1624047346
transform 1 0 45356 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_493
timestamp 1624047346
transform 1 0 46460 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1624047346
transform 1 0 47564 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1624047346
transform 1 0 48300 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_514
timestamp 1624047346
transform 1 0 48392 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_526
timestamp 1624047346
transform 1 0 49496 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_538
timestamp 1624047346
transform 1 0 50600 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_550
timestamp 1624047346
transform 1 0 51704 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1624047346
transform 1 0 53544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_562
timestamp 1624047346
transform 1 0 52808 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_571
timestamp 1624047346
transform 1 0 53636 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_583
timestamp 1624047346
transform 1 0 54740 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_595
timestamp 1624047346
transform 1 0 55844 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output215
timestamp 1624047346
transform 1 0 57868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_607
timestamp 1624047346
transform 1 0 56948 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_615
timestamp 1624047346
transform 1 0 57684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1624047346
transform 1 0 58236 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624047346
transform -1 0 58880 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624047346
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624047346
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624047346
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1624047346
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624047346
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1624047346
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1624047346
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_54
timestamp 1624047346
transform 1 0 6072 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_66
timestamp 1624047346
transform 1 0 7176 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_78
timestamp 1624047346
transform 1 0 8280 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1624047346
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_87
timestamp 1624047346
transform 1 0 9108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1624047346
transform 1 0 10212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_111
timestamp 1624047346
transform 1 0 11316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_123
timestamp 1624047346
transform 1 0 12420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1624047346
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_135
timestamp 1624047346
transform 1 0 13524 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_144
timestamp 1624047346
transform 1 0 14352 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_156
timestamp 1624047346
transform 1 0 15456 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_168
timestamp 1624047346
transform 1 0 16560 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_180
timestamp 1624047346
transform 1 0 17664 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1624047346
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_192
timestamp 1624047346
transform 1 0 18768 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1624047346
transform 1 0 19596 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_213
timestamp 1624047346
transform 1 0 20700 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_225
timestamp 1624047346
transform 1 0 21804 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_237
timestamp 1624047346
transform 1 0 22908 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_249
timestamp 1624047346
transform 1 0 24012 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1624047346
transform 1 0 24748 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_258
timestamp 1624047346
transform 1 0 24840 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_270
timestamp 1624047346
transform 1 0 25944 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_282
timestamp 1624047346
transform 1 0 27048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_294
timestamp 1624047346
transform 1 0 28152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1624047346
transform 1 0 29992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_306
timestamp 1624047346
transform 1 0 29256 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_315
timestamp 1624047346
transform 1 0 30084 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_327
timestamp 1624047346
transform 1 0 31188 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_339
timestamp 1624047346
transform 1 0 32292 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_351
timestamp 1624047346
transform 1 0 33396 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_363
timestamp 1624047346
transform 1 0 34500 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1624047346
transform 1 0 35236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_372
timestamp 1624047346
transform 1 0 35328 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_384
timestamp 1624047346
transform 1 0 36432 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_396
timestamp 1624047346
transform 1 0 37536 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_408
timestamp 1624047346
transform 1 0 38640 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_420
timestamp 1624047346
transform 1 0 39744 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1624047346
transform 1 0 40480 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_429
timestamp 1624047346
transform 1 0 40572 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_441
timestamp 1624047346
transform 1 0 41676 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_453
timestamp 1624047346
transform 1 0 42780 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_465
timestamp 1624047346
transform 1 0 43884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1624047346
transform 1 0 45724 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1624047346
transform 1 0 44988 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_486
timestamp 1624047346
transform 1 0 45816 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_498
timestamp 1624047346
transform 1 0 46920 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_510
timestamp 1624047346
transform 1 0 48024 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_522
timestamp 1624047346
transform 1 0 49128 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_534
timestamp 1624047346
transform 1 0 50232 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1624047346
transform 1 0 50968 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_543
timestamp 1624047346
transform 1 0 51060 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_555
timestamp 1624047346
transform 1 0 52164 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_567
timestamp 1624047346
transform 1 0 53268 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_579
timestamp 1624047346
transform 1 0 54372 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1624047346
transform 1 0 56212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_591
timestamp 1624047346
transform 1 0 55476 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_600
timestamp 1624047346
transform 1 0 56304 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input67
timestamp 1624047346
transform -1 0 58236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1624047346
transform -1 0 57500 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_608
timestamp 1624047346
transform 1 0 57040 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_613
timestamp 1624047346
transform 1 0 57500 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_621
timestamp 1624047346
transform 1 0 58236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624047346
transform -1 0 58880 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1624047346
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624047346
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624047346
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output230
timestamp 1624047346
transform -1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__S
timestamp 1624047346
transform -1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1624047346
transform -1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1624047346
transform 1 0 1748 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_13
timestamp 1624047346
transform 1 0 2300 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_5
timestamp 1624047346
transform 1 0 1564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1624047346
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A0
timestamp 1624047346
transform -1 0 3312 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1624047346
transform 1 0 3404 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_18
timestamp 1624047346
transform 1 0 2760 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1624047346
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_28
timestamp 1624047346
transform 1 0 3680 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1624047346
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1624047346
transform 1 0 4508 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_49
timestamp 1624047346
transform 1 0 5612 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1624047346
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1624047346
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_58
timestamp 1624047346
transform 1 0 6440 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_54
timestamp 1624047346
transform 1 0 6072 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_66
timestamp 1624047346
transform 1 0 7176 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_70
timestamp 1624047346
transform 1 0 7544 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_82
timestamp 1624047346
transform 1 0 8648 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_78
timestamp 1624047346
transform 1 0 8280 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _082_
timestamp 1624047346
transform -1 0 10580 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1624047346
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_94
timestamp 1624047346
transform 1 0 9752 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_87
timestamp 1624047346
transform 1 0 9108 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_95
timestamp 1624047346
transform 1 0 9844 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_103
timestamp 1624047346
transform 1 0 10580 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_102
timestamp 1624047346
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1624047346
transform -1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _081_
timestamp 1624047346
transform -1 0 11408 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_112
timestamp 1624047346
transform 1 0 11408 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1624047346
transform 1 0 11500 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1624047346
transform 1 0 11776 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1624047346
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_115
timestamp 1624047346
transform 1 0 11684 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_105
timestamp 1624047346
transform 1 0 10764 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _088_
timestamp 1624047346
transform -1 0 13064 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1624047346
transform 1 0 13432 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1624047346
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_118
timestamp 1624047346
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_124
timestamp 1624047346
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_130
timestamp 1624047346
transform 1 0 13064 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1624047346
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_139
timestamp 1624047346
transform 1 0 13892 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_151
timestamp 1624047346
transform 1 0 14996 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_136
timestamp 1624047346
transform 1 0 13616 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_142
timestamp 1624047346
transform 1 0 14168 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_144
timestamp 1624047346
transform 1 0 14352 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_163
timestamp 1624047346
transform 1 0 16100 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_156
timestamp 1624047346
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_168
timestamp 1624047346
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1624047346
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_172
timestamp 1624047346
transform 1 0 16928 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1624047346
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1624047346
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1624047346
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1624047346
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1624047346
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_201
timestamp 1624047346
transform 1 0 19596 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1624047346
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1624047346
transform 1 0 20700 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1624047346
transform 1 0 22080 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_220
timestamp 1624047346
transform 1 0 21344 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_229
timestamp 1624047346
transform 1 0 22172 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_225
timestamp 1624047346
transform 1 0 21804 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_241
timestamp 1624047346
transform 1 0 23276 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1624047346
transform 1 0 22908 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_249
timestamp 1624047346
transform 1 0 24012 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1624047346
transform 1 0 24748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_253
timestamp 1624047346
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_265
timestamp 1624047346
transform 1 0 25484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_258
timestamp 1624047346
transform 1 0 24840 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1624047346
transform 1 0 27324 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_277
timestamp 1624047346
transform 1 0 26588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_286
timestamp 1624047346
transform 1 0 27416 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_270
timestamp 1624047346
transform 1 0 25944 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_282
timestamp 1624047346
transform 1 0 27048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_298
timestamp 1624047346
transform 1 0 28520 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_294
timestamp 1624047346
transform 1 0 28152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1624047346
transform 1 0 29992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_310
timestamp 1624047346
transform 1 0 29624 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_306
timestamp 1624047346
transform 1 0 29256 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_315
timestamp 1624047346
transform 1 0 30084 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_322
timestamp 1624047346
transform 1 0 30728 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_334
timestamp 1624047346
transform 1 0 31832 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_327
timestamp 1624047346
transform 1 0 31188 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1624047346
transform 1 0 32568 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_343
timestamp 1624047346
transform 1 0 32660 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_339
timestamp 1624047346
transform 1 0 32292 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_351
timestamp 1624047346
transform 1 0 33396 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_355
timestamp 1624047346
transform 1 0 33764 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1624047346
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_363
timestamp 1624047346
transform 1 0 34500 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1624047346
transform 1 0 35236 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1624047346
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_372
timestamp 1624047346
transform 1 0 35328 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_384
timestamp 1624047346
transform 1 0 36432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1624047346
transform 1 0 37812 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_391
timestamp 1624047346
transform 1 0 37076 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_400
timestamp 1624047346
transform 1 0 37904 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_396
timestamp 1624047346
transform 1 0 37536 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_412
timestamp 1624047346
transform 1 0 39008 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_408
timestamp 1624047346
transform 1 0 38640 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_420
timestamp 1624047346
transform 1 0 39744 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1624047346
transform 1 0 40480 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_424
timestamp 1624047346
transform 1 0 40112 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_436
timestamp 1624047346
transform 1 0 41216 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_429
timestamp 1624047346
transform 1 0 40572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_448
timestamp 1624047346
transform 1 0 42320 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_441
timestamp 1624047346
transform 1 0 41676 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_453
timestamp 1624047346
transform 1 0 42780 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1624047346
transform 1 0 43056 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_457
timestamp 1624047346
transform 1 0 43148 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_469
timestamp 1624047346
transform 1 0 44252 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_465
timestamp 1624047346
transform 1 0 43884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1624047346
transform 1 0 45724 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_481
timestamp 1624047346
transform 1 0 45356 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_477
timestamp 1624047346
transform 1 0 44988 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_486
timestamp 1624047346
transform 1 0 45816 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_493
timestamp 1624047346
transform 1 0 46460 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1624047346
transform 1 0 47564 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_498
timestamp 1624047346
transform 1 0 46920 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1624047346
transform 1 0 48300 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_514
timestamp 1624047346
transform 1 0 48392 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_510
timestamp 1624047346
transform 1 0 48024 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_526
timestamp 1624047346
transform 1 0 49496 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_538
timestamp 1624047346
transform 1 0 50600 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_522
timestamp 1624047346
transform 1 0 49128 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_534
timestamp 1624047346
transform 1 0 50232 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1624047346
transform 1 0 50968 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_550
timestamp 1624047346
transform 1 0 51704 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_543
timestamp 1624047346
transform 1 0 51060 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_555
timestamp 1624047346
transform 1 0 52164 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1624047346
transform 1 0 53544 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_562
timestamp 1624047346
transform 1 0 52808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_571
timestamp 1624047346
transform 1 0 53636 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_567
timestamp 1624047346
transform 1 0 53268 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_583
timestamp 1624047346
transform 1 0 54740 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_579
timestamp 1624047346
transform 1 0 54372 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1624047346
transform 1 0 56212 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_595
timestamp 1624047346
transform 1 0 55844 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_591
timestamp 1624047346
transform 1 0 55476 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_600
timestamp 1624047346
transform 1 0 56304 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input102
timestamp 1624047346
transform -1 0 58236 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1624047346
transform -1 0 57500 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_607
timestamp 1624047346
transform 1 0 56948 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_613
timestamp 1624047346
transform 1 0 57500 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_621
timestamp 1624047346
transform 1 0 58236 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_612
timestamp 1624047346
transform 1 0 57408 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624047346
transform -1 0 58880 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624047346
transform -1 0 58880 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_624
timestamp 1624047346
transform 1 0 58512 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624047346
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1624047346
transform -1 0 1656 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624047346
transform -1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_6
timestamp 1624047346
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_12
timestamp 1624047346
transform 1 0 2208 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_24
timestamp 1624047346
transform 1 0 3312 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_36
timestamp 1624047346
transform 1 0 4416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_48
timestamp 1624047346
transform 1 0 5520 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1624047346
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_56
timestamp 1624047346
transform 1 0 6256 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_58
timestamp 1624047346
transform 1 0 6440 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_70
timestamp 1624047346
transform 1 0 7544 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_82
timestamp 1624047346
transform 1 0 8648 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _188_
timestamp 1624047346
transform -1 0 10856 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_21_94
timestamp 1624047346
transform 1 0 9752 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_100
timestamp 1624047346
transform 1 0 10304 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1624047346
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1624047346
transform 1 0 11684 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_106
timestamp 1624047346
transform 1 0 10856 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_117
timestamp 1624047346
transform 1 0 11868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _191_
timestamp 1624047346
transform 1 0 13432 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_21_129
timestamp 1624047346
transform 1 0 12972 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_133
timestamp 1624047346
transform 1 0 13340 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__191__A
timestamp 1624047346
transform 1 0 14260 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_139
timestamp 1624047346
transform 1 0 13892 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_145
timestamp 1624047346
transform 1 0 14444 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_157
timestamp 1624047346
transform 1 0 15548 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1624047346
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1624047346
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_172
timestamp 1624047346
transform 1 0 16928 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1624047346
transform 1 0 18032 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1624047346
transform 1 0 19136 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1624047346
transform 1 0 20240 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _106_
timestamp 1624047346
transform -1 0 23092 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1624047346
transform 1 0 22080 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_220
timestamp 1624047346
transform 1 0 21344 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_229
timestamp 1624047346
transform 1 0 22172 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_233
timestamp 1624047346
transform 1 0 22540 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1624047346
transform 1 0 23460 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_239
timestamp 1624047346
transform 1 0 23092 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1624047346
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1624047346
transform 1 0 24748 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1624047346
transform 1 0 25852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1624047346
transform 1 0 27324 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1624047346
transform 1 0 26956 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_286
timestamp 1624047346
transform 1 0 27416 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_298
timestamp 1624047346
transform 1 0 28520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_310
timestamp 1624047346
transform 1 0 29624 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_322
timestamp 1624047346
transform 1 0 30728 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_334
timestamp 1624047346
transform 1 0 31832 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1624047346
transform 1 0 32568 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_343
timestamp 1624047346
transform 1 0 32660 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _100_
timestamp 1624047346
transform -1 0 35972 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1624047346
transform 1 0 34592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_355
timestamp 1624047346
transform 1 0 33764 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_363
timestamp 1624047346
transform 1 0 34500 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_366
timestamp 1624047346
transform 1 0 34776 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1624047346
transform 1 0 35972 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1624047346
transform 1 0 37812 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_391
timestamp 1624047346
transform 1 0 37076 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_400
timestamp 1624047346
transform 1 0 37904 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_412
timestamp 1624047346
transform 1 0 39008 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_424
timestamp 1624047346
transform 1 0 40112 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_436
timestamp 1624047346
transform 1 0 41216 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_448
timestamp 1624047346
transform 1 0 42320 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1624047346
transform 1 0 43056 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_457
timestamp 1624047346
transform 1 0 43148 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_469
timestamp 1624047346
transform 1 0 44252 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_481
timestamp 1624047346
transform 1 0 45356 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_493
timestamp 1624047346
transform 1 0 46460 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_505
timestamp 1624047346
transform 1 0 47564 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1624047346
transform 1 0 48300 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_514
timestamp 1624047346
transform 1 0 48392 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_526
timestamp 1624047346
transform 1 0 49496 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_538
timestamp 1624047346
transform 1 0 50600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_550
timestamp 1624047346
transform 1 0 51704 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1624047346
transform 1 0 53544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_562
timestamp 1624047346
transform 1 0 52808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_571
timestamp 1624047346
transform 1 0 53636 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_583
timestamp 1624047346
transform 1 0 54740 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_595
timestamp 1624047346
transform 1 0 55844 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_607
timestamp 1624047346
transform 1 0 56948 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_619
timestamp 1624047346
transform 1 0 58052 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624047346
transform -1 0 58880 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624047346
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624047346
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624047346
transform -1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1624047346
transform 1 0 1656 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_12
timestamp 1624047346
transform 1 0 2208 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1624047346
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1624047346
transform 1 0 3312 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_28
timestamp 1624047346
transform 1 0 3680 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1624047346
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_42
timestamp 1624047346
transform 1 0 4968 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_54
timestamp 1624047346
transform 1 0 6072 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_66
timestamp 1624047346
transform 1 0 7176 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_78
timestamp 1624047346
transform 1 0 8280 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1624047346
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_87
timestamp 1624047346
transform 1 0 9108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_99
timestamp 1624047346
transform 1 0 10212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_111
timestamp 1624047346
transform 1 0 11316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_123
timestamp 1624047346
transform 1 0 12420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1624047346
transform -1 0 14996 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1624047346
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1624047346
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_144
timestamp 1624047346
transform 1 0 14352 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_151
timestamp 1624047346
transform 1 0 14996 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1624047346
transform -1 0 15548 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_157
timestamp 1624047346
transform 1 0 15548 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_169
timestamp 1624047346
transform 1 0 16652 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_181
timestamp 1624047346
transform 1 0 17756 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1624047346
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_193
timestamp 1624047346
transform 1 0 18860 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_199
timestamp 1624047346
transform 1 0 19412 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_201
timestamp 1624047346
transform 1 0 19596 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_213
timestamp 1624047346
transform 1 0 20700 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp 1624047346
transform 1 0 22448 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_225
timestamp 1624047346
transform 1 0 21804 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_231
timestamp 1624047346
transform 1 0 22356 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_235
timestamp 1624047346
transform 1 0 22724 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _098_
timestamp 1624047346
transform -1 0 23828 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_247
timestamp 1624047346
transform 1 0 23828 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1624047346
transform 1 0 24748 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_255
timestamp 1624047346
transform 1 0 24564 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_258
timestamp 1624047346
transform 1 0 24840 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_270
timestamp 1624047346
transform 1 0 25944 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_282
timestamp 1624047346
transform 1 0 27048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_294
timestamp 1624047346
transform 1 0 28152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1624047346
transform 1 0 29992 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_306
timestamp 1624047346
transform 1 0 29256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_315
timestamp 1624047346
transform 1 0 30084 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_327
timestamp 1624047346
transform 1 0 31188 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_339
timestamp 1624047346
transform 1 0 32292 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_351
timestamp 1624047346
transform 1 0 33396 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_363
timestamp 1624047346
transform 1 0 34500 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1624047346
transform 1 0 35236 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_372
timestamp 1624047346
transform 1 0 35328 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_384
timestamp 1624047346
transform 1 0 36432 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp 1624047346
transform -1 0 37168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_388
timestamp 1624047346
transform 1 0 36800 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_392
timestamp 1624047346
transform 1 0 37168 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_404
timestamp 1624047346
transform 1 0 38272 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_416
timestamp 1624047346
transform 1 0 39376 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1624047346
transform 1 0 40480 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_429
timestamp 1624047346
transform 1 0 40572 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_441
timestamp 1624047346
transform 1 0 41676 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_453
timestamp 1624047346
transform 1 0 42780 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_465
timestamp 1624047346
transform 1 0 43884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1624047346
transform 1 0 45724 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_477
timestamp 1624047346
transform 1 0 44988 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_486
timestamp 1624047346
transform 1 0 45816 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_498
timestamp 1624047346
transform 1 0 46920 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_510
timestamp 1624047346
transform 1 0 48024 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_522
timestamp 1624047346
transform 1 0 49128 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_534
timestamp 1624047346
transform 1 0 50232 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1624047346
transform 1 0 50968 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__S
timestamp 1624047346
transform 1 0 51888 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_543
timestamp 1624047346
transform 1 0 51060 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_551
timestamp 1624047346
transform 1 0 51796 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_554
timestamp 1624047346
transform 1 0 52072 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _257_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 53544 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_570
timestamp 1624047346
transform 1 0 53544 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_582
timestamp 1624047346
transform 1 0 54648 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1624047346
transform 1 0 56212 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_594
timestamp 1624047346
transform 1 0 55752 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_598
timestamp 1624047346
transform 1 0 56120 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_600
timestamp 1624047346
transform 1 0 56304 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1624047346
transform 1 0 57960 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624047346
transform -1 0 57592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_614
timestamp 1624047346
transform 1 0 57592 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1624047346
transform 1 0 58236 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624047346
transform -1 0 58880 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624047346
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624047346
transform -1 0 1564 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_5
timestamp 1624047346
transform 1 0 1564 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_17
timestamp 1624047346
transform 1 0 2668 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_29
timestamp 1624047346
transform 1 0 3772 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_41
timestamp 1624047346
transform 1 0 4876 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1624047346
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_53
timestamp 1624047346
transform 1 0 5980 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_58
timestamp 1624047346
transform 1 0 6440 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_70
timestamp 1624047346
transform 1 0 7544 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_82
timestamp 1624047346
transform 1 0 8648 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_94
timestamp 1624047346
transform 1 0 9752 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1624047346
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_106
timestamp 1624047346
transform 1 0 10856 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_115
timestamp 1624047346
transform 1 0 11684 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_127
timestamp 1624047346
transform 1 0 12788 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_139
timestamp 1624047346
transform 1 0 13892 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_151
timestamp 1624047346
transform 1 0 14996 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_163
timestamp 1624047346
transform 1 0 16100 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _111_
timestamp 1624047346
transform 1 0 17572 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1624047346
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_172
timestamp 1624047346
transform 1 0 16928 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_178
timestamp 1624047346
transform 1 0 17480 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__B
timestamp 1624047346
transform -1 0 18952 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_188
timestamp 1624047346
transform 1 0 18400 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_194
timestamp 1624047346
transform 1 0 18952 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_206
timestamp 1624047346
transform 1 0 20056 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_218
timestamp 1624047346
transform 1 0 21160 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1624047346
transform 1 0 22080 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_226
timestamp 1624047346
transform 1 0 21896 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_229
timestamp 1624047346
transform 1 0 22172 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_241
timestamp 1624047346
transform 1 0 23276 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_253
timestamp 1624047346
transform 1 0 24380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_265
timestamp 1624047346
transform 1 0 25484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1624047346
transform 1 0 27324 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_277
timestamp 1624047346
transform 1 0 26588 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_286
timestamp 1624047346
transform 1 0 27416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_298
timestamp 1624047346
transform 1 0 28520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_310
timestamp 1624047346
transform 1 0 29624 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_322
timestamp 1624047346
transform 1 0 30728 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_334
timestamp 1624047346
transform 1 0 31832 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1624047346
transform 1 0 32568 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_343
timestamp 1624047346
transform 1 0 32660 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_355
timestamp 1624047346
transform 1 0 33764 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1624047346
transform 1 0 34868 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _246_
timestamp 1624047346
transform -1 0 37076 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_23_379
timestamp 1624047346
transform 1 0 35972 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_385
timestamp 1624047346
transform 1 0 36524 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1624047346
transform 1 0 37812 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_391
timestamp 1624047346
transform 1 0 37076 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_400
timestamp 1624047346
transform 1 0 37904 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_412
timestamp 1624047346
transform 1 0 39008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_424
timestamp 1624047346
transform 1 0 40112 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_436
timestamp 1624047346
transform 1 0 41216 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_448
timestamp 1624047346
transform 1 0 42320 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1624047346
transform 1 0 43056 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_457
timestamp 1624047346
transform 1 0 43148 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_469
timestamp 1624047346
transform 1 0 44252 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_481
timestamp 1624047346
transform 1 0 45356 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_493
timestamp 1624047346
transform 1 0 46460 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_505
timestamp 1624047346
transform 1 0 47564 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1624047346
transform 1 0 48300 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_514
timestamp 1624047346
transform 1 0 48392 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_526
timestamp 1624047346
transform 1 0 49496 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_538
timestamp 1624047346
transform 1 0 50600 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_550
timestamp 1624047346
transform 1 0 51704 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1624047346
transform 1 0 53544 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_562
timestamp 1624047346
transform 1 0 52808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_571
timestamp 1624047346
transform 1 0 53636 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_583
timestamp 1624047346
transform 1 0 54740 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_595
timestamp 1624047346
transform 1 0 55844 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1624047346
transform -1 0 58236 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1624047346
transform -1 0 57500 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_607
timestamp 1624047346
transform 1 0 56948 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_613
timestamp 1624047346
transform 1 0 57500 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_621
timestamp 1624047346
transform 1 0 58236 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624047346
transform -1 0 58880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624047346
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1624047346
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_7
timestamp 1624047346
transform 1 0 1748 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1624047346
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_19
timestamp 1624047346
transform 1 0 2852 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1624047346
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1624047346
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_42
timestamp 1624047346
transform 1 0 4968 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_54
timestamp 1624047346
transform 1 0 6072 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_66
timestamp 1624047346
transform 1 0 7176 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_78
timestamp 1624047346
transform 1 0 8280 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1624047346
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_87
timestamp 1624047346
transform 1 0 9108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_99
timestamp 1624047346
transform 1 0 10212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_111
timestamp 1624047346
transform 1 0 11316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_123
timestamp 1624047346
transform 1 0 12420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1624047346
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_135
timestamp 1624047346
transform 1 0 13524 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_144
timestamp 1624047346
transform 1 0 14352 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_156
timestamp 1624047346
transform 1 0 15456 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_168
timestamp 1624047346
transform 1 0 16560 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _113_
timestamp 1624047346
transform -1 0 18032 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_24_176
timestamp 1624047346
transform 1 0 17296 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_184
timestamp 1624047346
transform 1 0 18032 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1624047346
transform 1 0 18768 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1624047346
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_196
timestamp 1624047346
transform 1 0 19136 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_201
timestamp 1624047346
transform 1 0 19596 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_213
timestamp 1624047346
transform 1 0 20700 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _202_
timestamp 1624047346
transform -1 0 22264 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_221
timestamp 1624047346
transform 1 0 21436 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_230
timestamp 1624047346
transform 1 0 22264 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_242
timestamp 1624047346
transform 1 0 23368 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 25208 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1624047346
transform 1 0 24748 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_254
timestamp 1624047346
transform 1 0 24472 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1624047346
transform 1 0 24840 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_268
timestamp 1624047346
transform 1 0 25760 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_280
timestamp 1624047346
transform 1 0 26864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1624047346
transform 1 0 28428 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_292
timestamp 1624047346
transform 1 0 27968 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_296
timestamp 1624047346
transform 1 0 28336 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_300
timestamp 1624047346
transform 1 0 28704 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1624047346
transform 1 0 29992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1624047346
transform -1 0 29256 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_306
timestamp 1624047346
transform 1 0 29256 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_315
timestamp 1624047346
transform 1 0 30084 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_327
timestamp 1624047346
transform 1 0 31188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _206_
timestamp 1624047346
transform 1 0 32844 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A
timestamp 1624047346
transform 1 0 32292 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_341
timestamp 1624047346
transform 1 0 32476 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_350
timestamp 1624047346
transform 1 0 33304 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__B
timestamp 1624047346
transform 1 0 33672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_356
timestamp 1624047346
transform 1 0 33856 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_368
timestamp 1624047346
transform 1 0 34960 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1624047346
transform 1 0 35236 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1624047346
transform -1 0 36248 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_372
timestamp 1624047346
transform 1 0 35328 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_382
timestamp 1624047346
transform 1 0 36248 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 1624047346
transform 1 0 37628 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__A
timestamp 1624047346
transform -1 0 37260 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_390
timestamp 1624047346
transform 1 0 36984 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_393
timestamp 1624047346
transform 1 0 37260 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_400
timestamp 1624047346
transform 1 0 37904 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_404
timestamp 1624047346
transform 1 0 38272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _249_
timestamp 1624047346
transform -1 0 39192 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_24_414
timestamp 1624047346
transform 1 0 39192 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _152_
timestamp 1624047346
transform 1 0 40940 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1624047346
transform 1 0 40480 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_426
timestamp 1624047346
transform 1 0 40296 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_429
timestamp 1624047346
transform 1 0 40572 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_442
timestamp 1624047346
transform 1 0 41768 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_454
timestamp 1624047346
transform 1 0 42872 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_466
timestamp 1624047346
transform 1 0 43976 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1624047346
transform 1 0 45724 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_478
timestamp 1624047346
transform 1 0 45080 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_484
timestamp 1624047346
transform 1 0 45632 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_486
timestamp 1624047346
transform 1 0 45816 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_498
timestamp 1624047346
transform 1 0 46920 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_510
timestamp 1624047346
transform 1 0 48024 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_522
timestamp 1624047346
transform 1 0 49128 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_534
timestamp 1624047346
transform 1 0 50232 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1624047346
transform 1 0 50968 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_543
timestamp 1624047346
transform 1 0 51060 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_555
timestamp 1624047346
transform 1 0 52164 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_567
timestamp 1624047346
transform 1 0 53268 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_579
timestamp 1624047346
transform 1 0 54372 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1624047346
transform 1 0 56212 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_591
timestamp 1624047346
transform 1 0 55476 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_600
timestamp 1624047346
transform 1 0 56304 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_612
timestamp 1624047346
transform 1 0 57408 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624047346
transform -1 0 58880 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_624
timestamp 1624047346
transform 1 0 58512 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624047346
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1624047346
transform -1 0 1564 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_5
timestamp 1624047346
transform 1 0 1564 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_17
timestamp 1624047346
transform 1 0 2668 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_29
timestamp 1624047346
transform 1 0 3772 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_41
timestamp 1624047346
transform 1 0 4876 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1624047346
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_53
timestamp 1624047346
transform 1 0 5980 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_58
timestamp 1624047346
transform 1 0 6440 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _095_
timestamp 1624047346
transform -1 0 8832 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_25_70
timestamp 1624047346
transform 1 0 7544 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_78
timestamp 1624047346
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_84
timestamp 1624047346
transform 1 0 8832 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1624047346
transform -1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_90
timestamp 1624047346
transform 1 0 9384 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1624047346
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_102
timestamp 1624047346
transform 1 0 10488 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_115
timestamp 1624047346
transform 1 0 11684 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_127
timestamp 1624047346
transform 1 0 12788 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_139
timestamp 1624047346
transform 1 0 13892 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_151
timestamp 1624047346
transform 1 0 14996 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_163
timestamp 1624047346
transform 1 0 16100 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1624047346
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_172
timestamp 1624047346
transform 1 0 16928 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1624047346
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1624047346
transform -1 0 18584 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_190
timestamp 1624047346
transform 1 0 18584 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_202
timestamp 1624047346
transform 1 0 19688 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _187_
timestamp 1624047346
transform -1 0 21436 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_214
timestamp 1624047346
transform 1 0 20792 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1624047346
transform 1 0 22080 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__A
timestamp 1624047346
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_221
timestamp 1624047346
transform 1 0 21436 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_227
timestamp 1624047346
transform 1 0 21988 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_229
timestamp 1624047346
transform 1 0 22172 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_234
timestamp 1624047346
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _204_
timestamp 1624047346
transform -1 0 23828 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_25_247
timestamp 1624047346
transform 1 0 23828 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  _209_
timestamp 1624047346
transform -1 0 26404 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_259
timestamp 1624047346
transform 1 0 24932 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_267
timestamp 1624047346
transform 1 0 25668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1624047346
transform 1 0 27324 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_275
timestamp 1624047346
transform 1 0 26404 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_283
timestamp 1624047346
transform 1 0 27140 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_286
timestamp 1624047346
transform 1 0 27416 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1624047346
transform -1 0 28704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1624047346
transform 1 0 28704 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _093_
timestamp 1624047346
transform 1 0 29072 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _208_
timestamp 1624047346
transform -1 0 30176 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_309
timestamp 1624047346
transform 1 0 29532 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1624047346
transform 1 0 30176 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1624047346
transform 1 0 30544 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_322
timestamp 1624047346
transform 1 0 30728 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_334
timestamp 1624047346
transform 1 0 31832 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1624047346
transform 1 0 32568 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1624047346
transform 1 0 32660 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_355
timestamp 1624047346
transform 1 0 33764 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_367
timestamp 1624047346
transform 1 0 34868 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1624047346
transform -1 0 36064 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_375
timestamp 1624047346
transform 1 0 35604 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_380
timestamp 1624047346
transform 1 0 36064 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _144_
timestamp 1624047346
transform 1 0 36892 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1624047346
transform 1 0 37812 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_388
timestamp 1624047346
transform 1 0 36800 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_395
timestamp 1624047346
transform 1 0 37444 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_400
timestamp 1624047346
transform 1 0 37904 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _227_
timestamp 1624047346
transform 1 0 38640 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_25_413
timestamp 1624047346
transform 1 0 39100 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _225_
timestamp 1624047346
transform 1 0 40388 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_425
timestamp 1624047346
transform 1 0 40204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_436
timestamp 1624047346
transform 1 0 41216 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_448
timestamp 1624047346
transform 1 0 42320 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _226_
timestamp 1624047346
transform -1 0 43976 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _228_
timestamp 1624047346
transform 1 0 44344 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1624047346
transform 1 0 43056 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_457
timestamp 1624047346
transform 1 0 43148 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_466
timestamp 1624047346
transform 1 0 43976 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_475
timestamp 1624047346
transform 1 0 44804 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_487
timestamp 1624047346
transform 1 0 45908 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_499
timestamp 1624047346
transform 1 0 47012 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1624047346
transform 1 0 48300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_511
timestamp 1624047346
transform 1 0 48116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_514
timestamp 1624047346
transform 1 0 48392 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_526
timestamp 1624047346
transform 1 0 49496 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_538
timestamp 1624047346
transform 1 0 50600 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_550
timestamp 1624047346
transform 1 0 51704 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1624047346
transform 1 0 53544 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_562
timestamp 1624047346
transform 1 0 52808 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_571
timestamp 1624047346
transform 1 0 53636 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_583
timestamp 1624047346
transform 1 0 54740 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_595
timestamp 1624047346
transform 1 0 55844 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_607
timestamp 1624047346
transform 1 0 56948 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_619
timestamp 1624047346
transform 1 0 58052 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624047346
transform -1 0 58880 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624047346
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624047346
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1624047346
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_7
timestamp 1624047346
transform 1 0 1748 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1624047346
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1624047346
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1624047346
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1624047346
transform 1 0 2852 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1624047346
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1624047346
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1624047346
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_42
timestamp 1624047346
transform 1 0 4968 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1624047346
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1624047346
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_54
timestamp 1624047346
transform 1 0 6072 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_66
timestamp 1624047346
transform 1 0 7176 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_51
timestamp 1624047346
transform 1 0 5796 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_58
timestamp 1624047346
transform 1 0 6440 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1624047346
transform 1 0 8004 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_78
timestamp 1624047346
transform 1 0 8280 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_70
timestamp 1624047346
transform 1 0 7544 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_74
timestamp 1624047346
transform 1 0 7912 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_78
timestamp 1624047346
transform 1 0 8280 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _195_
timestamp 1624047346
transform -1 0 10672 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1624047346
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_87
timestamp 1624047346
transform 1 0 9108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_90
timestamp 1624047346
transform 1 0 9384 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1624047346
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A
timestamp 1624047346
transform 1 0 11040 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1624047346
transform 1 0 10672 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_110
timestamp 1624047346
transform 1 0 11224 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_102
timestamp 1624047346
transform 1 0 10488 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_115
timestamp 1624047346
transform 1 0 11684 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_122
timestamp 1624047346
transform 1 0 12328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_134
timestamp 1624047346
transform 1 0 13432 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_127
timestamp 1624047346
transform 1 0 12788 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1624047346
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_142
timestamp 1624047346
transform 1 0 14168 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_144
timestamp 1624047346
transform 1 0 14352 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_139
timestamp 1624047346
transform 1 0 13892 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_151
timestamp 1624047346
transform 1 0 14996 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_156
timestamp 1624047346
transform 1 0 15456 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_168
timestamp 1624047346
transform 1 0 16560 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_163
timestamp 1624047346
transform 1 0 16100 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1624047346
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_180
timestamp 1624047346
transform 1 0 17664 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_172
timestamp 1624047346
transform 1 0 16928 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1624047346
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1624047346
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_192
timestamp 1624047346
transform 1 0 18768 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_201
timestamp 1624047346
transform 1 0 19596 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1624047346
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _186_
timestamp 1624047346
transform 1 0 21068 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A
timestamp 1624047346
transform 1 0 20516 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_209
timestamp 1624047346
transform 1 0 20332 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1624047346
transform 1 0 20700 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1624047346
transform 1 0 20240 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _192_
timestamp 1624047346
transform 1 0 21712 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _197_
timestamp 1624047346
transform 1 0 22632 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1624047346
transform 1 0 22080 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_220
timestamp 1624047346
transform 1 0 21344 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_230
timestamp 1624047346
transform 1 0 22264 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_220
timestamp 1624047346
transform 1 0 21344 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_229
timestamp 1624047346
transform 1 0 22172 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_240
timestamp 1624047346
transform 1 0 23184 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_252
timestamp 1624047346
transform 1 0 24288 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_241
timestamp 1624047346
transform 1 0 23276 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_259
timestamp 1624047346
transform 1 0 24932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1624047346
transform 1 0 24380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_258
timestamp 1624047346
transform 1 0 24840 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_256
timestamp 1624047346
transform 1 0 24656 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1624047346
transform 1 0 24748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1624047346
transform 1 0 24748 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_266
timestamp 1624047346
transform 1 0 25576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_264
timestamp 1624047346
transform 1 0 25392 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _079_
timestamp 1624047346
transform -1 0 25760 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 1624047346
transform 1 0 25300 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_268
timestamp 1624047346
transform 1 0 25760 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  _117_
timestamp 1624047346
transform -1 0 26772 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _214_
timestamp 1624047346
transform -1 0 26864 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1624047346
transform 1 0 27324 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_280
timestamp 1624047346
transform 1 0 26864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_279
timestamp 1624047346
transform 1 0 26772 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_286
timestamp 1624047346
transform 1 0 27416 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1624047346
transform 1 0 28520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_292
timestamp 1624047346
transform 1 0 27968 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_300
timestamp 1624047346
transform 1 0 28704 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_298
timestamp 1624047346
transform 1 0 28520 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _194_
timestamp 1624047346
transform 1 0 29072 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1624047346
transform 1 0 29992 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_309
timestamp 1624047346
transform 1 0 29532 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_313
timestamp 1624047346
transform 1 0 29900 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_315
timestamp 1624047346
transform 1 0 30084 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_310
timestamp 1624047346
transform 1 0 29624 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_327
timestamp 1624047346
transform 1 0 31188 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_322
timestamp 1624047346
transform 1 0 30728 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_334
timestamp 1624047346
transform 1 0 31832 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1624047346
transform 1 0 32568 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_339
timestamp 1624047346
transform 1 0 32292 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_351
timestamp 1624047346
transform 1 0 33396 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_343
timestamp 1624047346
transform 1 0 32660 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_363
timestamp 1624047346
transform 1 0 34500 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_355
timestamp 1624047346
transform 1 0 33764 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1624047346
transform 1 0 34868 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _135_
timestamp 1624047346
transform 1 0 36248 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1624047346
transform 1 0 35236 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_372
timestamp 1624047346
transform 1 0 35328 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_384
timestamp 1624047346
transform 1 0 36432 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_27_379
timestamp 1624047346
transform 1 0 35972 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _219_
timestamp 1624047346
transform 1 0 37076 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _224_
timestamp 1624047346
transform 1 0 37996 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1624047346
transform 1 0 37812 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_390
timestamp 1624047346
transform 1 0 36984 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_397
timestamp 1624047346
transform 1 0 37628 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_388
timestamp 1624047346
transform 1 0 36800 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_396
timestamp 1624047346
transform 1 0 37536 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_400
timestamp 1624047346
transform 1 0 37904 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_405
timestamp 1624047346
transform 1 0 38364 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_417
timestamp 1624047346
transform 1 0 39468 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_412
timestamp 1624047346
transform 1 0 39008 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1624047346
transform 1 0 40480 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_425
timestamp 1624047346
transform 1 0 40204 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_429
timestamp 1624047346
transform 1 0 40572 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_424
timestamp 1624047346
transform 1 0 40112 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_436
timestamp 1624047346
transform 1 0 41216 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_441
timestamp 1624047346
transform 1 0 41676 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_453
timestamp 1624047346
transform 1 0 42780 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_448
timestamp 1624047346
transform 1 0 42320 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1624047346
transform -1 0 44712 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1624047346
transform 1 0 43056 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_465
timestamp 1624047346
transform 1 0 43884 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_457
timestamp 1624047346
transform 1 0 43148 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_469
timestamp 1624047346
transform 1 0 44252 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1624047346
transform 1 0 45724 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1624047346
transform -1 0 45264 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_474
timestamp 1624047346
transform 1 0 44712 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_480
timestamp 1624047346
transform 1 0 45264 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_484
timestamp 1624047346
transform 1 0 45632 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_486
timestamp 1624047346
transform 1 0 45816 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_481
timestamp 1624047346
transform 1 0 45356 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_498
timestamp 1624047346
transform 1 0 46920 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_493
timestamp 1624047346
transform 1 0 46460 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_505
timestamp 1624047346
transform 1 0 47564 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1624047346
transform 1 0 48300 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_510
timestamp 1624047346
transform 1 0 48024 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_514
timestamp 1624047346
transform 1 0 48392 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_522
timestamp 1624047346
transform 1 0 49128 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_534
timestamp 1624047346
transform 1 0 50232 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_526
timestamp 1624047346
transform 1 0 49496 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_538
timestamp 1624047346
transform 1 0 50600 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1624047346
transform 1 0 50968 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_543
timestamp 1624047346
transform 1 0 51060 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_555
timestamp 1624047346
transform 1 0 52164 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_550
timestamp 1624047346
transform 1 0 51704 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1624047346
transform 1 0 53544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_567
timestamp 1624047346
transform 1 0 53268 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_562
timestamp 1624047346
transform 1 0 52808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_571
timestamp 1624047346
transform 1 0 53636 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__S
timestamp 1624047346
transform 1 0 54372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_579
timestamp 1624047346
transform 1 0 54372 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_581
timestamp 1624047346
transform 1 0 54556 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1624047346
transform 1 0 56212 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_591
timestamp 1624047346
transform 1 0 55476 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_600
timestamp 1624047346
transform 1 0 56304 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_593
timestamp 1624047346
transform 1 0 55660 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_605
timestamp 1624047346
transform 1 0 56764 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1624047346
transform -1 0 58236 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output140
timestamp 1624047346
transform 1 0 57868 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1624047346
transform -1 0 57500 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_612
timestamp 1624047346
transform 1 0 57408 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_616
timestamp 1624047346
transform 1 0 57776 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1624047346
transform 1 0 58236 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_613
timestamp 1624047346
transform 1 0 57500 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1624047346
transform 1 0 58236 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624047346
transform -1 0 58880 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624047346
transform -1 0 58880 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624047346
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output181
timestamp 1624047346
transform -1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output181_A
timestamp 1624047346
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_7
timestamp 1624047346
transform 1 0 1748 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_13
timestamp 1624047346
transform 1 0 2300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1624047346
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_25
timestamp 1624047346
transform 1 0 3404 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1624047346
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_42
timestamp 1624047346
transform 1 0 4968 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_54
timestamp 1624047346
transform 1 0 6072 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_66
timestamp 1624047346
transform 1 0 7176 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_78
timestamp 1624047346
transform 1 0 8280 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1624047346
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_87
timestamp 1624047346
transform 1 0 9108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_99
timestamp 1624047346
transform 1 0 10212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_111
timestamp 1624047346
transform 1 0 11316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_123
timestamp 1624047346
transform 1 0 12420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1624047346
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_135
timestamp 1624047346
transform 1 0 13524 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_144
timestamp 1624047346
transform 1 0 14352 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_156
timestamp 1624047346
transform 1 0 15456 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_168
timestamp 1624047346
transform 1 0 16560 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_180
timestamp 1624047346
transform 1 0 17664 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1624047346
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_192
timestamp 1624047346
transform 1 0 18768 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_201
timestamp 1624047346
transform 1 0 19596 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_213
timestamp 1624047346
transform 1 0 20700 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_225
timestamp 1624047346
transform 1 0 21804 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_237
timestamp 1624047346
transform 1 0 22908 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_249
timestamp 1624047346
transform 1 0 24012 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1624047346
transform 1 0 24748 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_258
timestamp 1624047346
transform 1 0 24840 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1624047346
transform 1 0 26220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1624047346
transform -1 0 27324 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_270
timestamp 1624047346
transform 1 0 25944 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_277
timestamp 1624047346
transform 1 0 26588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_285
timestamp 1624047346
transform 1 0 27324 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1624047346
transform 1 0 27692 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_293
timestamp 1624047346
transform 1 0 28060 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1624047346
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_305
timestamp 1624047346
transform 1 0 29164 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_313
timestamp 1624047346
transform 1 0 29900 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1624047346
transform 1 0 30084 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1624047346
transform 1 0 31188 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1624047346
transform 1 0 32292 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1624047346
transform 1 0 33396 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_363
timestamp 1624047346
transform 1 0 34500 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1624047346
transform 1 0 35236 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_372
timestamp 1624047346
transform 1 0 35328 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_384
timestamp 1624047346
transform 1 0 36432 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_396
timestamp 1624047346
transform 1 0 37536 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_408
timestamp 1624047346
transform 1 0 38640 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_420
timestamp 1624047346
transform 1 0 39744 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1624047346
transform 1 0 40480 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_429
timestamp 1624047346
transform 1 0 40572 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_441
timestamp 1624047346
transform 1 0 41676 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_453
timestamp 1624047346
transform 1 0 42780 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_465
timestamp 1624047346
transform 1 0 43884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1624047346
transform 1 0 45724 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_477
timestamp 1624047346
transform 1 0 44988 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_486
timestamp 1624047346
transform 1 0 45816 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_498
timestamp 1624047346
transform 1 0 46920 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_510
timestamp 1624047346
transform 1 0 48024 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_522
timestamp 1624047346
transform 1 0 49128 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_534
timestamp 1624047346
transform 1 0 50232 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1624047346
transform 1 0 50968 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_543
timestamp 1624047346
transform 1 0 51060 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_555
timestamp 1624047346
transform 1 0 52164 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_567
timestamp 1624047346
transform 1 0 53268 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1624047346
transform 1 0 54740 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A0
timestamp 1624047346
transform -1 0 54372 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_575
timestamp 1624047346
transform 1 0 54004 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_579
timestamp 1624047346
transform 1 0 54372 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1624047346
transform 1 0 56212 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_592
timestamp 1624047346
transform 1 0 55568 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_598
timestamp 1624047346
transform 1 0 56120 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_600
timestamp 1624047346
transform 1 0 56304 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1624047346
transform 1 0 57960 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624047346
transform -1 0 57592 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_614
timestamp 1624047346
transform 1 0 57592 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_621
timestamp 1624047346
transform 1 0 58236 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624047346
transform -1 0 58880 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624047346
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1624047346
transform -1 0 1656 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1624047346
transform -1 0 2208 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__S
timestamp 1624047346
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_6
timestamp 1624047346
transform 1 0 1656 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_12
timestamp 1624047346
transform 1 0 2208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_18
timestamp 1624047346
transform 1 0 2760 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_30
timestamp 1624047346
transform 1 0 3864 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_42
timestamp 1624047346
transform 1 0 4968 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1624047346
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_54
timestamp 1624047346
transform 1 0 6072 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_58
timestamp 1624047346
transform 1 0 6440 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_70
timestamp 1624047346
transform 1 0 7544 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1624047346
transform 1 0 8648 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1624047346
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1624047346
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_106
timestamp 1624047346
transform 1 0 10856 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_115
timestamp 1624047346
transform 1 0 11684 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_127
timestamp 1624047346
transform 1 0 12788 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_139
timestamp 1624047346
transform 1 0 13892 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1624047346
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_163
timestamp 1624047346
transform 1 0 16100 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1624047346
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_172
timestamp 1624047346
transform 1 0 16928 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1624047346
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1624047346
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1624047346
transform 1 0 20240 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1624047346
transform 1 0 22080 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_220
timestamp 1624047346
transform 1 0 21344 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_229
timestamp 1624047346
transform 1 0 22172 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_241
timestamp 1624047346
transform 1 0 23276 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_253
timestamp 1624047346
transform 1 0 24380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_265
timestamp 1624047346
transform 1 0 25484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1624047346
transform 1 0 27324 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_277
timestamp 1624047346
transform 1 0 26588 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_286
timestamp 1624047346
transform 1 0 27416 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_298
timestamp 1624047346
transform 1 0 28520 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_310
timestamp 1624047346
transform 1 0 29624 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_322
timestamp 1624047346
transform 1 0 30728 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_334
timestamp 1624047346
transform 1 0 31832 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1624047346
transform 1 0 32568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_343
timestamp 1624047346
transform 1 0 32660 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_355
timestamp 1624047346
transform 1 0 33764 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1624047346
transform 1 0 34868 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1624047346
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1624047346
transform 1 0 37812 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_391
timestamp 1624047346
transform 1 0 37076 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_400
timestamp 1624047346
transform 1 0 37904 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_412
timestamp 1624047346
transform 1 0 39008 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_424
timestamp 1624047346
transform 1 0 40112 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_436
timestamp 1624047346
transform 1 0 41216 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_448
timestamp 1624047346
transform 1 0 42320 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1624047346
transform 1 0 43056 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_457
timestamp 1624047346
transform 1 0 43148 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_469
timestamp 1624047346
transform 1 0 44252 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_481
timestamp 1624047346
transform 1 0 45356 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_493
timestamp 1624047346
transform 1 0 46460 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1624047346
transform 1 0 47564 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1624047346
transform 1 0 48300 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_514
timestamp 1624047346
transform 1 0 48392 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_526
timestamp 1624047346
transform 1 0 49496 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_538
timestamp 1624047346
transform 1 0 50600 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_550
timestamp 1624047346
transform 1 0 51704 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1624047346
transform 1 0 53544 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_562
timestamp 1624047346
transform 1 0 52808 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_571
timestamp 1624047346
transform 1 0 53636 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_583
timestamp 1624047346
transform 1 0 54740 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_595
timestamp 1624047346
transform 1 0 55844 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_607
timestamp 1624047346
transform 1 0 56948 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_619
timestamp 1624047346
transform 1 0 58052 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624047346
transform -1 0 58880 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _266_
timestamp 1624047346
transform 1 0 1932 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624047346
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624047346
transform -1 0 1564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_5
timestamp 1624047346
transform 1 0 1564 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1624047346
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__266__A1
timestamp 1624047346
transform -1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_18
timestamp 1624047346
transform 1 0 2760 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1624047346
transform 1 0 3312 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_28
timestamp 1624047346
transform 1 0 3680 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_30
timestamp 1624047346
transform 1 0 3864 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_42
timestamp 1624047346
transform 1 0 4968 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_54
timestamp 1624047346
transform 1 0 6072 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_66
timestamp 1624047346
transform 1 0 7176 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_78
timestamp 1624047346
transform 1 0 8280 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1624047346
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_87
timestamp 1624047346
transform 1 0 9108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_99
timestamp 1624047346
transform 1 0 10212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_111
timestamp 1624047346
transform 1 0 11316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_123
timestamp 1624047346
transform 1 0 12420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1624047346
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_135
timestamp 1624047346
transform 1 0 13524 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_144
timestamp 1624047346
transform 1 0 14352 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_156
timestamp 1624047346
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_168
timestamp 1624047346
transform 1 0 16560 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1624047346
transform 1 0 17664 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1624047346
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_192
timestamp 1624047346
transform 1 0 18768 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1624047346
transform 1 0 19596 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_213
timestamp 1624047346
transform 1 0 20700 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_225
timestamp 1624047346
transform 1 0 21804 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_237
timestamp 1624047346
transform 1 0 22908 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_249
timestamp 1624047346
transform 1 0 24012 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1624047346
transform 1 0 24748 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_258
timestamp 1624047346
transform 1 0 24840 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _128_
timestamp 1624047346
transform 1 0 27416 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _130_
timestamp 1624047346
transform 1 0 26404 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_270
timestamp 1624047346
transform 1 0 25944 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1624047346
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_278
timestamp 1624047346
transform 1 0 26680 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_295
timestamp 1624047346
transform 1 0 28244 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1624047346
transform 1 0 29992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_307
timestamp 1624047346
transform 1 0 29348 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_313
timestamp 1624047346
transform 1 0 29900 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_315
timestamp 1624047346
transform 1 0 30084 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_327
timestamp 1624047346
transform 1 0 31188 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1624047346
transform 1 0 32292 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1624047346
transform 1 0 33396 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_363
timestamp 1624047346
transform 1 0 34500 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1624047346
transform 1 0 35236 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1624047346
transform 1 0 35328 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1624047346
transform 1 0 36432 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_396
timestamp 1624047346
transform 1 0 37536 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_408
timestamp 1624047346
transform 1 0 38640 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_420
timestamp 1624047346
transform 1 0 39744 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1624047346
transform 1 0 40480 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_429
timestamp 1624047346
transform 1 0 40572 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_441
timestamp 1624047346
transform 1 0 41676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_453
timestamp 1624047346
transform 1 0 42780 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_465
timestamp 1624047346
transform 1 0 43884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1624047346
transform 1 0 45724 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_477
timestamp 1624047346
transform 1 0 44988 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_486
timestamp 1624047346
transform 1 0 45816 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_498
timestamp 1624047346
transform 1 0 46920 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_510
timestamp 1624047346
transform 1 0 48024 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_522
timestamp 1624047346
transform 1 0 49128 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_534
timestamp 1624047346
transform 1 0 50232 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1624047346
transform 1 0 50968 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_543
timestamp 1624047346
transform 1 0 51060 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_555
timestamp 1624047346
transform 1 0 52164 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_567
timestamp 1624047346
transform 1 0 53268 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_579
timestamp 1624047346
transform 1 0 54372 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1624047346
transform 1 0 56212 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_591
timestamp 1624047346
transform 1 0 55476 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_600
timestamp 1624047346
transform 1 0 56304 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_612
timestamp 1624047346
transform 1 0 57408 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624047346
transform -1 0 58880 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_624
timestamp 1624047346
transform 1 0 58512 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1624047346
transform 1 0 2208 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624047346
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1624047346
transform -1 0 1656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_6
timestamp 1624047346
transform 1 0 1656 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1624047346
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1624047346
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1624047346
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1624047346
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_51
timestamp 1624047346
transform 1 0 5796 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_58
timestamp 1624047346
transform 1 0 6440 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1624047346
transform 1 0 8648 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_70
timestamp 1624047346
transform 1 0 7544 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_85
timestamp 1624047346
transform 1 0 8924 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_97
timestamp 1624047346
transform 1 0 10028 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1624047346
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_109
timestamp 1624047346
transform 1 0 11132 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 1624047346
transform 1 0 11500 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_115
timestamp 1624047346
transform 1 0 11684 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_127
timestamp 1624047346
transform 1 0 12788 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_139
timestamp 1624047346
transform 1 0 13892 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_151
timestamp 1624047346
transform 1 0 14996 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1624047346
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_165
timestamp 1624047346
transform 1 0 16284 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1624047346
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_172
timestamp 1624047346
transform 1 0 16928 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1624047346
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1624047346
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1624047346
transform 1 0 20240 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1624047346
transform 1 0 22080 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_220
timestamp 1624047346
transform 1 0 21344 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1624047346
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_241
timestamp 1624047346
transform 1 0 23276 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_253
timestamp 1624047346
transform 1 0 24380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_265
timestamp 1624047346
transform 1 0 25484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1624047346
transform 1 0 27324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_277
timestamp 1624047346
transform 1 0 26588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1624047346
transform 1 0 27416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_298
timestamp 1624047346
transform 1 0 28520 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_310
timestamp 1624047346
transform 1 0 29624 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_322
timestamp 1624047346
transform 1 0 30728 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_334
timestamp 1624047346
transform 1 0 31832 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1624047346
transform 1 0 32568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A
timestamp 1624047346
transform 1 0 32660 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_345
timestamp 1624047346
transform 1 0 32844 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_357
timestamp 1624047346
transform 1 0 33948 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_369
timestamp 1624047346
transform 1 0 35052 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_381
timestamp 1624047346
transform 1 0 36156 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1624047346
transform 1 0 37812 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1624047346
transform 1 0 37260 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_400
timestamp 1624047346
transform 1 0 37904 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_412
timestamp 1624047346
transform 1 0 39008 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_424
timestamp 1624047346
transform 1 0 40112 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_436
timestamp 1624047346
transform 1 0 41216 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_448
timestamp 1624047346
transform 1 0 42320 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1624047346
transform 1 0 43056 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_457
timestamp 1624047346
transform 1 0 43148 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_469
timestamp 1624047346
transform 1 0 44252 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_481
timestamp 1624047346
transform 1 0 45356 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_493
timestamp 1624047346
transform 1 0 46460 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_505
timestamp 1624047346
transform 1 0 47564 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1624047346
transform 1 0 48300 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_514
timestamp 1624047346
transform 1 0 48392 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_526
timestamp 1624047346
transform 1 0 49496 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_538
timestamp 1624047346
transform 1 0 50600 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_550
timestamp 1624047346
transform 1 0 51704 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1624047346
transform 1 0 53544 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_562
timestamp 1624047346
transform 1 0 52808 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_571
timestamp 1624047346
transform 1 0 53636 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_583
timestamp 1624047346
transform 1 0 54740 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_595
timestamp 1624047346
transform 1 0 55844 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1624047346
transform 1 0 57868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output130_A
timestamp 1624047346
transform -1 0 57500 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_607
timestamp 1624047346
transform 1 0 56948 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_613
timestamp 1624047346
transform 1 0 57500 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_621
timestamp 1624047346
transform 1 0 58236 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624047346
transform -1 0 58880 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _211_
timestamp 1624047346
transform 1 0 2300 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624047346
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1624047346
transform 1 0 1380 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_11
timestamp 1624047346
transform 1 0 2116 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_16
timestamp 1624047346
transform 1 0 2576 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _212_
timestamp 1624047346
transform -1 0 3220 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1624047346
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1624047346
transform 1 0 3864 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_23
timestamp 1624047346
transform 1 0 3220 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1624047346
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1624047346
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1624047346
transform 1 0 6256 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1624047346
transform 1 0 7360 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_80
timestamp 1624047346
transform 1 0 8464 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1624047346
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_87
timestamp 1624047346
transform 1 0 9108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_99
timestamp 1624047346
transform 1 0 10212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_111
timestamp 1624047346
transform 1 0 11316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_123
timestamp 1624047346
transform 1 0 12420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1624047346
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_135
timestamp 1624047346
transform 1 0 13524 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_144
timestamp 1624047346
transform 1 0 14352 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_8  _121_
timestamp 1624047346
transform -1 0 18032 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_1  _123_
timestamp 1624047346
transform 1 0 15824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_156
timestamp 1624047346
transform 1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_163
timestamp 1624047346
transform 1 0 16100 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_167
timestamp 1624047346
transform 1 0 16468 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_184
timestamp 1624047346
transform 1 0 18032 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1624047346
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1624047346
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_190
timestamp 1624047346
transform 1 0 18584 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_198
timestamp 1624047346
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1624047346
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_213
timestamp 1624047346
transform 1 0 20700 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp 1624047346
transform 1 0 21804 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1624047346
transform -1 0 22632 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1624047346
transform 1 0 22080 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_234
timestamp 1624047346
transform 1 0 22632 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_246
timestamp 1624047346
transform 1 0 23736 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1624047346
transform 1 0 24748 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_254
timestamp 1624047346
transform 1 0 24472 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_258
timestamp 1624047346
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_270
timestamp 1624047346
transform 1 0 25944 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_282
timestamp 1624047346
transform 1 0 27048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_294
timestamp 1624047346
transform 1 0 28152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1624047346
transform 1 0 29992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_306
timestamp 1624047346
transform 1 0 29256 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_315
timestamp 1624047346
transform 1 0 30084 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1624047346
transform -1 0 32200 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _232_
timestamp 1624047346
transform 1 0 31096 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_32_323
timestamp 1624047346
transform 1 0 30820 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_331
timestamp 1624047346
transform 1 0 31556 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _161_
timestamp 1624047346
transform 1 0 32568 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1624047346
transform 1 0 32200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_345
timestamp 1624047346
transform 1 0 32844 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_357
timestamp 1624047346
transform 1 0 33948 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_369
timestamp 1624047346
transform 1 0 35052 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _175_
timestamp 1624047346
transform 1 0 36340 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1624047346
transform 1 0 35236 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__A
timestamp 1624047346
transform 1 0 35788 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_372
timestamp 1624047346
transform 1 0 35328 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_376
timestamp 1624047346
transform 1 0 35696 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_379
timestamp 1624047346
transform 1 0 35972 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_386
timestamp 1624047346
transform 1 0 36616 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _242_
timestamp 1624047346
transform 1 0 36984 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_32_395
timestamp 1624047346
transform 1 0 37444 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_407
timestamp 1624047346
transform 1 0 38548 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_419
timestamp 1624047346
transform 1 0 39652 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1624047346
transform 1 0 40480 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_427
timestamp 1624047346
transform 1 0 40388 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_429
timestamp 1624047346
transform 1 0 40572 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_441
timestamp 1624047346
transform 1 0 41676 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_453
timestamp 1624047346
transform 1 0 42780 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_465
timestamp 1624047346
transform 1 0 43884 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1624047346
transform 1 0 45724 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_477
timestamp 1624047346
transform 1 0 44988 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_486
timestamp 1624047346
transform 1 0 45816 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_498
timestamp 1624047346
transform 1 0 46920 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_510
timestamp 1624047346
transform 1 0 48024 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_522
timestamp 1624047346
transform 1 0 49128 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_534
timestamp 1624047346
transform 1 0 50232 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1624047346
transform 1 0 50968 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_543
timestamp 1624047346
transform 1 0 51060 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_555
timestamp 1624047346
transform 1 0 52164 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_567
timestamp 1624047346
transform 1 0 53268 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_579
timestamp 1624047346
transform 1 0 54372 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1624047346
transform 1 0 56212 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_591
timestamp 1624047346
transform 1 0 55476 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_600
timestamp 1624047346
transform 1 0 56304 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output151
timestamp 1624047346
transform 1 0 57868 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output151_A
timestamp 1624047346
transform -1 0 57500 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_608
timestamp 1624047346
transform 1 0 57040 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1624047346
transform 1 0 57500 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1624047346
transform 1 0 58236 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624047346
transform -1 0 58880 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624047346
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1624047346
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1624047346
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output157
timestamp 1624047346
transform -1 0 1748 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624047346
transform -1 0 2208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1624047346
transform -1 0 2760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_6
timestamp 1624047346
transform 1 0 1656 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_12
timestamp 1624047346
transform 1 0 2208 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_7
timestamp 1624047346
transform 1 0 1748 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1624047346
transform 1 0 3772 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_18
timestamp 1624047346
transform 1 0 2760 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_30
timestamp 1624047346
transform 1 0 3864 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_19
timestamp 1624047346
transform 1 0 2852 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_27
timestamp 1624047346
transform 1 0 3588 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_30
timestamp 1624047346
transform 1 0 3864 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_42
timestamp 1624047346
transform 1 0 4968 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_42
timestamp 1624047346
transform 1 0 4968 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1624047346
transform 1 0 6348 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_54
timestamp 1624047346
transform 1 0 6072 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_58
timestamp 1624047346
transform 1 0 6440 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_54
timestamp 1624047346
transform 1 0 6072 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1624047346
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_70
timestamp 1624047346
transform 1 0 7544 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_82
timestamp 1624047346
transform 1 0 8648 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_78
timestamp 1624047346
transform 1 0 8280 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1624047346
transform 1 0 9016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1624047346
transform 1 0 9752 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_87
timestamp 1624047346
transform 1 0 9108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_99
timestamp 1624047346
transform 1 0 10212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1624047346
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_106
timestamp 1624047346
transform 1 0 10856 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_115
timestamp 1624047346
transform 1 0 11684 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_111
timestamp 1624047346
transform 1 0 11316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_127
timestamp 1624047346
transform 1 0 12788 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_123
timestamp 1624047346
transform 1 0 12420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1624047346
transform 1 0 14260 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_139
timestamp 1624047346
transform 1 0 13892 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_151
timestamp 1624047346
transform 1 0 14996 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_135
timestamp 1624047346
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_144
timestamp 1624047346
transform 1 0 14352 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_163
timestamp 1624047346
transform 1 0 16100 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_156
timestamp 1624047346
transform 1 0 15456 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1624047346
transform 1 0 16560 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1624047346
transform 1 0 16836 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_172
timestamp 1624047346
transform 1 0 16928 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1624047346
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_180
timestamp 1624047346
transform 1 0 17664 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1624047346
transform 1 0 19504 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1624047346
transform 1 0 19136 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_192
timestamp 1624047346
transform 1 0 18768 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1624047346
transform 1 0 19596 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1624047346
transform -1 0 20240 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A
timestamp 1624047346
transform -1 0 20792 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1624047346
transform 1 0 20240 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_208
timestamp 1624047346
transform 1 0 20240 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_214
timestamp 1624047346
transform 1 0 20792 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _238_
timestamp 1624047346
transform -1 0 23460 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1624047346
transform 1 0 22080 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1624047346
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1624047346
transform 1 0 22172 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_233
timestamp 1624047346
transform 1 0 22540 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_226
timestamp 1624047346
transform 1 0 21896 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_243
timestamp 1624047346
transform 1 0 23460 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_238
timestamp 1624047346
transform 1 0 23000 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_250
timestamp 1624047346
transform 1 0 24104 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1624047346
transform 1 0 24748 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_255
timestamp 1624047346
transform 1 0 24564 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_267
timestamp 1624047346
transform 1 0 25668 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_256
timestamp 1624047346
transform 1 0 24656 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1624047346
transform 1 0 24840 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1624047346
transform 1 0 27324 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_279
timestamp 1624047346
transform 1 0 26772 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_286
timestamp 1624047346
transform 1 0 27416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_270
timestamp 1624047346
transform 1 0 25944 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_282
timestamp 1624047346
transform 1 0 27048 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _233_
timestamp 1624047346
transform -1 0 28520 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _235_
timestamp 1624047346
transform -1 0 29440 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_298
timestamp 1624047346
transform 1 0 28520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_288
timestamp 1624047346
transform 1 0 27600 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_298
timestamp 1624047346
transform 1 0 28520 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1624047346
transform 1 0 29992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_310
timestamp 1624047346
transform 1 0 29624 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_308
timestamp 1624047346
transform 1 0 29440 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_315
timestamp 1624047346
transform 1 0 30084 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_319
timestamp 1624047346
transform 1 0 30452 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _162_
timestamp 1624047346
transform 1 0 31372 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _230_
timestamp 1624047346
transform -1 0 31096 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _234_
timestamp 1624047346
transform 1 0 31648 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_33_322
timestamp 1624047346
transform 1 0 30728 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_328
timestamp 1624047346
transform 1 0 31280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_334
timestamp 1624047346
transform 1 0 31832 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_326
timestamp 1624047346
transform 1 0 31096 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1624047346
transform 1 0 32568 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_343
timestamp 1624047346
transform 1 0 32660 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_341
timestamp 1624047346
transform 1 0 32476 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_353
timestamp 1624047346
transform 1 0 33580 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_355
timestamp 1624047346
transform 1 0 33764 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1624047346
transform 1 0 34868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_365
timestamp 1624047346
transform 1 0 34684 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _180_
timestamp 1624047346
transform -1 0 36616 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _241_
timestamp 1624047346
transform 1 0 36248 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1624047346
transform 1 0 35236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_379
timestamp 1624047346
transform 1 0 35972 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_372
timestamp 1624047346
transform 1 0 35328 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_376
timestamp 1624047346
transform 1 0 35696 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_386
timestamp 1624047346
transform 1 0 36616 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _174_
timestamp 1624047346
transform -1 0 37444 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _176_
timestamp 1624047346
transform 1 0 37812 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1624047346
transform -1 0 38548 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1624047346
transform 1 0 37812 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_391
timestamp 1624047346
transform 1 0 37076 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_400
timestamp 1624047346
transform 1 0 37904 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_395
timestamp 1624047346
transform 1 0 37444 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_404
timestamp 1624047346
transform 1 0 38272 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _173_
timestamp 1624047346
transform -1 0 38916 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__A
timestamp 1624047346
transform -1 0 39100 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_407
timestamp 1624047346
transform 1 0 38548 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_413
timestamp 1624047346
transform 1 0 39100 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_411
timestamp 1624047346
transform 1 0 38916 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1624047346
transform 1 0 40480 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_425
timestamp 1624047346
transform 1 0 40204 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_437
timestamp 1624047346
transform 1 0 41308 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_423
timestamp 1624047346
transform 1 0 40020 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_427
timestamp 1624047346
transform 1 0 40388 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_429
timestamp 1624047346
transform 1 0 40572 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_449
timestamp 1624047346
transform 1 0 42412 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_441
timestamp 1624047346
transform 1 0 41676 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_453
timestamp 1624047346
transform 1 0 42780 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1624047346
transform 1 0 43056 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_455
timestamp 1624047346
transform 1 0 42964 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_457
timestamp 1624047346
transform 1 0 43148 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_469
timestamp 1624047346
transform 1 0 44252 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_465
timestamp 1624047346
transform 1 0 43884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1624047346
transform 1 0 45724 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_481
timestamp 1624047346
transform 1 0 45356 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_477
timestamp 1624047346
transform 1 0 44988 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_486
timestamp 1624047346
transform 1 0 45816 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A0
timestamp 1624047346
transform 1 0 47196 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__S
timestamp 1624047346
transform 1 0 47380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_493
timestamp 1624047346
transform 1 0 46460 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_501
timestamp 1624047346
transform 1 0 47196 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1624047346
transform 1 0 47564 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_498
timestamp 1624047346
transform 1 0 46920 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_503
timestamp 1624047346
transform 1 0 47380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1624047346
transform 1 0 47748 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1624047346
transform 1 0 48300 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_514
timestamp 1624047346
transform 1 0 48392 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_516
timestamp 1624047346
transform 1 0 48576 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_526
timestamp 1624047346
transform 1 0 49496 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_538
timestamp 1624047346
transform 1 0 50600 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_528
timestamp 1624047346
transform 1 0 49680 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1624047346
transform 1 0 50968 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_550
timestamp 1624047346
transform 1 0 51704 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_540
timestamp 1624047346
transform 1 0 50784 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_543
timestamp 1624047346
transform 1 0 51060 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_555
timestamp 1624047346
transform 1 0 52164 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1624047346
transform 1 0 53544 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_562
timestamp 1624047346
transform 1 0 52808 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_571
timestamp 1624047346
transform 1 0 53636 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_567
timestamp 1624047346
transform 1 0 53268 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_583
timestamp 1624047346
transform 1 0 54740 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_579
timestamp 1624047346
transform 1 0 54372 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1624047346
transform 1 0 56212 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_595
timestamp 1624047346
transform 1 0 55844 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_591
timestamp 1624047346
transform 1 0 55476 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_600
timestamp 1624047346
transform 1 0 56304 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1624047346
transform 1 0 57960 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1624047346
transform -1 0 57592 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_607
timestamp 1624047346
transform 1 0 56948 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_619
timestamp 1624047346
transform 1 0 58052 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_614
timestamp 1624047346
transform 1 0 57592 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_621
timestamp 1624047346
transform 1 0 58236 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624047346
transform -1 0 58880 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1624047346
transform -1 0 58880 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1624047346
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1624047346
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1624047346
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1624047346
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1624047346
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1624047346
transform 1 0 6348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_51
timestamp 1624047346
transform 1 0 5796 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_58
timestamp 1624047346
transform 1 0 6440 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_70
timestamp 1624047346
transform 1 0 7544 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1624047346
transform 1 0 8648 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1624047346
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1624047346
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_106
timestamp 1624047346
transform 1 0 10856 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1624047346
transform 1 0 11684 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_127
timestamp 1624047346
transform 1 0 12788 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_139
timestamp 1624047346
transform 1 0 13892 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_151
timestamp 1624047346
transform 1 0 14996 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_163
timestamp 1624047346
transform 1 0 16100 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1624047346
transform 1 0 16836 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_172
timestamp 1624047346
transform 1 0 16928 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1624047346
transform 1 0 18032 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_196
timestamp 1624047346
transform 1 0 19136 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_202
timestamp 1624047346
transform 1 0 19688 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _156_
timestamp 1624047346
transform 1 0 20424 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _231_
timestamp 1624047346
transform 1 0 19780 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_206
timestamp 1624047346
transform 1 0 20056 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_213
timestamp 1624047346
transform 1 0 20700 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1624047346
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1624047346
transform 1 0 21804 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_229
timestamp 1624047346
transform 1 0 22172 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_241
timestamp 1624047346
transform 1 0 23276 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_253
timestamp 1624047346
transform 1 0 24380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_265
timestamp 1624047346
transform 1 0 25484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1624047346
transform 1 0 27324 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_277
timestamp 1624047346
transform 1 0 26588 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_286
timestamp 1624047346
transform 1 0 27416 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _229_
timestamp 1624047346
transform 1 0 28704 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_298
timestamp 1624047346
transform 1 0 28520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_303
timestamp 1624047346
transform 1 0 28980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1624047346
transform 1 0 30452 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1624047346
transform 1 0 29348 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_309
timestamp 1624047346
transform 1 0 29532 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_317
timestamp 1624047346
transform 1 0 30268 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _158_
timestamp 1624047346
transform -1 0 31464 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_323
timestamp 1624047346
transform 1 0 30820 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_330
timestamp 1624047346
transform 1 0 31464 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1624047346
transform 1 0 32568 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_343
timestamp 1624047346
transform 1 0 32660 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_355
timestamp 1624047346
transform 1 0 33764 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_367
timestamp 1624047346
transform 1 0 34868 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _172_
timestamp 1624047346
transform 1 0 35880 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _243_
timestamp 1624047346
transform -1 0 37076 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_35_375
timestamp 1624047346
transform 1 0 35604 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_382
timestamp 1624047346
transform 1 0 36248 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _178_
timestamp 1624047346
transform 1 0 38272 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1624047346
transform 1 0 37812 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_391
timestamp 1624047346
transform 1 0 37076 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_400
timestamp 1624047346
transform 1 0 37904 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_413
timestamp 1624047346
transform 1 0 39100 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_425
timestamp 1624047346
transform 1 0 40204 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_437
timestamp 1624047346
transform 1 0 41308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_449
timestamp 1624047346
transform 1 0 42412 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1624047346
transform 1 0 43056 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_455
timestamp 1624047346
transform 1 0 42964 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_457
timestamp 1624047346
transform 1 0 43148 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_469
timestamp 1624047346
transform 1 0 44252 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_481
timestamp 1624047346
transform 1 0 45356 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_493
timestamp 1624047346
transform 1 0 46460 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_505
timestamp 1624047346
transform 1 0 47564 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1624047346
transform 1 0 48300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_514
timestamp 1624047346
transform 1 0 48392 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_526
timestamp 1624047346
transform 1 0 49496 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_538
timestamp 1624047346
transform 1 0 50600 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_550
timestamp 1624047346
transform 1 0 51704 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1624047346
transform 1 0 53544 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_562
timestamp 1624047346
transform 1 0 52808 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_571
timestamp 1624047346
transform 1 0 53636 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_583
timestamp 1624047346
transform 1 0 54740 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_595
timestamp 1624047346
transform 1 0 55844 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_607
timestamp 1624047346
transform 1 0 56948 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_619
timestamp 1624047346
transform 1 0 58052 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1624047346
transform -1 0 58880 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1624047346
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1624047346
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1624047346
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1624047346
transform 1 0 3772 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_27
timestamp 1624047346
transform 1 0 3588 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_30
timestamp 1624047346
transform 1 0 3864 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_42
timestamp 1624047346
transform 1 0 4968 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_54
timestamp 1624047346
transform 1 0 6072 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_66
timestamp 1624047346
transform 1 0 7176 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_78
timestamp 1624047346
transform 1 0 8280 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1624047346
transform 1 0 9016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_87
timestamp 1624047346
transform 1 0 9108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_99
timestamp 1624047346
transform 1 0 10212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_111
timestamp 1624047346
transform 1 0 11316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_123
timestamp 1624047346
transform 1 0 12420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1624047346
transform 1 0 14260 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_135
timestamp 1624047346
transform 1 0 13524 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_144
timestamp 1624047346
transform 1 0 14352 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_156
timestamp 1624047346
transform 1 0 15456 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_168
timestamp 1624047346
transform 1 0 16560 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_180
timestamp 1624047346
transform 1 0 17664 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1624047346
transform 1 0 19504 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_192
timestamp 1624047346
transform 1 0 18768 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1624047346
transform 1 0 19596 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_213
timestamp 1624047346
transform 1 0 20700 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1624047346
transform 1 0 21804 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_237
timestamp 1624047346
transform 1 0 22908 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_249
timestamp 1624047346
transform 1 0 24012 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1624047346
transform 1 0 24748 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1624047346
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _160_
timestamp 1624047346
transform -1 0 27508 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_270
timestamp 1624047346
transform 1 0 25944 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_282
timestamp 1624047346
transform 1 0 27048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_287
timestamp 1624047346
transform 1 0 27508 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_299
timestamp 1624047346
transform 1 0 28612 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1624047346
transform 1 0 29992 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_311
timestamp 1624047346
transform 1 0 29716 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_315
timestamp 1624047346
transform 1 0 30084 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_327
timestamp 1624047346
transform 1 0 31188 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_339
timestamp 1624047346
transform 1 0 32292 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_351
timestamp 1624047346
transform 1 0 33396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_363
timestamp 1624047346
transform 1 0 34500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _240_
timestamp 1624047346
transform 1 0 36156 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1624047346
transform 1 0 35236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_372
timestamp 1624047346
transform 1 0 35328 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_380
timestamp 1624047346
transform 1 0 36064 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_385
timestamp 1624047346
transform 1 0 36524 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _245_
timestamp 1624047346
transform 1 0 36892 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_393
timestamp 1624047346
transform 1 0 37260 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_405
timestamp 1624047346
transform 1 0 38364 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_417
timestamp 1624047346
transform 1 0 39468 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1624047346
transform 1 0 40480 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_425
timestamp 1624047346
transform 1 0 40204 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_429
timestamp 1624047346
transform 1 0 40572 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_441
timestamp 1624047346
transform 1 0 41676 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_453
timestamp 1624047346
transform 1 0 42780 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_465
timestamp 1624047346
transform 1 0 43884 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1624047346
transform 1 0 45724 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_477
timestamp 1624047346
transform 1 0 44988 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_486
timestamp 1624047346
transform 1 0 45816 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_498
timestamp 1624047346
transform 1 0 46920 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_510
timestamp 1624047346
transform 1 0 48024 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_522
timestamp 1624047346
transform 1 0 49128 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_534
timestamp 1624047346
transform 1 0 50232 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1624047346
transform 1 0 50968 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_543
timestamp 1624047346
transform 1 0 51060 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_555
timestamp 1624047346
transform 1 0 52164 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_567
timestamp 1624047346
transform 1 0 53268 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_579
timestamp 1624047346
transform 1 0 54372 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1624047346
transform 1 0 56212 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_591
timestamp 1624047346
transform 1 0 55476 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_600
timestamp 1624047346
transform 1 0 56304 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output199
timestamp 1624047346
transform 1 0 57868 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output199_A
timestamp 1624047346
transform 1 0 57316 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_608
timestamp 1624047346
transform 1 0 57040 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_613
timestamp 1624047346
transform 1 0 57500 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_621
timestamp 1624047346
transform 1 0 58236 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1624047346
transform -1 0 58880 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1624047346
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output197
timestamp 1624047346
transform -1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output197_A
timestamp 1624047346
transform -1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_7
timestamp 1624047346
transform 1 0 1748 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_13
timestamp 1624047346
transform 1 0 2300 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater247_A
timestamp 1624047346
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_25
timestamp 1624047346
transform 1 0 3404 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_31
timestamp 1624047346
transform 1 0 3956 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_34
timestamp 1624047346
transform 1 0 4232 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_46
timestamp 1624047346
transform 1 0 5336 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1624047346
transform 1 0 6348 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_54
timestamp 1624047346
transform 1 0 6072 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_58
timestamp 1624047346
transform 1 0 6440 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_70
timestamp 1624047346
transform 1 0 7544 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_82
timestamp 1624047346
transform 1 0 8648 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_94
timestamp 1624047346
transform 1 0 9752 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1624047346
transform 1 0 11592 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_106
timestamp 1624047346
transform 1 0 10856 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_115
timestamp 1624047346
transform 1 0 11684 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_127
timestamp 1624047346
transform 1 0 12788 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1624047346
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1624047346
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_163
timestamp 1624047346
transform 1 0 16100 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1624047346
transform 1 0 16836 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_172
timestamp 1624047346
transform 1 0 16928 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1624047346
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1624047346
transform 1 0 19136 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_2  _171_
timestamp 1624047346
transform -1 0 21528 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_37_208
timestamp 1624047346
transform 1 0 20240 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_216
timestamp 1624047346
transform 1 0 20976 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1624047346
transform 1 0 22080 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_222
timestamp 1624047346
transform 1 0 21528 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_229
timestamp 1624047346
transform 1 0 22172 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_241
timestamp 1624047346
transform 1 0 23276 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_253
timestamp 1624047346
transform 1 0 24380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_265
timestamp 1624047346
transform 1 0 25484 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _159_
timestamp 1624047346
transform 1 0 26404 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1624047346
transform 1 0 27324 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_273
timestamp 1624047346
transform 1 0 26220 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_278
timestamp 1624047346
transform 1 0 26680 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_284
timestamp 1624047346
transform 1 0 27232 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_286
timestamp 1624047346
transform 1 0 27416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1624047346
transform 1 0 28520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_310
timestamp 1624047346
transform 1 0 29624 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_322
timestamp 1624047346
transform 1 0 30728 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_334
timestamp 1624047346
transform 1 0 31832 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1624047346
transform 1 0 32568 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_343
timestamp 1624047346
transform 1 0 32660 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__179__A
timestamp 1624047346
transform 1 0 34868 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_355
timestamp 1624047346
transform 1 0 33764 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_369
timestamp 1624047346
transform 1 0 35052 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp 1624047346
transform 1 0 35420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _244_
timestamp 1624047346
transform 1 0 36432 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_376
timestamp 1624047346
transform 1 0 35696 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_387
timestamp 1624047346
transform 1 0 36708 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1624047346
transform 1 0 37812 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_400
timestamp 1624047346
transform 1 0 37904 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_412
timestamp 1624047346
transform 1 0 39008 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_424
timestamp 1624047346
transform 1 0 40112 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_436
timestamp 1624047346
transform 1 0 41216 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_448
timestamp 1624047346
transform 1 0 42320 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1624047346
transform 1 0 43056 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_457
timestamp 1624047346
transform 1 0 43148 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_469
timestamp 1624047346
transform 1 0 44252 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_481
timestamp 1624047346
transform 1 0 45356 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_493
timestamp 1624047346
transform 1 0 46460 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_505
timestamp 1624047346
transform 1 0 47564 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1624047346
transform 1 0 48300 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_514
timestamp 1624047346
transform 1 0 48392 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_526
timestamp 1624047346
transform 1 0 49496 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_538
timestamp 1624047346
transform 1 0 50600 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_550
timestamp 1624047346
transform 1 0 51704 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1624047346
transform 1 0 53544 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_562
timestamp 1624047346
transform 1 0 52808 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_571
timestamp 1624047346
transform 1 0 53636 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_583
timestamp 1624047346
transform 1 0 54740 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_595
timestamp 1624047346
transform 1 0 55844 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624047346
transform -1 0 58236 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624047346
transform -1 0 57592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_607
timestamp 1624047346
transform 1 0 56948 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_611
timestamp 1624047346
transform 1 0 57316 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_614
timestamp 1624047346
transform 1 0 57592 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_621
timestamp 1624047346
transform 1 0 58236 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1624047346
transform -1 0 58880 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1624047346
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output240
timestamp 1624047346
transform -1 0 1748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output240_A
timestamp 1624047346
transform 1 0 2116 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_7
timestamp 1624047346
transform 1 0 1748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_13
timestamp 1624047346
transform 1 0 2300 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1624047346
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_25
timestamp 1624047346
transform 1 0 3404 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_30
timestamp 1624047346
transform 1 0 3864 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  repeater247 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform -1 0 5336 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_46
timestamp 1624047346
transform 1 0 5336 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_58
timestamp 1624047346
transform 1 0 6440 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_70
timestamp 1624047346
transform 1 0 7544 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_82
timestamp 1624047346
transform 1 0 8648 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1624047346
transform 1 0 9016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_87
timestamp 1624047346
transform 1 0 9108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_99
timestamp 1624047346
transform 1 0 10212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_111
timestamp 1624047346
transform 1 0 11316 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_123
timestamp 1624047346
transform 1 0 12420 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1624047346
transform 1 0 14260 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_135
timestamp 1624047346
transform 1 0 13524 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_144
timestamp 1624047346
transform 1 0 14352 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_156
timestamp 1624047346
transform 1 0 15456 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1624047346
transform 1 0 16560 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1624047346
transform 1 0 17664 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1624047346
transform 1 0 19504 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_192
timestamp 1624047346
transform 1 0 18768 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_201
timestamp 1624047346
transform 1 0 19596 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _170_
timestamp 1624047346
transform 1 0 20608 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A
timestamp 1624047346
transform -1 0 20240 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_205
timestamp 1624047346
transform 1 0 19964 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_208
timestamp 1624047346
transform 1 0 20240 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_215
timestamp 1624047346
transform 1 0 20884 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _239_
timestamp 1624047346
transform -1 0 21896 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__decap_12  FILLER_38_226
timestamp 1624047346
transform 1 0 21896 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_238
timestamp 1624047346
transform 1 0 23000 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_250
timestamp 1624047346
transform 1 0 24104 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1624047346
transform 1 0 24748 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_256
timestamp 1624047346
transform 1 0 24656 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_258
timestamp 1624047346
transform 1 0 24840 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1624047346
transform -1 0 27784 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_270
timestamp 1624047346
transform 1 0 25944 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_282
timestamp 1624047346
transform 1 0 27048 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_290
timestamp 1624047346
transform 1 0 27784 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_302
timestamp 1624047346
transform 1 0 28888 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1624047346
transform 1 0 29992 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_315
timestamp 1624047346
transform 1 0 30084 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_327
timestamp 1624047346
transform 1 0 31188 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_339
timestamp 1624047346
transform 1 0 32292 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_351
timestamp 1624047346
transform 1 0 33396 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_363
timestamp 1624047346
transform 1 0 34500 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1624047346
transform 1 0 35236 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_372
timestamp 1624047346
transform 1 0 35328 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_384
timestamp 1624047346
transform 1 0 36432 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_396
timestamp 1624047346
transform 1 0 37536 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_408
timestamp 1624047346
transform 1 0 38640 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_420
timestamp 1624047346
transform 1 0 39744 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1624047346
transform 1 0 40480 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_429
timestamp 1624047346
transform 1 0 40572 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_441
timestamp 1624047346
transform 1 0 41676 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_453
timestamp 1624047346
transform 1 0 42780 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_465
timestamp 1624047346
transform 1 0 43884 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1624047346
transform 1 0 45724 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1624047346
transform 1 0 44988 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_486
timestamp 1624047346
transform 1 0 45816 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_498
timestamp 1624047346
transform 1 0 46920 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_510
timestamp 1624047346
transform 1 0 48024 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_522
timestamp 1624047346
transform 1 0 49128 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_534
timestamp 1624047346
transform 1 0 50232 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1624047346
transform 1 0 50968 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_543
timestamp 1624047346
transform 1 0 51060 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_555
timestamp 1624047346
transform 1 0 52164 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_567
timestamp 1624047346
transform 1 0 53268 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_579
timestamp 1624047346
transform 1 0 54372 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1624047346
transform 1 0 56212 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_591
timestamp 1624047346
transform 1 0 55476 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_600
timestamp 1624047346
transform 1 0 56304 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_612
timestamp 1624047346
transform 1 0 57408 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1624047346
transform -1 0 58880 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_624
timestamp 1624047346
transform 1 0 58512 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1624047346
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1624047346
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1624047346
transform -1 0 1748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1624047346
transform -1 0 2300 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1624047346
transform 1 0 1748 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_13
timestamp 1624047346
transform 1 0 2300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1624047346
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1624047346
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1624047346
transform 1 0 3772 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_25
timestamp 1624047346
transform 1 0 3404 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1624047346
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_30
timestamp 1624047346
transform 1 0 3864 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_37
timestamp 1624047346
transform 1 0 4508 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_49
timestamp 1624047346
transform 1 0 5612 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_42
timestamp 1624047346
transform 1 0 4968 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1624047346
transform 1 0 6348 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_58
timestamp 1624047346
transform 1 0 6440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_54
timestamp 1624047346
transform 1 0 6072 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_66
timestamp 1624047346
transform 1 0 7176 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_70
timestamp 1624047346
transform 1 0 7544 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_82
timestamp 1624047346
transform 1 0 8648 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_78
timestamp 1624047346
transform 1 0 8280 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1624047346
transform 1 0 9016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_94
timestamp 1624047346
transform 1 0 9752 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_87
timestamp 1624047346
transform 1 0 9108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_99
timestamp 1624047346
transform 1 0 10212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1624047346
transform 1 0 11592 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_106
timestamp 1624047346
transform 1 0 10856 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_115
timestamp 1624047346
transform 1 0 11684 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_111
timestamp 1624047346
transform 1 0 11316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_127
timestamp 1624047346
transform 1 0 12788 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_123
timestamp 1624047346
transform 1 0 12420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1624047346
transform 1 0 14260 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_139
timestamp 1624047346
transform 1 0 13892 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_151
timestamp 1624047346
transform 1 0 14996 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_135
timestamp 1624047346
transform 1 0 13524 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_144
timestamp 1624047346
transform 1 0 14352 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_163
timestamp 1624047346
transform 1 0 16100 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_156
timestamp 1624047346
transform 1 0 15456 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_168
timestamp 1624047346
transform 1 0 16560 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1624047346
transform 1 0 16836 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_172
timestamp 1624047346
transform 1 0 16928 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1624047346
transform 1 0 18032 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_180
timestamp 1624047346
transform 1 0 17664 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1624047346
transform 1 0 19504 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1624047346
transform 1 0 19136 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_192
timestamp 1624047346
transform 1 0 18768 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1624047346
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1624047346
transform 1 0 20240 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_213
timestamp 1624047346
transform 1 0 20700 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _169_
timestamp 1624047346
transform 1 0 22540 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _236_
timestamp 1624047346
transform -1 0 22908 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1624047346
transform 1 0 22080 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_220
timestamp 1624047346
transform 1 0 21344 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_229
timestamp 1624047346
transform 1 0 22172 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_225
timestamp 1624047346
transform 1 0 21804 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_231
timestamp 1624047346
transform 1 0 22356 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_236
timestamp 1624047346
transform 1 0 22816 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_248
timestamp 1624047346
transform 1 0 23920 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_237
timestamp 1624047346
transform 1 0 22908 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_249
timestamp 1624047346
transform 1 0 24012 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _165_
timestamp 1624047346
transform 1 0 25760 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1624047346
transform 1 0 24748 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_260
timestamp 1624047346
transform 1 0 25024 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1624047346
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1624047346
transform 1 0 27324 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_273
timestamp 1624047346
transform 1 0 26220 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1624047346
transform 1 0 27416 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_270
timestamp 1624047346
transform 1 0 25944 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_282
timestamp 1624047346
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _167_
timestamp 1624047346
transform -1 0 28428 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _237_
timestamp 1624047346
transform -1 0 28612 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_39_299
timestamp 1624047346
transform 1 0 28612 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_297
timestamp 1624047346
transform 1 0 28428 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1624047346
transform 1 0 29992 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_311
timestamp 1624047346
transform 1 0 29716 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_309
timestamp 1624047346
transform 1 0 29532 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_313
timestamp 1624047346
transform 1 0 29900 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_315
timestamp 1624047346
transform 1 0 30084 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_323
timestamp 1624047346
transform 1 0 30820 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_335
timestamp 1624047346
transform 1 0 31924 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_327
timestamp 1624047346
transform 1 0 31188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1624047346
transform 1 0 32568 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1624047346
transform 1 0 32476 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_343
timestamp 1624047346
transform 1 0 32660 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_339
timestamp 1624047346
transform 1 0 32292 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_351
timestamp 1624047346
transform 1 0 33396 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_355
timestamp 1624047346
transform 1 0 33764 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1624047346
transform 1 0 34868 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_363
timestamp 1624047346
transform 1 0 34500 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1624047346
transform 1 0 36708 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1624047346
transform 1 0 35236 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_379
timestamp 1624047346
transform 1 0 35972 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_372
timestamp 1624047346
transform 1 0 35328 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_384
timestamp 1624047346
transform 1 0 36432 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _185_
timestamp 1624047346
transform 1 0 37720 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1624047346
transform 1 0 37812 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_391
timestamp 1624047346
transform 1 0 37076 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_400
timestamp 1624047346
transform 1 0 37904 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_396
timestamp 1624047346
transform 1 0 37536 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 1624047346
transform -1 0 39192 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp 1624047346
transform -1 0 39836 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1624047346
transform 1 0 39192 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_412
timestamp 1624047346
transform 1 0 39008 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_416
timestamp 1624047346
transform 1 0 39376 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_407
timestamp 1624047346
transform 1 0 38548 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_414
timestamp 1624047346
transform 1 0 39192 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1624047346
transform 1 0 40480 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A
timestamp 1624047346
transform -1 0 40756 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_428
timestamp 1624047346
transform 1 0 40480 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_421
timestamp 1624047346
transform 1 0 39836 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_427
timestamp 1624047346
transform 1 0 40388 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_431
timestamp 1624047346
transform 1 0 40756 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_440
timestamp 1624047346
transform 1 0 41584 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_452
timestamp 1624047346
transform 1 0 42688 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_443
timestamp 1624047346
transform 1 0 41860 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1624047346
transform 1 0 43056 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_457
timestamp 1624047346
transform 1 0 43148 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_469
timestamp 1624047346
transform 1 0 44252 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_455
timestamp 1624047346
transform 1 0 42964 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_467
timestamp 1624047346
transform 1 0 44068 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1624047346
transform 1 0 45724 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_481
timestamp 1624047346
transform 1 0 45356 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_479
timestamp 1624047346
transform 1 0 45172 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_40_486
timestamp 1624047346
transform 1 0 45816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_493
timestamp 1624047346
transform 1 0 46460 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_505
timestamp 1624047346
transform 1 0 47564 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_498
timestamp 1624047346
transform 1 0 46920 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1624047346
transform 1 0 48300 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_514
timestamp 1624047346
transform 1 0 48392 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_510
timestamp 1624047346
transform 1 0 48024 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_526
timestamp 1624047346
transform 1 0 49496 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_538
timestamp 1624047346
transform 1 0 50600 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_522
timestamp 1624047346
transform 1 0 49128 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_534
timestamp 1624047346
transform 1 0 50232 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1624047346
transform 1 0 50968 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_550
timestamp 1624047346
transform 1 0 51704 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_543
timestamp 1624047346
transform 1 0 51060 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_555
timestamp 1624047346
transform 1 0 52164 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1624047346
transform 1 0 53544 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_562
timestamp 1624047346
transform 1 0 52808 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_571
timestamp 1624047346
transform 1 0 53636 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_567
timestamp 1624047346
transform 1 0 53268 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_583
timestamp 1624047346
transform 1 0 54740 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_579
timestamp 1624047346
transform 1 0 54372 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1624047346
transform 1 0 56212 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output216_A
timestamp 1624047346
transform -1 0 57040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_595
timestamp 1624047346
transform 1 0 55844 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_591
timestamp 1624047346
transform 1 0 55476 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_600
timestamp 1624047346
transform 1 0 56304 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_608
timestamp 1624047346
transform 1 0 57040 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_607
timestamp 1624047346
transform 1 0 56948 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_614
timestamp 1624047346
transform 1 0 57592 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_614
timestamp 1624047346
transform 1 0 57592 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_611
timestamp 1624047346
transform 1 0 57316 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1624047346
transform -1 0 57592 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1624047346
transform -1 0 57592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 1624047346
transform -1 0 58236 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1624047346
transform -1 0 58236 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1624047346
transform 1 0 58236 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_621
timestamp 1624047346
transform 1 0 58236 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1624047346
transform -1 0 58880 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1624047346
transform -1 0 58880 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1624047346
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1624047346
transform -1 0 1564 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output236_A
timestamp 1624047346
transform -1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_5
timestamp 1624047346
transform 1 0 1564 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_11
timestamp 1624047346
transform 1 0 2116 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1624047346
transform 1 0 3220 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1624047346
transform 1 0 4324 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1624047346
transform 1 0 5428 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1624047346
transform 1 0 6348 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_55
timestamp 1624047346
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_58
timestamp 1624047346
transform 1 0 6440 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_70
timestamp 1624047346
transform 1 0 7544 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_82
timestamp 1624047346
transform 1 0 8648 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_94
timestamp 1624047346
transform 1 0 9752 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1624047346
transform 1 0 11592 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_106
timestamp 1624047346
transform 1 0 10856 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_115
timestamp 1624047346
transform 1 0 11684 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_127
timestamp 1624047346
transform 1 0 12788 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1624047346
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_151
timestamp 1624047346
transform 1 0 14996 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_163
timestamp 1624047346
transform 1 0 16100 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1624047346
transform 1 0 16836 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_172
timestamp 1624047346
transform 1 0 16928 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1624047346
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1624047346
transform 1 0 19136 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1624047346
transform 1 0 20240 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1624047346
transform 1 0 22080 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_220
timestamp 1624047346
transform 1 0 21344 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_229
timestamp 1624047346
transform 1 0 22172 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1624047346
transform -1 0 23644 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_241
timestamp 1624047346
transform 1 0 23276 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1624047346
transform 1 0 23644 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1624047346
transform 1 0 24748 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_269
timestamp 1624047346
transform 1 0 25852 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1624047346
transform 1 0 27324 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_281
timestamp 1624047346
transform 1 0 26956 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_286
timestamp 1624047346
transform 1 0 27416 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _166_
timestamp 1624047346
transform -1 0 29072 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_298
timestamp 1624047346
transform 1 0 28520 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_304
timestamp 1624047346
transform 1 0 29072 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_316
timestamp 1624047346
transform 1 0 30176 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_328
timestamp 1624047346
transform 1 0 31280 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1624047346
transform 1 0 32568 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_340
timestamp 1624047346
transform 1 0 32384 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_343
timestamp 1624047346
transform 1 0 32660 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1624047346
transform -1 0 34592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_355
timestamp 1624047346
transform 1 0 33764 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_361
timestamp 1624047346
transform 1 0 34316 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_364
timestamp 1624047346
transform 1 0 34592 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1624047346
transform 1 0 36616 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_376
timestamp 1624047346
transform 1 0 35696 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_384
timestamp 1624047346
transform 1 0 36432 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1624047346
transform 1 0 37812 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A
timestamp 1624047346
transform 1 0 37168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A
timestamp 1624047346
transform -1 0 38088 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_388
timestamp 1624047346
transform 1 0 36800 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_394
timestamp 1624047346
transform 1 0 37352 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_398
timestamp 1624047346
transform 1 0 37720 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_402
timestamp 1624047346
transform 1 0 38088 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__A
timestamp 1624047346
transform -1 0 38640 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__B
timestamp 1624047346
transform -1 0 39192 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__B
timestamp 1624047346
transform -1 0 39744 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_408
timestamp 1624047346
transform 1 0 38640 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_414
timestamp 1624047346
transform 1 0 39192 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_420
timestamp 1624047346
transform 1 0 39744 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__S
timestamp 1624047346
transform 1 0 40112 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_426
timestamp 1624047346
transform 1 0 40296 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_438
timestamp 1624047346
transform 1 0 41400 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_450
timestamp 1624047346
transform 1 0 42504 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1624047346
transform 1 0 43056 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_457
timestamp 1624047346
transform 1 0 43148 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_469
timestamp 1624047346
transform 1 0 44252 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_481
timestamp 1624047346
transform 1 0 45356 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_493
timestamp 1624047346
transform 1 0 46460 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_505
timestamp 1624047346
transform 1 0 47564 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1624047346
transform 1 0 48300 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_514
timestamp 1624047346
transform 1 0 48392 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_526
timestamp 1624047346
transform 1 0 49496 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_538
timestamp 1624047346
transform 1 0 50600 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_550
timestamp 1624047346
transform 1 0 51704 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1624047346
transform 1 0 53544 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_562
timestamp 1624047346
transform 1 0 52808 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_571
timestamp 1624047346
transform 1 0 53636 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_583
timestamp 1624047346
transform 1 0 54740 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output200_A
timestamp 1624047346
transform 1 0 56856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__S
timestamp 1624047346
transform 1 0 56304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_595
timestamp 1624047346
transform 1 0 55844 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_599
timestamp 1624047346
transform 1 0 56212 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_602
timestamp 1624047346
transform 1 0 56488 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1624047346
transform -1 0 58236 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624047346
transform -1 0 57592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_608
timestamp 1624047346
transform 1 0 57040 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_614
timestamp 1624047346
transform 1 0 57592 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_621
timestamp 1624047346
transform 1 0 58236 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1624047346
transform -1 0 58880 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1624047346
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output211
timestamp 1624047346
transform -1 0 1748 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1624047346
transform -1 0 2300 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_7
timestamp 1624047346
transform 1 0 1748 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_13
timestamp 1624047346
transform 1 0 2300 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1624047346
transform 1 0 3772 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output227_A
timestamp 1624047346
transform -1 0 2852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_19
timestamp 1624047346
transform 1 0 2852 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_27
timestamp 1624047346
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_30
timestamp 1624047346
transform 1 0 3864 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_42
timestamp 1624047346
transform 1 0 4968 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_54
timestamp 1624047346
transform 1 0 6072 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_66
timestamp 1624047346
transform 1 0 7176 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_78
timestamp 1624047346
transform 1 0 8280 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1624047346
transform 1 0 9016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__A1
timestamp 1624047346
transform -1 0 10120 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_87
timestamp 1624047346
transform 1 0 9108 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_95
timestamp 1624047346
transform 1 0 9844 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_98
timestamp 1624047346
transform 1 0 10120 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_110
timestamp 1624047346
transform 1 0 11224 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_122
timestamp 1624047346
transform 1 0 12328 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_134
timestamp 1624047346
transform 1 0 13432 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1624047346
transform 1 0 14260 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_142
timestamp 1624047346
transform 1 0 14168 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_144
timestamp 1624047346
transform 1 0 14352 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_156
timestamp 1624047346
transform 1 0 15456 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_168
timestamp 1624047346
transform 1 0 16560 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1624047346
transform -1 0 17940 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__S
timestamp 1624047346
transform 1 0 16928 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_174
timestamp 1624047346
transform 1 0 17112 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_180
timestamp 1624047346
transform 1 0 17664 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_183
timestamp 1624047346
transform 1 0 17940 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1624047346
transform 1 0 19504 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__S
timestamp 1624047346
transform 1 0 18768 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_191
timestamp 1624047346
transform 1 0 18676 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_194
timestamp 1624047346
transform 1 0 18952 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_201
timestamp 1624047346
transform 1 0 19596 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_213
timestamp 1624047346
transform 1 0 20700 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_225
timestamp 1624047346
transform 1 0 21804 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_237
timestamp 1624047346
transform 1 0 22908 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_249
timestamp 1624047346
transform 1 0 24012 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1624047346
transform 1 0 24748 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_258
timestamp 1624047346
transform 1 0 24840 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_270
timestamp 1624047346
transform 1 0 25944 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_282
timestamp 1624047346
transform 1 0 27048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_294
timestamp 1624047346
transform 1 0 28152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1624047346
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_306
timestamp 1624047346
transform 1 0 29256 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_315
timestamp 1624047346
transform 1 0 30084 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_327
timestamp 1624047346
transform 1 0 31188 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__S
timestamp 1624047346
transform 1 0 33396 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1624047346
transform 1 0 32292 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_353
timestamp 1624047346
transform 1 0 33580 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__A
timestamp 1624047346
transform 1 0 34224 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_359
timestamp 1624047346
transform 1 0 34132 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_362
timestamp 1624047346
transform 1 0 34408 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_370
timestamp 1624047346
transform 1 0 35144 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1624047346
transform 1 0 35236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__223__A
timestamp 1624047346
transform 1 0 36064 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1624047346
transform -1 0 35696 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_372
timestamp 1624047346
transform 1 0 35328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_376
timestamp 1624047346
transform 1 0 35696 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_382
timestamp 1624047346
transform 1 0 36248 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _251_
timestamp 1624047346
transform 1 0 38180 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__B
timestamp 1624047346
transform 1 0 37628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1624047346
transform 1 0 36892 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_388
timestamp 1624047346
transform 1 0 36800 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_391
timestamp 1624047346
transform 1 0 37076 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_399
timestamp 1624047346
transform 1 0 37812 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _247_
timestamp 1624047346
transform -1 0 39284 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A1
timestamp 1624047346
transform -1 0 39836 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_408
timestamp 1624047346
transform 1 0 38640 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_415
timestamp 1624047346
transform 1 0 39284 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1624047346
transform 1 0 40480 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__S
timestamp 1624047346
transform 1 0 40572 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_421
timestamp 1624047346
transform 1 0 39836 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_427
timestamp 1624047346
transform 1 0 40388 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_431
timestamp 1624047346
transform 1 0 40756 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_443
timestamp 1624047346
transform 1 0 41860 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_455
timestamp 1624047346
transform 1 0 42964 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_467
timestamp 1624047346
transform 1 0 44068 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1624047346
transform 1 0 45724 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_479
timestamp 1624047346
transform 1 0 45172 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_486
timestamp 1624047346
transform 1 0 45816 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_498
timestamp 1624047346
transform 1 0 46920 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_510
timestamp 1624047346
transform 1 0 48024 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_522
timestamp 1624047346
transform 1 0 49128 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_534
timestamp 1624047346
transform 1 0 50232 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1624047346
transform 1 0 50968 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_543
timestamp 1624047346
transform 1 0 51060 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_555
timestamp 1624047346
transform 1 0 52164 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_567
timestamp 1624047346
transform 1 0 53268 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_579
timestamp 1624047346
transform 1 0 54372 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1624047346
transform 1 0 56212 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624047346
transform -1 0 56856 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output169_A
timestamp 1624047346
transform 1 0 55660 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_591
timestamp 1624047346
transform 1 0 55476 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_595
timestamp 1624047346
transform 1 0 55844 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_600
timestamp 1624047346
transform 1 0 56304 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_606
timestamp 1624047346
transform 1 0 56856 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1624047346
transform -1 0 57500 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output216
timestamp 1624047346
transform 1 0 57868 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1624047346
transform 1 0 57500 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1624047346
transform 1 0 58236 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1624047346
transform -1 0 58880 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1624047346
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output158
timestamp 1624047346
transform -1 0 1748 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1624047346
transform -1 0 2760 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_7
timestamp 1624047346
transform 1 0 1748 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1624047346
transform 1 0 2484 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1624047346
transform 1 0 3404 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_18
timestamp 1624047346
transform 1 0 2760 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_24
timestamp 1624047346
transform 1 0 3312 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1624047346
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A1
timestamp 1624047346
transform 1 0 5060 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__S
timestamp 1624047346
transform 1 0 5612 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_39
timestamp 1624047346
transform 1 0 4692 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_45
timestamp 1624047346
transform 1 0 5244 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1624047346
transform 1 0 6348 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_51
timestamp 1624047346
transform 1 0 5796 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_58
timestamp 1624047346
transform 1 0 6440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__278__S
timestamp 1624047346
transform 1 0 8648 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_70
timestamp 1624047346
transform 1 0 7544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_84
timestamp 1624047346
transform 1 0 8832 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _086_
timestamp 1624047346
transform 1 0 9752 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1624047346
transform 1 0 10396 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1624047346
transform 1 0 9200 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_90
timestamp 1624047346
transform 1 0 9384 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_97
timestamp 1624047346
transform 1 0 10028 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1624047346
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A
timestamp 1624047346
transform 1 0 11684 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__S
timestamp 1624047346
transform 1 0 10948 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_103
timestamp 1624047346
transform 1 0 10580 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_109
timestamp 1624047346
transform 1 0 11132 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_113
timestamp 1624047346
transform 1 0 11500 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_117
timestamp 1624047346
transform 1 0 11868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_129
timestamp 1624047346
transform 1 0 12972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_141
timestamp 1624047346
transform 1 0 14076 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_153
timestamp 1624047346
transform 1 0 15180 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_165
timestamp 1624047346
transform 1 0 16284 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1624047346
transform 1 0 16836 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1624047346
transform 1 0 17480 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__A0
timestamp 1624047346
transform 1 0 16928 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_174
timestamp 1624047346
transform 1 0 17112 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_181
timestamp 1624047346
transform 1 0 17756 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_185
timestamp 1624047346
transform 1 0 18124 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _083_
timestamp 1624047346
transform 1 0 19412 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624047346
transform -1 0 18400 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__B
timestamp 1624047346
transform 1 0 18768 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_188
timestamp 1624047346
transform 1 0 18400 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_194
timestamp 1624047346
transform 1 0 18952 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_198
timestamp 1624047346
transform 1 0 19320 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1624047346
transform 1 0 19688 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__189__A
timestamp 1624047346
transform -1 0 21344 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__276__A0
timestamp 1624047346
transform -1 0 20240 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_208
timestamp 1624047346
transform 1 0 20240 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_216
timestamp 1624047346
transform 1 0 20976 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1624047346
transform 1 0 22080 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_220
timestamp 1624047346
transform 1 0 21344 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_229
timestamp 1624047346
transform 1 0 22172 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output152_A
timestamp 1624047346
transform 1 0 23552 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_241
timestamp 1624047346
transform 1 0 23276 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_246
timestamp 1624047346
transform 1 0 23736 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_258
timestamp 1624047346
transform 1 0 24840 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _134_
timestamp 1624047346
transform -1 0 26956 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1624047346
transform 1 0 27324 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_270
timestamp 1624047346
transform 1 0 25944 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1624047346
transform 1 0 26956 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_286
timestamp 1624047346
transform 1 0 27416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_298
timestamp 1624047346
transform 1 0 28520 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__S
timestamp 1624047346
transform 1 0 29256 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_308
timestamp 1624047346
transform 1 0 29440 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_320
timestamp 1624047346
transform 1 0 30544 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_332
timestamp 1624047346
transform 1 0 31648 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1624047346
transform 1 0 32568 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A1
timestamp 1624047346
transform -1 0 33488 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__S
timestamp 1624047346
transform 1 0 32660 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_340
timestamp 1624047346
transform 1 0 32384 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_345
timestamp 1624047346
transform 1 0 32844 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_349
timestamp 1624047346
transform 1 0 33212 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_352
timestamp 1624047346
transform 1 0 33488 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1624047346
transform -1 0 35236 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624047346
transform -1 0 34592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1624047346
transform -1 0 34040 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_358
timestamp 1624047346
transform 1 0 34040 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_364
timestamp 1624047346
transform 1 0 34592 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624047346
transform -1 0 36800 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1624047346
transform -1 0 35788 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_371
timestamp 1624047346
transform 1 0 35236 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_377
timestamp 1624047346
transform 1 0 35788 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_385
timestamp 1624047346
transform 1 0 36524 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_1  _183_
timestamp 1624047346
transform 1 0 37168 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _250_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624047346
transform 1 0 38272 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1624047346
transform 1 0 37812 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1624047346
transform 1 0 36800 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_395
timestamp 1624047346
transform 1 0 37444 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_400
timestamp 1624047346
transform 1 0 37904 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1624047346
transform -1 0 39376 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__270__A0
timestamp 1624047346
transform 1 0 39744 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_409
timestamp 1624047346
transform 1 0 38732 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_413
timestamp 1624047346
transform 1 0 39100 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_416
timestamp 1624047346
transform 1 0 39376 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624047346
transform -1 0 41124 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__282__A1
timestamp 1624047346
transform 1 0 40296 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_422
timestamp 1624047346
transform 1 0 39928 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_428
timestamp 1624047346
transform 1 0 40480 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_432
timestamp 1624047346
transform 1 0 40848 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_435
timestamp 1624047346
transform 1 0 41124 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1624047346
transform -1 0 41676 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_441
timestamp 1624047346
transform 1 0 41676 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_453
timestamp 1624047346
transform 1 0 42780 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1624047346
transform 1 0 43056 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_457
timestamp 1624047346
transform 1 0 43148 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_469
timestamp 1624047346
transform 1 0 44252 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_481
timestamp 1624047346
transform 1 0 45356 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_493
timestamp 1624047346
transform 1 0 46460 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1624047346
transform 1 0 47564 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1624047346
transform 1 0 48300 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_514
timestamp 1624047346
transform 1 0 48392 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_526
timestamp 1624047346
transform 1 0 49496 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_538
timestamp 1624047346
transform 1 0 50600 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_550
timestamp 1624047346
transform 1 0 51704 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1624047346
transform 1 0 53544 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_562
timestamp 1624047346
transform 1 0 52808 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_571
timestamp 1624047346
transform 1 0 53636 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output205_A
timestamp 1624047346
transform 1 0 54924 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_583
timestamp 1624047346
transform 1 0 54740 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_587
timestamp 1624047346
transform 1 0 55108 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624047346
transform -1 0 56764 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A0
timestamp 1624047346
transform -1 0 56212 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output143_A
timestamp 1624047346
transform -1 0 55660 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_593
timestamp 1624047346
transform 1 0 55660 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_599
timestamp 1624047346
transform 1 0 56212 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_605
timestamp 1624047346
transform 1 0 56764 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _269_
timestamp 1624047346
transform 1 0 57132 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_43_618
timestamp 1624047346
transform 1 0 57960 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1624047346
transform -1 0 58880 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_624
timestamp 1624047346
transform 1 0 58512 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1624047346
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1624047346
transform 1 0 2300 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output236
timestamp 1624047346
transform -1 0 1748 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_7
timestamp 1624047346
transform 1 0 1748 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_16
timestamp 1624047346
transform 1 0 2576 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1624047346
transform 1 0 3772 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624047346
transform -1 0 3128 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1624047346
transform 1 0 3128 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_28
timestamp 1624047346
transform 1 0 3680 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_30
timestamp 1624047346
transform 1 0 3864 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output233
timestamp 1624047346
transform -1 0 4600 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624047346
transform -1 0 5336 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A0
timestamp 1624047346
transform -1 0 5888 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_38
timestamp 1624047346
transform 1 0 4600 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_46
timestamp 1624047346
transform 1 0 5336 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__S
timestamp 1624047346
transform 1 0 6256 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_52
timestamp 1624047346
transform 1 0 5888 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_58
timestamp 1624047346
transform 1 0 6440 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_66
timestamp 1624047346
transform 1 0 7176 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1624047346
transform -1 0 7544 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1624047346
transform -1 0 8648 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output210_A
timestamp 1624047346
transform -1 0 8096 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_70
timestamp 1624047346
transform 1 0 7544 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_76
timestamp 1624047346
transform 1 0 8096 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_82
timestamp 1624047346
transform 1 0 8648 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 1624047346
transform 1 0 10212 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1624047346
transform 1 0 9016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output231
timestamp 1624047346
transform -1 0 9844 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_87
timestamp 1624047346
transform 1 0 9108 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_95
timestamp 1624047346
transform 1 0 9844 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _283_
timestamp 1624047346
transform 1 0 11132 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_44_102
timestamp 1624047346
transform 1 0 10488 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_108
timestamp 1624047346
transform 1 0 11040 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1624047346
transform 1 0 12328 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624047346
transform -1 0 13156 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_118
timestamp 1624047346
transform 1 0 11960 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_125
timestamp 1624047346
transform 1 0 12604 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_131
timestamp 1624047346
transform 1 0 13156 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1624047346
transform 1 0 14260 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 1624047346
transform 1 0 13524 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_137
timestamp 1624047346
transform 1 0 13708 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_44_144
timestamp 1624047346
transform 1 0 14352 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624047346
transform -1 0 16008 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1624047346
transform -1 0 16560 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output214_A
timestamp 1624047346
transform 1 0 15272 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_152
timestamp 1624047346
transform 1 0 15088 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_156
timestamp 1624047346
transform 1 0 15456 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_162
timestamp 1624047346
transform 1 0 16008 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_168
timestamp 1624047346
transform 1 0 16560 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _115_
timestamp 1624047346
transform -1 0 18032 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _203_
timestamp 1624047346
transform 1 0 16928 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_175
timestamp 1624047346
transform 1 0 17204 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_184
timestamp 1624047346
transform 1 0 18032 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1624047346
transform 1 0 19504 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1624047346
transform 1 0 18860 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1624047346
transform -1 0 19780 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_192
timestamp 1624047346
transform 1 0 18768 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_196
timestamp 1624047346
transform 1 0 19136 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output222
timestamp 1624047346
transform -1 0 20608 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output229
timestamp 1624047346
transform -1 0 21528 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_203
timestamp 1624047346
transform 1 0 19780 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_207
timestamp 1624047346
transform 1 0 20148 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_212
timestamp 1624047346
transform 1 0 20608 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp 1624047346
transform 1 0 22264 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_222
timestamp 1624047346
transform 1 0 21528 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_233
timestamp 1624047346
transform 1 0 22540 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1624047346
transform -1 0 23920 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A
timestamp 1624047346
transform 1 0 23092 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_241
timestamp 1624047346
transform 1 0 23276 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_245
timestamp 1624047346
transform 1 0 23644 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_248
timestamp 1624047346
transform 1 0 23920 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1624047346
transform 1 0 24748 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624047346
transform -1 0 25944 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A
timestamp 1624047346
transform -1 0 25392 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_256
timestamp 1624047346
transform 1 0 24656 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_258
timestamp 1624047346
transform 1 0 24840 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_264
timestamp 1624047346
transform 1 0 25392 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _133_
timestamp 1624047346
transform -1 0 27232 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1624047346
transform -1 0 26588 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_270
timestamp 1624047346
transform 1 0 25944 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_277
timestamp 1624047346
transform 1 0 26588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_284
timestamp 1624047346
transform 1 0 27232 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output192
timestamp 1624047346
transform -1 0 27968 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1624047346
transform -1 0 28520 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_292
timestamp 1624047346
transform 1 0 27968 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_298
timestamp 1624047346
transform 1 0 28520 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _131_
timestamp 1624047346
transform -1 0 29624 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1624047346
transform 1 0 29992 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1624047346
transform 1 0 30452 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_306
timestamp 1624047346
transform 1 0 29256 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_310
timestamp 1624047346
transform 1 0 29624 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_315
timestamp 1624047346
transform 1 0 30084 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624047346
transform -1 0 32200 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1624047346
transform -1 0 31280 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_322
timestamp 1624047346
transform 1 0 30728 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_328
timestamp 1624047346
transform 1 0 31280 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  output235
timestamp 1624047346
transform -1 0 33488 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__A0
timestamp 1624047346
transform -1 0 32752 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_338
timestamp 1624047346
transform 1 0 32200 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_344
timestamp 1624047346
transform 1 0 32752 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_352
timestamp 1624047346
transform 1 0 33488 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1624047346
transform 1 0 34592 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1624047346
transform -1 0 34224 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_356
timestamp 1624047346
transform 1 0 33856 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1624047346
transform 1 0 34224 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_367
timestamp 1624047346
transform 1 0 34868 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1624047346
transform 1 0 35696 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1624047346
transform 1 0 35236 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1624047346
transform 1 0 36340 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_372
timestamp 1624047346
transform 1 0 35328 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_379
timestamp 1624047346
transform 1 0 35972 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_386
timestamp 1624047346
transform 1 0 36616 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _207_
timestamp 1624047346
transform 1 0 37352 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _270_
timestamp 1624047346
transform 1 0 38180 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_44_399
timestamp 1624047346
transform 1 0 37812 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1624047346
transform -1 0 39652 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_412
timestamp 1624047346
transform 1 0 39008 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_419
timestamp 1624047346
transform 1 0 39652 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1624047346
transform 1 0 40480 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 1624047346
transform -1 0 41216 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_427
timestamp 1624047346
transform 1 0 40388 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_429
timestamp 1624047346
transform 1 0 40572 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_436
timestamp 1624047346
transform 1 0 41216 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624047346
transform -1 0 41768 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output225_A
timestamp 1624047346
transform 1 0 42228 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_442
timestamp 1624047346
transform 1 0 41768 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_446
timestamp 1624047346
transform 1 0 42136 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_449
timestamp 1624047346
transform 1 0 42412 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output208_A
timestamp 1624047346
transform 1 0 44436 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_461
timestamp 1624047346
transform 1 0 43516 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_469
timestamp 1624047346
transform 1 0 44252 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1624047346
transform 1 0 45724 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output139_A
timestamp 1624047346
transform -1 0 46000 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_473
timestamp 1624047346
transform 1 0 44620 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_488
timestamp 1624047346
transform 1 0 46000 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_500
timestamp 1624047346
transform 1 0 47104 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_512
timestamp 1624047346
transform 1 0 48208 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output162_A
timestamp 1624047346
transform -1 0 49588 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output202_A
timestamp 1624047346
transform -1 0 50140 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_524
timestamp 1624047346
transform 1 0 49312 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_527
timestamp 1624047346
transform 1 0 49588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_533
timestamp 1624047346
transform 1 0 50140 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1624047346
transform 1 0 50968 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1624047346
transform -1 0 51612 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_541
timestamp 1624047346
transform 1 0 50876 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_543
timestamp 1624047346
transform 1 0 51060 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_549
timestamp 1624047346
transform 1 0 51612 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_561
timestamp 1624047346
transform 1 0 52716 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1624047346
transform -1 0 55292 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output145_A
timestamp 1624047346
transform 1 0 54556 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_573
timestamp 1624047346
transform 1 0 53820 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_583
timestamp 1624047346
transform 1 0 54740 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_589
timestamp 1624047346
transform 1 0 55292 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1624047346
transform 1 0 56212 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output205
timestamp 1624047346
transform -1 0 57040 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1624047346
transform -1 0 55844 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_595
timestamp 1624047346
transform 1 0 55844 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_600
timestamp 1624047346
transform 1 0 56304 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output200
timestamp 1624047346
transform 1 0 57868 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_608
timestamp 1624047346
transform 1 0 57040 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_616
timestamp 1624047346
transform 1 0 57776 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_621
timestamp 1624047346
transform 1 0 58236 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1624047346
transform -1 0 58880 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1624047346
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input99
timestamp 1624047346
transform 1 0 1380 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output227
timestamp 1624047346
transform -1 0 2484 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_7
timestamp 1624047346
transform 1 0 1748 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_15
timestamp 1624047346
transform 1 0 2484 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _279_
timestamp 1624047346
transform 1 0 4140 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1624047346
transform -1 0 3128 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624047346
transform -1 0 3680 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_22
timestamp 1624047346
transform 1 0 3128 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_28
timestamp 1624047346
transform 1 0 3680 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_32
timestamp 1624047346
transform 1 0 4048 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1624047346
transform 1 0 5336 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_42
timestamp 1624047346
transform 1 0 4968 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_49
timestamp 1624047346
transform 1 0 5612 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1624047346
transform 1 0 6348 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output210
timestamp 1624047346
transform -1 0 7176 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_58
timestamp 1624047346
transform 1 0 6440 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_66
timestamp 1624047346
transform 1 0 7176 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 1624047346
transform 1 0 7544 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 1624047346
transform 1 0 8464 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_73
timestamp 1624047346
transform 1 0 7820 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_79
timestamp 1624047346
transform 1 0 8372 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_83
timestamp 1624047346
transform 1 0 8740 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _190_
timestamp 1624047346
transform -1 0 11224 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1624047346
transform -1 0 9936 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_96
timestamp 1624047346
transform 1 0 9936 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_100
timestamp 1624047346
transform 1 0 10304 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1624047346
transform 1 0 11592 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_110
timestamp 1624047346
transform 1 0 11224 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_115
timestamp 1624047346
transform 1 0 11684 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1624047346
transform 1 0 12052 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1624047346
transform -1 0 13156 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_122
timestamp 1624047346
transform 1 0 12328 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_131
timestamp 1624047346
transform 1 0 13156 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1624047346
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624047346
transform -1 0 13708 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1624047346
transform -1 0 15088 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_137
timestamp 1624047346
transform 1 0 13708 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_146
timestamp 1624047346
transform 1 0 14536 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1624047346
transform -1 0 16468 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1624047346
transform -1 0 15824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_152
timestamp 1624047346
transform 1 0 15088 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_156
timestamp 1624047346
transform 1 0 15456 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_160
timestamp 1624047346
transform 1 0 15824 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_167
timestamp 1624047346
transform 1 0 16468 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _264_
timestamp 1624047346
transform -1 0 18124 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1624047346
transform 1 0 16836 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_172
timestamp 1624047346
transform 1 0 16928 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_185
timestamp 1624047346
transform 1 0 18124 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp 1624047346
transform -1 0 19780 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_45_193
timestamp 1624047346
transform 1 0 18860 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _189_
timestamp 1624047346
transform -1 0 21160 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_45_203
timestamp 1624047346
transform 1 0 19780 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_218
timestamp 1624047346
transform 1 0 21160 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1624047346
transform 1 0 22080 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output196
timestamp 1624047346
transform -1 0 22908 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1624047346
transform -1 0 21712 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_224
timestamp 1624047346
transform 1 0 21712 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_229
timestamp 1624047346
transform 1 0 22172 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _201_
timestamp 1624047346
transform 1 0 23276 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1624047346
transform 1 0 23920 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_237
timestamp 1624047346
transform 1 0 22908 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_244
timestamp 1624047346
transform 1 0 23552 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_251
timestamp 1624047346
transform 1 0 24196 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input94
timestamp 1624047346
transform 1 0 25300 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1624047346
transform -1 0 24932 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_259
timestamp 1624047346
transform 1 0 24932 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_266
timestamp 1624047346
transform 1 0 25576 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _218_
timestamp 1624047346
transform -1 0 26220 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1624047346
transform 1 0 27324 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output209
timestamp 1624047346
transform 1 0 26588 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_273
timestamp 1624047346
transform 1 0 26220 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1624047346
transform 1 0 26956 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_286
timestamp 1624047346
transform 1 0 27416 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _217_
timestamp 1624047346
transform 1 0 27784 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  output195
timestamp 1624047346
transform 1 0 28704 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_295
timestamp 1624047346
transform 1 0 28244 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_299
timestamp 1624047346
transform 1 0 28612 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _274_
timestamp 1624047346
transform 1 0 29440 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_304
timestamp 1624047346
transform 1 0 29072 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_317
timestamp 1624047346
transform 1 0 30268 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1624047346
transform -1 0 32016 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output190
timestamp 1624047346
transform -1 0 31188 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_327
timestamp 1624047346
transform 1 0 31188 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_336
timestamp 1624047346
transform 1 0 32016 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _254_
timestamp 1624047346
transform 1 0 33028 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1624047346
transform 1 0 32568 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_343
timestamp 1624047346
transform 1 0 32660 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _198_
timestamp 1624047346
transform 1 0 34408 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_45_356
timestamp 1624047346
transform 1 0 33856 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_367
timestamp 1624047346
transform 1 0 34868 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _143_
timestamp 1624047346
transform -1 0 36892 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _223_
timestamp 1624047346
transform 1 0 35236 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_45_380
timestamp 1624047346
transform 1 0 36064 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1624047346
transform 1 0 37812 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1624047346
transform -1 0 38548 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624047346
transform -1 0 37444 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_389
timestamp 1624047346
transform 1 0 36892 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_395
timestamp 1624047346
transform 1 0 37444 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_400
timestamp 1624047346
transform 1 0 37904 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  repeater246
timestamp 1624047346
transform -1 0 40020 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_407
timestamp 1624047346
transform 1 0 38548 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1624047346
transform 1 0 41124 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output221
timestamp 1624047346
transform -1 0 40756 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_423
timestamp 1624047346
transform 1 0 40020 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_431
timestamp 1624047346
transform 1 0 40756 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output225
timestamp 1624047346
transform -1 0 42228 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_438
timestamp 1624047346
transform 1 0 41400 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_442
timestamp 1624047346
transform 1 0 41768 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_447
timestamp 1624047346
transform 1 0 42228 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1624047346
transform 1 0 43056 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1624047346
transform 1 0 44068 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater246_A
timestamp 1624047346
transform -1 0 43332 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_455
timestamp 1624047346
transform 1 0 42964 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_459
timestamp 1624047346
transform 1 0 43332 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_469
timestamp 1624047346
transform 1 0 44252 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1624047346
transform -1 0 45632 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output208
timestamp 1624047346
transform -1 0 44988 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624047346
transform -1 0 46184 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_477
timestamp 1624047346
transform 1 0 44988 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_484
timestamp 1624047346
transform 1 0 45632 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output244
timestamp 1624047346
transform 1 0 47564 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_490
timestamp 1624047346
transform 1 0 46184 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_502
timestamp 1624047346
transform 1 0 47288 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1624047346
transform 1 0 48300 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624047346
transform -1 0 48852 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_509
timestamp 1624047346
transform 1 0 47932 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_514
timestamp 1624047346
transform 1 0 48392 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_519
timestamp 1624047346
transform 1 0 48852 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output184
timestamp 1624047346
transform -1 0 50508 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output202
timestamp 1624047346
transform 1 0 49404 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_529
timestamp 1624047346
transform 1 0 49772 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_537
timestamp 1624047346
transform 1 0 50508 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  output212
timestamp 1624047346
transform -1 0 51428 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624047346
transform -1 0 52256 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_547
timestamp 1624047346
transform 1 0 51428 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_553
timestamp 1624047346
transform 1 0 51980 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1624047346
transform 1 0 53544 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624047346
transform -1 0 53912 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_556
timestamp 1624047346
transform 1 0 52256 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_568
timestamp 1624047346
transform 1 0 53360 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_571
timestamp 1624047346
transform 1 0 53636 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1624047346
transform -1 0 55108 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1624047346
transform 1 0 54372 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_574
timestamp 1624047346
transform 1 0 53912 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_578
timestamp 1624047346
transform 1 0 54280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_581
timestamp 1624047346
transform 1 0 54556 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_587
timestamp 1624047346
transform 1 0 55108 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input116
timestamp 1624047346
transform -1 0 55752 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output169
timestamp 1624047346
transform -1 0 56488 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_594
timestamp 1624047346
transform 1 0 55752 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_602
timestamp 1624047346
transform 1 0 56488 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1624047346
transform -1 0 58236 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output145
timestamp 1624047346
transform 1 0 57132 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_608
timestamp 1624047346
transform 1 0 57040 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_613
timestamp 1624047346
transform 1 0 57500 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1624047346
transform 1 0 58236 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1624047346
transform -1 0 58880 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1624047346
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1624047346
transform 1 0 1380 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output167
timestamp 1624047346
transform 1 0 2300 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_7
timestamp 1624047346
transform 1 0 1748 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1624047346
transform 1 0 3772 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output146
timestamp 1624047346
transform -1 0 3404 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_17
timestamp 1624047346
transform 1 0 2668 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_25
timestamp 1624047346
transform 1 0 3404 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_30
timestamp 1624047346
transform 1 0 3864 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp 1624047346
transform 1 0 4232 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output177
timestamp 1624047346
transform -1 0 5888 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_43
timestamp 1624047346
transform 1 0 5060 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_47
timestamp 1624047346
transform 1 0 5428 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1624047346
transform 1 0 6440 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output191
timestamp 1624047346
transform -1 0 7268 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_52
timestamp 1624047346
transform 1 0 5888 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_59
timestamp 1624047346
transform 1 0 6532 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_67
timestamp 1624047346
transform 1 0 7268 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1624047346
transform 1 0 7820 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1624047346
transform -1 0 8740 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_77
timestamp 1624047346
transform 1 0 8188 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_83
timestamp 1624047346
transform 1 0 8740 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1624047346
transform 1 0 9108 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output136
timestamp 1624047346
transform -1 0 10028 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1624047346
transform 1 0 9200 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_92
timestamp 1624047346
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_97
timestamp 1624047346
transform 1 0 10028 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1624047346
transform 1 0 11776 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624047346
transform -1 0 10948 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624047346
transform -1 0 12052 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_107
timestamp 1624047346
transform 1 0 10948 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_115
timestamp 1624047346
transform 1 0 11684 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output137
timestamp 1624047346
transform -1 0 12788 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output136_A
timestamp 1624047346
transform 1 0 13156 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_119
timestamp 1624047346
transform 1 0 12052 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_127
timestamp 1624047346
transform 1 0 12788 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_133
timestamp 1624047346
transform 1 0 13340 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1624047346
transform 1 0 14444 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1624047346
transform -1 0 14076 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output214
timestamp 1624047346
transform -1 0 15272 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1624047346
transform 1 0 14076 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_146
timestamp 1624047346
transform 1 0 14536 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output163
timestamp 1624047346
transform 1 0 16376 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output206
timestamp 1624047346
transform 1 0 15640 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_154
timestamp 1624047346
transform 1 0 15272 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_162
timestamp 1624047346
transform 1 0 16008 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _109_
timestamp 1624047346
transform -1 0 18032 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1624047346
transform 1 0 17112 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_170
timestamp 1624047346
transform 1 0 16744 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_175
timestamp 1624047346
transform 1 0 17204 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_184
timestamp 1624047346
transform 1 0 18032 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1624047346
transform 1 0 18400 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output141
timestamp 1624047346
transform 1 0 19044 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1624047346
transform 1 0 18676 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_199
timestamp 1624047346
transform 1 0 19412 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _084_
timestamp 1624047346
transform 1 0 20240 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1624047346
transform 1 0 19780 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output189
timestamp 1624047346
transform -1 0 21436 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_204
timestamp 1624047346
transform 1 0 19872 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_213
timestamp 1624047346
transform 1 0 20700 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1624047346
transform 1 0 22448 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 1624047346
transform 1 0 21804 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1624047346
transform -1 0 22724 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_221
timestamp 1624047346
transform 1 0 21436 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1624047346
transform 1 0 22080 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_235
timestamp 1624047346
transform 1 0 22724 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1624047346
transform -1 0 24288 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output152
timestamp 1624047346
transform 1 0 23184 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_239
timestamp 1624047346
transform 1 0 23092 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_244
timestamp 1624047346
transform 1 0 23552 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_252
timestamp 1624047346
transform 1 0 24288 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1624047346
transform 1 0 25116 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1624047346
transform -1 0 25944 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_260
timestamp 1624047346
transform 1 0 25024 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_262
timestamp 1624047346
transform 1 0 25208 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _132_
timestamp 1624047346
transform -1 0 27232 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__decap_8  FILLER_46_270
timestamp 1624047346
transform 1 0 25944 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_278
timestamp 1624047346
transform 1 0 26680 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_284
timestamp 1624047346
transform 1 0 27232 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1624047346
transform 1 0 27784 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1624047346
transform 1 0 28520 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624047346
transform -1 0 28152 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_291
timestamp 1624047346
transform 1 0 27876 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_294
timestamp 1624047346
transform 1 0 28152 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_302
timestamp 1624047346
transform 1 0 28888 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1624047346
transform 1 0 30452 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1624047346
transform 1 0 29716 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_310
timestamp 1624047346
transform 1 0 29624 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_315
timestamp 1624047346
transform 1 0 30084 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output170
timestamp 1624047346
transform 1 0 31464 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__274__A0
timestamp 1624047346
transform -1 0 30728 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_322
timestamp 1624047346
transform 1 0 30728 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_334
timestamp 1624047346
transform 1 0 31832 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_2  _260_
timestamp 1624047346
transform 1 0 33580 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1624047346
transform 1 0 33120 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output166
timestamp 1624047346
transform -1 0 32568 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_342
timestamp 1624047346
transform 1 0 32568 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_349
timestamp 1624047346
transform 1 0 33212 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624047346
transform -1 0 35144 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_362
timestamp 1624047346
transform 1 0 34408 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_370
timestamp 1624047346
transform 1 0 35144 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1624047346
transform 1 0 35788 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output135
timestamp 1624047346
transform -1 0 36616 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_376
timestamp 1624047346
transform 1 0 35696 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_378
timestamp 1624047346
transform 1 0 35880 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_386
timestamp 1624047346
transform 1 0 36616 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _205_
timestamp 1624047346
transform -1 0 37812 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__decap_6  FILLER_46_399
timestamp 1624047346
transform 1 0 37812 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_2  _282_
timestamp 1624047346
transform 1 0 38916 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1624047346
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_405
timestamp 1624047346
transform 1 0 38364 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_407
timestamp 1624047346
transform 1 0 38548 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_420
timestamp 1624047346
transform 1 0 39744 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1624047346
transform 1 0 41124 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output153
timestamp 1624047346
transform -1 0 40480 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_428
timestamp 1624047346
transform 1 0 40480 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_434
timestamp 1624047346
transform 1 0 41032 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_436
timestamp 1624047346
transform 1 0 41216 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1624047346
transform 1 0 41584 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output203
timestamp 1624047346
transform 1 0 42320 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_444
timestamp 1624047346
transform 1 0 41952 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_452
timestamp 1624047346
transform 1 0 42688 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1624047346
transform 1 0 43792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1624047346
transform -1 0 44620 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output138
timestamp 1624047346
transform -1 0 43424 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_460
timestamp 1624047346
transform 1 0 43424 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_465
timestamp 1624047346
transform 1 0 43884 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output139
timestamp 1624047346
transform 1 0 45724 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output156
timestamp 1624047346
transform 1 0 44988 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_473
timestamp 1624047346
transform 1 0 44620 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_481
timestamp 1624047346
transform 1 0 45356 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1624047346
transform 1 0 46460 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1624047346
transform -1 0 47288 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_489
timestamp 1624047346
transform 1 0 46092 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_494
timestamp 1624047346
transform 1 0 46552 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_502
timestamp 1624047346
transform 1 0 47288 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1624047346
transform -1 0 48668 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624047346
transform -1 0 47840 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_508
timestamp 1624047346
transform 1 0 47840 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_512
timestamp 1624047346
transform 1 0 48208 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_517
timestamp 1624047346
transform 1 0 48668 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_521
timestamp 1624047346
transform 1 0 49036 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1624047346
transform 1 0 49128 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output162
timestamp 1624047346
transform -1 0 49956 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output179
timestamp 1624047346
transform 1 0 50324 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_523
timestamp 1624047346
transform 1 0 49220 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_531
timestamp 1624047346
transform 1 0 49956 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1624047346
transform 1 0 51796 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1624047346
transform -1 0 51428 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_539
timestamp 1624047346
transform 1 0 50692 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_547
timestamp 1624047346
transform 1 0 51428 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_552
timestamp 1624047346
transform 1 0 51888 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1624047346
transform -1 0 52624 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624047346
transform -1 0 53728 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_560
timestamp 1624047346
transform 1 0 52624 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_572
timestamp 1624047346
transform 1 0 53728 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1624047346
transform 1 0 54464 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624047346
transform -1 0 55292 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_581
timestamp 1624047346
transform 1 0 54556 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_589
timestamp 1624047346
transform 1 0 55292 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1624047346
transform -1 0 56028 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output143
timestamp 1624047346
transform -1 0 56764 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_597
timestamp 1624047346
transform 1 0 56028 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_605
timestamp 1624047346
transform 1 0 56764 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1624047346
transform 1 0 57132 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1624047346
transform -1 0 58236 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_610
timestamp 1624047346
transform 1 0 57224 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_614
timestamp 1624047346
transform 1 0 57592 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_621
timestamp 1624047346
transform 1 0 58236 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1624047346
transform -1 0 58880 0 -1 27744
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 23808 800 23928 6 core_a_data_addr_o[0]
port 0 nsew signal tristate
rlabel metal2 s 54298 29200 54354 30000 6 core_a_data_addr_o[1]
port 1 nsew signal tristate
rlabel metal2 s 43718 29200 43774 30000 6 core_a_data_addr_o[2]
port 2 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 core_a_data_addr_o[3]
port 3 nsew signal tristate
rlabel metal2 s 56138 0 56194 800 6 core_a_data_addr_o[4]
port 4 nsew signal tristate
rlabel metal2 s 29918 29200 29974 30000 6 core_a_data_addr_o[5]
port 5 nsew signal tristate
rlabel metal2 s 10598 29200 10654 30000 6 core_a_data_addr_o[6]
port 6 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 core_a_data_addr_o[7]
port 7 nsew signal tristate
rlabel metal2 s 55218 29200 55274 30000 6 core_a_data_addr_o[8]
port 8 nsew signal tristate
rlabel metal3 s 59200 9528 60000 9648 6 core_a_data_addr_o[9]
port 9 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 core_a_data_be_o[0]
port 10 nsew signal tristate
rlabel metal2 s 23938 29200 23994 30000 6 core_a_data_be_o[1]
port 11 nsew signal tristate
rlabel metal2 s 13818 29200 13874 30000 6 core_a_data_be_o[2]
port 12 nsew signal tristate
rlabel metal3 s 59200 19048 60000 19168 6 core_a_data_be_o[3]
port 13 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 core_a_data_rdata_i[0]
port 14 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 core_a_data_rdata_i[10]
port 15 nsew signal input
rlabel metal3 s 59200 22448 60000 22568 6 core_a_data_rdata_i[11]
port 16 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 core_a_data_rdata_i[12]
port 17 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 core_a_data_rdata_i[13]
port 18 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 core_a_data_rdata_i[14]
port 19 nsew signal input
rlabel metal2 s 51998 29200 52054 30000 6 core_a_data_rdata_i[15]
port 20 nsew signal input
rlabel metal2 s 57978 29200 58034 30000 6 core_a_data_rdata_i[16]
port 21 nsew signal input
rlabel metal3 s 59200 2728 60000 2848 6 core_a_data_rdata_i[17]
port 22 nsew signal input
rlabel metal3 s 59200 26528 60000 26648 6 core_a_data_rdata_i[18]
port 23 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 core_a_data_rdata_i[19]
port 24 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 core_a_data_rdata_i[1]
port 25 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 core_a_data_rdata_i[20]
port 26 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 core_a_data_rdata_i[21]
port 27 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 core_a_data_rdata_i[22]
port 28 nsew signal input
rlabel metal2 s 28538 29200 28594 30000 6 core_a_data_rdata_i[23]
port 29 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 core_a_data_rdata_i[24]
port 30 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 core_a_data_rdata_i[25]
port 31 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 core_a_data_rdata_i[26]
port 32 nsew signal input
rlabel metal2 s 31758 29200 31814 30000 6 core_a_data_rdata_i[27]
port 33 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 core_a_data_rdata_i[28]
port 34 nsew signal input
rlabel metal2 s 41418 29200 41474 30000 6 core_a_data_rdata_i[29]
port 35 nsew signal input
rlabel metal2 s 11978 29200 12034 30000 6 core_a_data_rdata_i[2]
port 36 nsew signal input
rlabel metal2 s 38658 29200 38714 30000 6 core_a_data_rdata_i[30]
port 37 nsew signal input
rlabel metal2 s 26698 29200 26754 30000 6 core_a_data_rdata_i[31]
port 38 nsew signal input
rlabel metal2 s 15658 29200 15714 30000 6 core_a_data_rdata_i[3]
port 39 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 core_a_data_rdata_i[4]
port 40 nsew signal input
rlabel metal3 s 59200 14288 60000 14408 6 core_a_data_rdata_i[5]
port 41 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 core_a_data_rdata_i[6]
port 42 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 core_a_data_rdata_i[7]
port 43 nsew signal input
rlabel metal2 s 45098 29200 45154 30000 6 core_a_data_rdata_i[8]
port 44 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 core_a_data_rdata_i[9]
port 45 nsew signal input
rlabel metal2 s 24398 29200 24454 30000 6 core_a_data_req_o
port 46 nsew signal tristate
rlabel metal2 s 11978 0 12034 800 6 core_a_data_rvalid_i
port 47 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 core_a_data_wdata_o[0]
port 48 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 core_a_data_wdata_o[10]
port 49 nsew signal tristate
rlabel metal2 s 54298 0 54354 800 6 core_a_data_wdata_o[11]
port 50 nsew signal tristate
rlabel metal2 s 35438 29200 35494 30000 6 core_a_data_wdata_o[12]
port 51 nsew signal tristate
rlabel metal2 s 9678 29200 9734 30000 6 core_a_data_wdata_o[13]
port 52 nsew signal tristate
rlabel metal2 s 12438 29200 12494 30000 6 core_a_data_wdata_o[14]
port 53 nsew signal tristate
rlabel metal2 s 43258 29200 43314 30000 6 core_a_data_wdata_o[15]
port 54 nsew signal tristate
rlabel metal2 s 46478 29200 46534 30000 6 core_a_data_wdata_o[16]
port 55 nsew signal tristate
rlabel metal3 s 59200 16328 60000 16448 6 core_a_data_wdata_o[17]
port 56 nsew signal tristate
rlabel metal2 s 19338 29200 19394 30000 6 core_a_data_wdata_o[18]
port 57 nsew signal tristate
rlabel metal2 s 31298 0 31354 800 6 core_a_data_wdata_o[19]
port 58 nsew signal tristate
rlabel metal2 s 54758 29200 54814 30000 6 core_a_data_wdata_o[1]
port 59 nsew signal tristate
rlabel metal2 s 37278 0 37334 800 6 core_a_data_wdata_o[20]
port 60 nsew signal tristate
rlabel metal2 s 57518 29200 57574 30000 6 core_a_data_wdata_o[21]
port 61 nsew signal tristate
rlabel metal2 s 3238 29200 3294 30000 6 core_a_data_wdata_o[22]
port 62 nsew signal tristate
rlabel metal2 s 23938 0 23994 800 6 core_a_data_wdata_o[23]
port 63 nsew signal tristate
rlabel metal3 s 59200 10208 60000 10328 6 core_a_data_wdata_o[24]
port 64 nsew signal tristate
rlabel metal2 s 21638 0 21694 800 6 core_a_data_wdata_o[25]
port 65 nsew signal tristate
rlabel metal2 s 23478 0 23534 800 6 core_a_data_wdata_o[26]
port 66 nsew signal tristate
rlabel metal3 s 59200 19728 60000 19848 6 core_a_data_wdata_o[27]
port 67 nsew signal tristate
rlabel metal2 s 25778 29200 25834 30000 6 core_a_data_wdata_o[28]
port 68 nsew signal tristate
rlabel metal2 s 37278 29200 37334 30000 6 core_a_data_wdata_o[29]
port 69 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 core_a_data_wdata_o[2]
port 70 nsew signal tristate
rlabel metal2 s 35438 0 35494 800 6 core_a_data_wdata_o[30]
port 71 nsew signal tristate
rlabel metal2 s 45558 29200 45614 30000 6 core_a_data_wdata_o[31]
port 72 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 core_a_data_wdata_o[3]
port 73 nsew signal tristate
rlabel metal3 s 0 25848 800 25968 6 core_a_data_wdata_o[4]
port 74 nsew signal tristate
rlabel metal2 s 25778 0 25834 800 6 core_a_data_wdata_o[5]
port 75 nsew signal tristate
rlabel metal2 s 20258 0 20314 800 6 core_a_data_wdata_o[6]
port 76 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 core_a_data_wdata_o[7]
port 77 nsew signal tristate
rlabel metal2 s 48778 29200 48834 30000 6 core_a_data_wdata_o[8]
port 78 nsew signal tristate
rlabel metal2 s 17958 29200 18014 30000 6 core_a_data_wdata_o[9]
port 79 nsew signal tristate
rlabel metal3 s 59200 8168 60000 8288 6 core_a_data_we_o
port 80 nsew signal tristate
rlabel metal2 s 2318 0 2374 800 6 core_b_data_addr_o[0]
port 81 nsew signal tristate
rlabel metal2 s 32218 29200 32274 30000 6 core_b_data_addr_o[1]
port 82 nsew signal tristate
rlabel metal2 s 2778 29200 2834 30000 6 core_b_data_addr_o[2]
port 83 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 core_b_data_addr_o[3]
port 84 nsew signal tristate
rlabel metal2 s 56138 29200 56194 30000 6 core_b_data_addr_o[4]
port 85 nsew signal tristate
rlabel metal2 s 36818 29200 36874 30000 6 core_b_data_addr_o[5]
port 86 nsew signal tristate
rlabel metal2 s 7838 0 7894 800 6 core_b_data_addr_o[6]
port 87 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 core_b_data_addr_o[7]
port 88 nsew signal tristate
rlabel metal2 s 58898 0 58954 800 6 core_b_data_addr_o[8]
port 89 nsew signal tristate
rlabel metal2 s 57518 0 57574 800 6 core_b_data_addr_o[9]
port 90 nsew signal tristate
rlabel metal2 s 25318 0 25374 800 6 core_b_data_be_o[0]
port 91 nsew signal tristate
rlabel metal2 s 18878 0 18934 800 6 core_b_data_be_o[1]
port 92 nsew signal tristate
rlabel metal2 s 5538 29200 5594 30000 6 core_b_data_be_o[2]
port 93 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 core_b_data_be_o[3]
port 94 nsew signal tristate
rlabel metal2 s 49698 0 49754 800 6 core_b_data_rdata_i[0]
port 95 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 core_b_data_rdata_i[10]
port 96 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 core_b_data_rdata_i[11]
port 97 nsew signal input
rlabel metal2 s 17038 29200 17094 30000 6 core_b_data_rdata_i[12]
port 98 nsew signal input
rlabel metal2 s 53378 29200 53434 30000 6 core_b_data_rdata_i[13]
port 99 nsew signal input
rlabel metal2 s 33598 29200 33654 30000 6 core_b_data_rdata_i[14]
port 100 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 core_b_data_rdata_i[15]
port 101 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 core_b_data_rdata_i[16]
port 102 nsew signal input
rlabel metal3 s 59200 25848 60000 25968 6 core_b_data_rdata_i[17]
port 103 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 core_b_data_rdata_i[18]
port 104 nsew signal input
rlabel metal2 s 40038 29200 40094 30000 6 core_b_data_rdata_i[19]
port 105 nsew signal input
rlabel metal2 s 938 29200 994 30000 6 core_b_data_rdata_i[1]
port 106 nsew signal input
rlabel metal3 s 59200 2048 60000 2168 6 core_b_data_rdata_i[20]
port 107 nsew signal input
rlabel metal3 s 59200 4088 60000 4208 6 core_b_data_rdata_i[21]
port 108 nsew signal input
rlabel metal2 s 36358 29200 36414 30000 6 core_b_data_rdata_i[22]
port 109 nsew signal input
rlabel metal3 s 59200 17688 60000 17808 6 core_b_data_rdata_i[23]
port 110 nsew signal input
rlabel metal2 s 12898 29200 12954 30000 6 core_b_data_rdata_i[24]
port 111 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 core_b_data_rdata_i[25]
port 112 nsew signal input
rlabel metal2 s 46938 29200 46994 30000 6 core_b_data_rdata_i[26]
port 113 nsew signal input
rlabel metal2 s 4618 29200 4674 30000 6 core_b_data_rdata_i[27]
port 114 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 core_b_data_rdata_i[28]
port 115 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 core_b_data_rdata_i[29]
port 116 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 core_b_data_rdata_i[2]
port 117 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 core_b_data_rdata_i[30]
port 118 nsew signal input
rlabel metal2 s 11058 29200 11114 30000 6 core_b_data_rdata_i[31]
port 119 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 core_b_data_rdata_i[3]
port 120 nsew signal input
rlabel metal2 s 48318 29200 48374 30000 6 core_b_data_rdata_i[4]
port 121 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 core_b_data_rdata_i[5]
port 122 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 core_b_data_rdata_i[6]
port 123 nsew signal input
rlabel metal3 s 59200 4768 60000 4888 6 core_b_data_rdata_i[7]
port 124 nsew signal input
rlabel metal2 s 34058 29200 34114 30000 6 core_b_data_rdata_i[8]
port 125 nsew signal input
rlabel metal3 s 59200 21088 60000 21208 6 core_b_data_rdata_i[9]
port 126 nsew signal input
rlabel metal2 s 52918 29200 52974 30000 6 core_b_data_req_o
port 127 nsew signal tristate
rlabel metal2 s 51538 29200 51594 30000 6 core_b_data_rvalid_i
port 128 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 core_b_data_wdata_o[0]
port 129 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 core_b_data_wdata_o[10]
port 130 nsew signal tristate
rlabel metal2 s 48318 0 48374 800 6 core_b_data_wdata_o[11]
port 131 nsew signal tristate
rlabel metal2 s 56598 0 56654 800 6 core_b_data_wdata_o[12]
port 132 nsew signal tristate
rlabel metal2 s 50158 29200 50214 30000 6 core_b_data_wdata_o[13]
port 133 nsew signal tristate
rlabel metal2 s 41878 0 41934 800 6 core_b_data_wdata_o[14]
port 134 nsew signal tristate
rlabel metal2 s 39578 0 39634 800 6 core_b_data_wdata_o[15]
port 135 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 core_b_data_wdata_o[16]
port 136 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 core_b_data_wdata_o[17]
port 137 nsew signal tristate
rlabel metal2 s 20718 29200 20774 30000 6 core_b_data_wdata_o[18]
port 138 nsew signal tristate
rlabel metal2 s 30838 29200 30894 30000 6 core_b_data_wdata_o[19]
port 139 nsew signal tristate
rlabel metal2 s 5998 29200 6054 30000 6 core_b_data_wdata_o[1]
port 140 nsew signal tristate
rlabel metal2 s 27618 29200 27674 30000 6 core_b_data_wdata_o[20]
port 141 nsew signal tristate
rlabel metal2 s 31758 0 31814 800 6 core_b_data_wdata_o[21]
port 142 nsew signal tristate
rlabel metal2 s 26698 0 26754 800 6 core_b_data_wdata_o[22]
port 143 nsew signal tristate
rlabel metal2 s 28998 29200 29054 30000 6 core_b_data_wdata_o[23]
port 144 nsew signal tristate
rlabel metal2 s 22558 29200 22614 30000 6 core_b_data_wdata_o[24]
port 145 nsew signal tristate
rlabel metal3 s 0 22448 800 22568 6 core_b_data_wdata_o[25]
port 146 nsew signal tristate
rlabel metal2 s 36358 0 36414 800 6 core_b_data_wdata_o[26]
port 147 nsew signal tristate
rlabel metal3 s 59200 21768 60000 21888 6 core_b_data_wdata_o[27]
port 148 nsew signal tristate
rlabel metal3 s 59200 28568 60000 28688 6 core_b_data_wdata_o[28]
port 149 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 core_b_data_wdata_o[29]
port 150 nsew signal tristate
rlabel metal2 s 49698 29200 49754 30000 6 core_b_data_wdata_o[2]
port 151 nsew signal tristate
rlabel metal2 s 42798 29200 42854 30000 6 core_b_data_wdata_o[30]
port 152 nsew signal tristate
rlabel metal2 s 28538 0 28594 800 6 core_b_data_wdata_o[31]
port 153 nsew signal tristate
rlabel metal2 s 56598 29200 56654 30000 6 core_b_data_wdata_o[3]
port 154 nsew signal tristate
rlabel metal2 s 16118 29200 16174 30000 6 core_b_data_wdata_o[4]
port 155 nsew signal tristate
rlabel metal2 s 51078 0 51134 800 6 core_b_data_wdata_o[5]
port 156 nsew signal tristate
rlabel metal2 s 44638 29200 44694 30000 6 core_b_data_wdata_o[6]
port 157 nsew signal tristate
rlabel metal2 s 27158 29200 27214 30000 6 core_b_data_wdata_o[7]
port 158 nsew signal tristate
rlabel metal2 s 6458 29200 6514 30000 6 core_b_data_wdata_o[8]
port 159 nsew signal tristate
rlabel metal3 s 0 25168 800 25288 6 core_b_data_wdata_o[9]
port 160 nsew signal tristate
rlabel metal2 s 51078 29200 51134 30000 6 core_b_data_we_o
port 161 nsew signal tristate
rlabel metal3 s 59200 12248 60000 12368 6 wb_data_addr_i[0]
port 162 nsew signal input
rlabel metal2 s 938 0 994 800 6 wb_data_addr_i[10]
port 163 nsew signal input
rlabel metal2 s 2318 29200 2374 30000 6 wb_data_addr_i[1]
port 164 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 wb_data_addr_i[2]
port 165 nsew signal input
rlabel metal3 s 59200 14968 60000 15088 6 wb_data_addr_i[3]
port 166 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wb_data_addr_i[4]
port 167 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wb_data_addr_i[5]
port 168 nsew signal input
rlabel metal2 s 7378 29200 7434 30000 6 wb_data_addr_i[6]
port 169 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wb_data_addr_i[7]
port 170 nsew signal input
rlabel metal2 s 7838 29200 7894 30000 6 wb_data_addr_i[8]
port 171 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wb_data_addr_i[9]
port 172 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wb_data_be_i[0]
port 173 nsew signal input
rlabel metal2 s 8758 29200 8814 30000 6 wb_data_be_i[1]
port 174 nsew signal input
rlabel metal2 s 17498 29200 17554 30000 6 wb_data_be_i[2]
port 175 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wb_data_be_i[3]
port 176 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wb_data_rdata_o[0]
port 177 nsew signal tristate
rlabel metal2 s 14738 29200 14794 30000 6 wb_data_rdata_o[10]
port 178 nsew signal tristate
rlabel metal3 s 59200 11568 60000 11688 6 wb_data_rdata_o[11]
port 179 nsew signal tristate
rlabel metal2 s 58438 29200 58494 30000 6 wb_data_rdata_o[12]
port 180 nsew signal tristate
rlabel metal2 s 40038 0 40094 800 6 wb_data_rdata_o[13]
port 181 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 wb_data_rdata_o[14]
port 182 nsew signal tristate
rlabel metal2 s 24858 0 24914 800 6 wb_data_rdata_o[15]
port 183 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 wb_data_rdata_o[16]
port 184 nsew signal tristate
rlabel metal2 s 39578 29200 39634 30000 6 wb_data_rdata_o[17]
port 185 nsew signal tristate
rlabel metal2 s 20258 29200 20314 30000 6 wb_data_rdata_o[18]
port 186 nsew signal tristate
rlabel metal2 s 51538 0 51594 800 6 wb_data_rdata_o[19]
port 187 nsew signal tristate
rlabel metal3 s 59200 5448 60000 5568 6 wb_data_rdata_o[1]
port 188 nsew signal tristate
rlabel metal2 s 41878 29200 41934 30000 6 wb_data_rdata_o[20]
port 189 nsew signal tristate
rlabel metal2 s 46478 0 46534 800 6 wb_data_rdata_o[21]
port 190 nsew signal tristate
rlabel metal2 s 1398 29200 1454 30000 6 wb_data_rdata_o[22]
port 191 nsew signal tristate
rlabel metal2 s 54758 0 54814 800 6 wb_data_rdata_o[23]
port 192 nsew signal tristate
rlabel metal2 s 21178 29200 21234 30000 6 wb_data_rdata_o[24]
port 193 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 wb_data_rdata_o[25]
port 194 nsew signal tristate
rlabel metal2 s 9218 29200 9274 30000 6 wb_data_rdata_o[26]
port 195 nsew signal tristate
rlabel metal2 s 478 0 534 800 6 wb_data_rdata_o[27]
port 196 nsew signal tristate
rlabel metal2 s 4158 29200 4214 30000 6 wb_data_rdata_o[28]
port 197 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 wb_data_rdata_o[29]
port 198 nsew signal tristate
rlabel metal2 s 33138 29200 33194 30000 6 wb_data_rdata_o[2]
port 199 nsew signal tristate
rlabel metal3 s 0 28568 800 28688 6 wb_data_rdata_o[30]
port 200 nsew signal tristate
rlabel metal2 s 11058 0 11114 800 6 wb_data_rdata_o[31]
port 201 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 wb_data_rdata_o[3]
port 202 nsew signal tristate
rlabel metal2 s 4618 0 4674 800 6 wb_data_rdata_o[4]
port 203 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 wb_data_rdata_o[5]
port 204 nsew signal tristate
rlabel metal2 s 50158 0 50214 800 6 wb_data_rdata_o[6]
port 205 nsew signal tristate
rlabel metal2 s 27158 0 27214 800 6 wb_data_rdata_o[7]
port 206 nsew signal tristate
rlabel metal2 s 30378 0 30434 800 6 wb_data_rdata_o[8]
port 207 nsew signal tristate
rlabel metal2 s 47858 29200 47914 30000 6 wb_data_rdata_o[9]
port 208 nsew signal tristate
rlabel metal2 s 44638 0 44694 800 6 wb_data_rvalid_o
port 209 nsew signal tristate
rlabel metal3 s 59200 17008 60000 17128 6 wb_data_wdata_i[0]
port 210 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 wb_data_wdata_i[10]
port 211 nsew signal input
rlabel metal3 s 59200 7488 60000 7608 6 wb_data_wdata_i[11]
port 212 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wb_data_wdata_i[12]
port 213 nsew signal input
rlabel metal2 s 14278 29200 14334 30000 6 wb_data_wdata_i[13]
port 214 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wb_data_wdata_i[14]
port 215 nsew signal input
rlabel metal3 s 59200 688 60000 808 6 wb_data_wdata_i[15]
port 216 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wb_data_wdata_i[16]
port 217 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 wb_data_wdata_i[17]
port 218 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_data_wdata_i[18]
port 219 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wb_data_wdata_i[19]
port 220 nsew signal input
rlabel metal3 s 59200 23808 60000 23928 6 wb_data_wdata_i[1]
port 221 nsew signal input
rlabel metal2 s 25318 29200 25374 30000 6 wb_data_wdata_i[20]
port 222 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 wb_data_wdata_i[21]
port 223 nsew signal input
rlabel metal2 s 23478 29200 23534 30000 6 wb_data_wdata_i[22]
port 224 nsew signal input
rlabel metal2 s 34978 29200 35034 30000 6 wb_data_wdata_i[23]
port 225 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wb_data_wdata_i[24]
port 226 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 wb_data_wdata_i[25]
port 227 nsew signal input
rlabel metal2 s 40498 29200 40554 30000 6 wb_data_wdata_i[26]
port 228 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wb_data_wdata_i[27]
port 229 nsew signal input
rlabel metal3 s 59200 12928 60000 13048 6 wb_data_wdata_i[28]
port 230 nsew signal input
rlabel metal2 s 22098 29200 22154 30000 6 wb_data_wdata_i[29]
port 231 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wb_data_wdata_i[2]
port 232 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wb_data_wdata_i[30]
port 233 nsew signal input
rlabel metal3 s 59200 24488 60000 24608 6 wb_data_wdata_i[31]
port 234 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 wb_data_wdata_i[3]
port 235 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wb_data_wdata_i[4]
port 236 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 wb_data_wdata_i[5]
port 237 nsew signal input
rlabel metal3 s 59200 6808 60000 6928 6 wb_data_wdata_i[6]
port 238 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wb_data_wdata_i[7]
port 239 nsew signal input
rlabel metal2 s 30378 29200 30434 30000 6 wb_data_wdata_i[8]
port 240 nsew signal input
rlabel metal2 s 38198 29200 38254 30000 6 wb_data_wdata_i[9]
port 241 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 wb_data_we_i
port 242 nsew signal input
rlabel metal2 s 18878 29200 18934 30000 6 wbs_cyc_i
port 243 nsew signal input
rlabel metal2 s 59358 29200 59414 30000 6 wbs_stb_i
port 244 nsew signal input
rlabel metal4 s 49104 2128 49424 27792 6 VPWR
port 245 nsew power bidirectional
rlabel metal4 s 29840 2128 30160 27792 6 VPWR
port 246 nsew power bidirectional
rlabel metal4 s 10576 2128 10896 27792 6 VPWR
port 247 nsew power bidirectional
rlabel metal5 s 1104 23341 58880 23661 6 VPWR
port 248 nsew power bidirectional
rlabel metal5 s 1104 14792 58880 15112 6 VPWR
port 249 nsew power bidirectional
rlabel metal5 s 1104 6243 58880 6563 6 VPWR
port 250 nsew power bidirectional
rlabel metal4 s 39472 2128 39792 27792 6 VGND
port 251 nsew ground bidirectional
rlabel metal4 s 20208 2128 20528 27792 6 VGND
port 252 nsew ground bidirectional
rlabel metal5 s 1104 19067 58880 19387 6 VGND
port 253 nsew ground bidirectional
rlabel metal5 s 1104 10517 58880 10837 6 VGND
port 254 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 30000
<< end >>
