magic
tech sky130A
magscale 1 2
timestamp 1624394029
<< obsli1 >>
rect 1104 2159 238832 239921
<< obsm1 >>
rect 474 1708 239278 240304
<< metal2 >>
rect 2318 241292 2374 242092
rect 5078 241292 5134 242092
rect 7838 241292 7894 242092
rect 10598 241292 10654 242092
rect 13358 241292 13414 242092
rect 16118 241292 16174 242092
rect 18878 241292 18934 242092
rect 21638 241292 21694 242092
rect 24398 241292 24454 242092
rect 27158 241292 27214 242092
rect 29918 241292 29974 242092
rect 32678 241292 32734 242092
rect 35438 241292 35494 242092
rect 38198 241292 38254 242092
rect 41418 241292 41474 242092
rect 44178 241292 44234 242092
rect 46938 241292 46994 242092
rect 49698 241292 49754 242092
rect 52458 241292 52514 242092
rect 55218 241292 55274 242092
rect 57978 241292 58034 242092
rect 60738 241292 60794 242092
rect 63498 241292 63554 242092
rect 66258 241292 66314 242092
rect 69018 241292 69074 242092
rect 71778 241292 71834 242092
rect 74538 241292 74594 242092
rect 77298 241292 77354 242092
rect 80518 241292 80574 242092
rect 83278 241292 83334 242092
rect 86038 241292 86094 242092
rect 88798 241292 88854 242092
rect 91558 241292 91614 242092
rect 94318 241292 94374 242092
rect 97078 241292 97134 242092
rect 99838 241292 99894 242092
rect 102598 241292 102654 242092
rect 105358 241292 105414 242092
rect 108118 241292 108174 242092
rect 110878 241292 110934 242092
rect 113638 241292 113694 242092
rect 116398 241292 116454 242092
rect 119618 241292 119674 242092
rect 122378 241292 122434 242092
rect 125138 241292 125194 242092
rect 127898 241292 127954 242092
rect 130658 241292 130714 242092
rect 133418 241292 133474 242092
rect 136178 241292 136234 242092
rect 138938 241292 138994 242092
rect 141698 241292 141754 242092
rect 144458 241292 144514 242092
rect 147218 241292 147274 242092
rect 149978 241292 150034 242092
rect 152738 241292 152794 242092
rect 155498 241292 155554 242092
rect 158258 241292 158314 242092
rect 161478 241292 161534 242092
rect 164238 241292 164294 242092
rect 166998 241292 167054 242092
rect 169758 241292 169814 242092
rect 172518 241292 172574 242092
rect 175278 241292 175334 242092
rect 178038 241292 178094 242092
rect 180798 241292 180854 242092
rect 183558 241292 183614 242092
rect 186318 241292 186374 242092
rect 189078 241292 189134 242092
rect 191838 241292 191894 242092
rect 194598 241292 194654 242092
rect 197358 241292 197414 242092
rect 200578 241292 200634 242092
rect 203338 241292 203394 242092
rect 206098 241292 206154 242092
rect 208858 241292 208914 242092
rect 211618 241292 211674 242092
rect 214378 241292 214434 242092
rect 217138 241292 217194 242092
rect 219898 241292 219954 242092
rect 222658 241292 222714 242092
rect 225418 241292 225474 242092
rect 228178 241292 228234 242092
rect 230938 241292 230994 242092
rect 233698 241292 233754 242092
rect 236458 241292 236514 242092
rect 239218 241292 239274 242092
rect 478 0 534 800
rect 3238 0 3294 800
rect 5998 0 6054 800
rect 8758 0 8814 800
rect 11518 0 11574 800
rect 14278 0 14334 800
rect 17038 0 17094 800
rect 19798 0 19854 800
rect 22558 0 22614 800
rect 25318 0 25374 800
rect 28078 0 28134 800
rect 30838 0 30894 800
rect 33598 0 33654 800
rect 36358 0 36414 800
rect 39118 0 39174 800
rect 42338 0 42394 800
rect 45098 0 45154 800
rect 47858 0 47914 800
rect 50618 0 50674 800
rect 53378 0 53434 800
rect 56138 0 56194 800
rect 58898 0 58954 800
rect 61658 0 61714 800
rect 64418 0 64474 800
rect 67178 0 67234 800
rect 69938 0 69994 800
rect 72698 0 72754 800
rect 75458 0 75514 800
rect 78218 0 78274 800
rect 81438 0 81494 800
rect 84198 0 84254 800
rect 86958 0 87014 800
rect 89718 0 89774 800
rect 92478 0 92534 800
rect 95238 0 95294 800
rect 97998 0 98054 800
rect 100758 0 100814 800
rect 103518 0 103574 800
rect 106278 0 106334 800
rect 109038 0 109094 800
rect 111798 0 111854 800
rect 114558 0 114614 800
rect 117318 0 117374 800
rect 120078 0 120134 800
rect 123298 0 123354 800
rect 126058 0 126114 800
rect 128818 0 128874 800
rect 131578 0 131634 800
rect 134338 0 134394 800
rect 137098 0 137154 800
rect 139858 0 139914 800
rect 142618 0 142674 800
rect 145378 0 145434 800
rect 148138 0 148194 800
rect 150898 0 150954 800
rect 153658 0 153714 800
rect 156418 0 156474 800
rect 159178 0 159234 800
rect 162398 0 162454 800
rect 165158 0 165214 800
rect 167918 0 167974 800
rect 170678 0 170734 800
rect 173438 0 173494 800
rect 176198 0 176254 800
rect 178958 0 179014 800
rect 181718 0 181774 800
rect 184478 0 184534 800
rect 187238 0 187294 800
rect 189998 0 190054 800
rect 192758 0 192814 800
rect 195518 0 195574 800
rect 198278 0 198334 800
rect 201498 0 201554 800
rect 204258 0 204314 800
rect 207018 0 207074 800
rect 209778 0 209834 800
rect 212538 0 212594 800
rect 215298 0 215354 800
rect 218058 0 218114 800
rect 220818 0 220874 800
rect 223578 0 223634 800
rect 226338 0 226394 800
rect 229098 0 229154 800
rect 231858 0 231914 800
rect 234618 0 234674 800
rect 237378 0 237434 800
<< obsm2 >>
rect 480 241236 2262 241292
rect 2430 241236 5022 241292
rect 5190 241236 7782 241292
rect 7950 241236 10542 241292
rect 10710 241236 13302 241292
rect 13470 241236 16062 241292
rect 16230 241236 18822 241292
rect 18990 241236 21582 241292
rect 21750 241236 24342 241292
rect 24510 241236 27102 241292
rect 27270 241236 29862 241292
rect 30030 241236 32622 241292
rect 32790 241236 35382 241292
rect 35550 241236 38142 241292
rect 38310 241236 41362 241292
rect 41530 241236 44122 241292
rect 44290 241236 46882 241292
rect 47050 241236 49642 241292
rect 49810 241236 52402 241292
rect 52570 241236 55162 241292
rect 55330 241236 57922 241292
rect 58090 241236 60682 241292
rect 60850 241236 63442 241292
rect 63610 241236 66202 241292
rect 66370 241236 68962 241292
rect 69130 241236 71722 241292
rect 71890 241236 74482 241292
rect 74650 241236 77242 241292
rect 77410 241236 80462 241292
rect 80630 241236 83222 241292
rect 83390 241236 85982 241292
rect 86150 241236 88742 241292
rect 88910 241236 91502 241292
rect 91670 241236 94262 241292
rect 94430 241236 97022 241292
rect 97190 241236 99782 241292
rect 99950 241236 102542 241292
rect 102710 241236 105302 241292
rect 105470 241236 108062 241292
rect 108230 241236 110822 241292
rect 110990 241236 113582 241292
rect 113750 241236 116342 241292
rect 116510 241236 119562 241292
rect 119730 241236 122322 241292
rect 122490 241236 125082 241292
rect 125250 241236 127842 241292
rect 128010 241236 130602 241292
rect 130770 241236 133362 241292
rect 133530 241236 136122 241292
rect 136290 241236 138882 241292
rect 139050 241236 141642 241292
rect 141810 241236 144402 241292
rect 144570 241236 147162 241292
rect 147330 241236 149922 241292
rect 150090 241236 152682 241292
rect 152850 241236 155442 241292
rect 155610 241236 158202 241292
rect 158370 241236 161422 241292
rect 161590 241236 164182 241292
rect 164350 241236 166942 241292
rect 167110 241236 169702 241292
rect 169870 241236 172462 241292
rect 172630 241236 175222 241292
rect 175390 241236 177982 241292
rect 178150 241236 180742 241292
rect 180910 241236 183502 241292
rect 183670 241236 186262 241292
rect 186430 241236 189022 241292
rect 189190 241236 191782 241292
rect 191950 241236 194542 241292
rect 194710 241236 197302 241292
rect 197470 241236 200522 241292
rect 200690 241236 203282 241292
rect 203450 241236 206042 241292
rect 206210 241236 208802 241292
rect 208970 241236 211562 241292
rect 211730 241236 214322 241292
rect 214490 241236 217082 241292
rect 217250 241236 219842 241292
rect 220010 241236 222602 241292
rect 222770 241236 225362 241292
rect 225530 241236 228122 241292
rect 228290 241236 230882 241292
rect 231050 241236 233642 241292
rect 233810 241236 236402 241292
rect 236570 241236 239162 241292
rect 480 856 239272 241236
rect 590 800 3182 856
rect 3350 800 5942 856
rect 6110 800 8702 856
rect 8870 800 11462 856
rect 11630 800 14222 856
rect 14390 800 16982 856
rect 17150 800 19742 856
rect 19910 800 22502 856
rect 22670 800 25262 856
rect 25430 800 28022 856
rect 28190 800 30782 856
rect 30950 800 33542 856
rect 33710 800 36302 856
rect 36470 800 39062 856
rect 39230 800 42282 856
rect 42450 800 45042 856
rect 45210 800 47802 856
rect 47970 800 50562 856
rect 50730 800 53322 856
rect 53490 800 56082 856
rect 56250 800 58842 856
rect 59010 800 61602 856
rect 61770 800 64362 856
rect 64530 800 67122 856
rect 67290 800 69882 856
rect 70050 800 72642 856
rect 72810 800 75402 856
rect 75570 800 78162 856
rect 78330 800 81382 856
rect 81550 800 84142 856
rect 84310 800 86902 856
rect 87070 800 89662 856
rect 89830 800 92422 856
rect 92590 800 95182 856
rect 95350 800 97942 856
rect 98110 800 100702 856
rect 100870 800 103462 856
rect 103630 800 106222 856
rect 106390 800 108982 856
rect 109150 800 111742 856
rect 111910 800 114502 856
rect 114670 800 117262 856
rect 117430 800 120022 856
rect 120190 800 123242 856
rect 123410 800 126002 856
rect 126170 800 128762 856
rect 128930 800 131522 856
rect 131690 800 134282 856
rect 134450 800 137042 856
rect 137210 800 139802 856
rect 139970 800 142562 856
rect 142730 800 145322 856
rect 145490 800 148082 856
rect 148250 800 150842 856
rect 151010 800 153602 856
rect 153770 800 156362 856
rect 156530 800 159122 856
rect 159290 800 162342 856
rect 162510 800 165102 856
rect 165270 800 167862 856
rect 168030 800 170622 856
rect 170790 800 173382 856
rect 173550 800 176142 856
rect 176310 800 178902 856
rect 179070 800 181662 856
rect 181830 800 184422 856
rect 184590 800 187182 856
rect 187350 800 189942 856
rect 190110 800 192702 856
rect 192870 800 195462 856
rect 195630 800 198222 856
rect 198390 800 201442 856
rect 201610 800 204202 856
rect 204370 800 206962 856
rect 207130 800 209722 856
rect 209890 800 212482 856
rect 212650 800 215242 856
rect 215410 800 218002 856
rect 218170 800 220762 856
rect 220930 800 223522 856
rect 223690 800 226282 856
rect 226450 800 229042 856
rect 229210 800 231802 856
rect 231970 800 234562 856
rect 234730 800 237322 856
rect 237490 800 239272 856
<< metal3 >>
rect 0 240048 800 240168
rect 239148 236648 239948 236768
rect 0 235288 800 235408
rect 239148 232568 239948 232688
rect 0 231208 800 231328
rect 239148 228488 239948 228608
rect 0 227128 800 227248
rect 239148 224408 239948 224528
rect 0 223048 800 223168
rect 239148 220328 239948 220448
rect 0 218968 800 219088
rect 239148 216248 239948 216368
rect 0 214888 800 215008
rect 239148 212168 239948 212288
rect 0 210808 800 210928
rect 239148 208088 239948 208208
rect 0 206728 800 206848
rect 239148 204008 239948 204128
rect 0 202648 800 202768
rect 239148 199928 239948 200048
rect 0 198568 800 198688
rect 239148 195848 239948 195968
rect 0 194488 800 194608
rect 239148 191768 239948 191888
rect 0 190408 800 190528
rect 239148 187688 239948 187808
rect 0 186328 800 186448
rect 239148 183608 239948 183728
rect 0 182248 800 182368
rect 239148 178848 239948 178968
rect 0 177488 800 177608
rect 239148 174768 239948 174888
rect 0 173408 800 173528
rect 239148 170688 239948 170808
rect 0 169328 800 169448
rect 239148 166608 239948 166728
rect 0 165248 800 165368
rect 239148 162528 239948 162648
rect 0 161168 800 161288
rect 239148 158448 239948 158568
rect 0 157088 800 157208
rect 239148 154368 239948 154488
rect 0 153008 800 153128
rect 239148 150288 239948 150408
rect 0 148928 800 149048
rect 239148 146208 239948 146328
rect 0 144848 800 144968
rect 239148 142128 239948 142248
rect 0 140768 800 140888
rect 239148 138048 239948 138168
rect 0 136688 800 136808
rect 239148 133968 239948 134088
rect 0 132608 800 132728
rect 239148 129888 239948 130008
rect 0 128528 800 128648
rect 239148 125808 239948 125928
rect 0 124448 800 124568
rect 239148 121048 239948 121168
rect 0 120368 800 120488
rect 239148 116968 239948 117088
rect 0 115608 800 115728
rect 239148 112888 239948 113008
rect 0 111528 800 111648
rect 239148 108808 239948 108928
rect 0 107448 800 107568
rect 239148 104728 239948 104848
rect 0 103368 800 103488
rect 239148 100648 239948 100768
rect 0 99288 800 99408
rect 239148 96568 239948 96688
rect 0 95208 800 95328
rect 239148 92488 239948 92608
rect 0 91128 800 91248
rect 239148 88408 239948 88528
rect 0 87048 800 87168
rect 239148 84328 239948 84448
rect 0 82968 800 83088
rect 239148 80248 239948 80368
rect 0 78888 800 79008
rect 239148 76168 239948 76288
rect 0 74808 800 74928
rect 239148 72088 239948 72208
rect 0 70728 800 70848
rect 239148 68008 239948 68128
rect 0 66648 800 66768
rect 239148 63928 239948 64048
rect 0 62568 800 62688
rect 239148 59168 239948 59288
rect 0 57808 800 57928
rect 239148 55088 239948 55208
rect 0 53728 800 53848
rect 239148 51008 239948 51128
rect 0 49648 800 49768
rect 239148 46928 239948 47048
rect 0 45568 800 45688
rect 239148 42848 239948 42968
rect 0 41488 800 41608
rect 239148 38768 239948 38888
rect 0 37408 800 37528
rect 239148 34688 239948 34808
rect 0 33328 800 33448
rect 239148 30608 239948 30728
rect 0 29248 800 29368
rect 239148 26528 239948 26648
rect 0 25168 800 25288
rect 239148 22448 239948 22568
rect 0 21088 800 21208
rect 239148 18368 239948 18488
rect 0 17008 800 17128
rect 239148 14288 239948 14408
rect 0 12928 800 13048
rect 239148 10208 239948 10328
rect 0 8848 800 8968
rect 239148 6128 239948 6248
rect 0 4768 800 4888
rect 239148 1368 239948 1488
<< obsm3 >>
rect 800 240248 239148 240549
rect 880 239968 239148 240248
rect 800 236848 239148 239968
rect 800 236568 239068 236848
rect 800 235488 239148 236568
rect 880 235208 239148 235488
rect 800 232768 239148 235208
rect 800 232488 239068 232768
rect 800 231408 239148 232488
rect 880 231128 239148 231408
rect 800 228688 239148 231128
rect 800 228408 239068 228688
rect 800 227328 239148 228408
rect 880 227048 239148 227328
rect 800 224608 239148 227048
rect 800 224328 239068 224608
rect 800 223248 239148 224328
rect 880 222968 239148 223248
rect 800 220528 239148 222968
rect 800 220248 239068 220528
rect 800 219168 239148 220248
rect 880 218888 239148 219168
rect 800 216448 239148 218888
rect 800 216168 239068 216448
rect 800 215088 239148 216168
rect 880 214808 239148 215088
rect 800 212368 239148 214808
rect 800 212088 239068 212368
rect 800 211008 239148 212088
rect 880 210728 239148 211008
rect 800 208288 239148 210728
rect 800 208008 239068 208288
rect 800 206928 239148 208008
rect 880 206648 239148 206928
rect 800 204208 239148 206648
rect 800 203928 239068 204208
rect 800 202848 239148 203928
rect 880 202568 239148 202848
rect 800 200128 239148 202568
rect 800 199848 239068 200128
rect 800 198768 239148 199848
rect 880 198488 239148 198768
rect 800 196048 239148 198488
rect 800 195768 239068 196048
rect 800 194688 239148 195768
rect 880 194408 239148 194688
rect 800 191968 239148 194408
rect 800 191688 239068 191968
rect 800 190608 239148 191688
rect 880 190328 239148 190608
rect 800 187888 239148 190328
rect 800 187608 239068 187888
rect 800 186528 239148 187608
rect 880 186248 239148 186528
rect 800 183808 239148 186248
rect 800 183528 239068 183808
rect 800 182448 239148 183528
rect 880 182168 239148 182448
rect 800 179048 239148 182168
rect 800 178768 239068 179048
rect 800 177688 239148 178768
rect 880 177408 239148 177688
rect 800 174968 239148 177408
rect 800 174688 239068 174968
rect 800 173608 239148 174688
rect 880 173328 239148 173608
rect 800 170888 239148 173328
rect 800 170608 239068 170888
rect 800 169528 239148 170608
rect 880 169248 239148 169528
rect 800 166808 239148 169248
rect 800 166528 239068 166808
rect 800 165448 239148 166528
rect 880 165168 239148 165448
rect 800 162728 239148 165168
rect 800 162448 239068 162728
rect 800 161368 239148 162448
rect 880 161088 239148 161368
rect 800 158648 239148 161088
rect 800 158368 239068 158648
rect 800 157288 239148 158368
rect 880 157008 239148 157288
rect 800 154568 239148 157008
rect 800 154288 239068 154568
rect 800 153208 239148 154288
rect 880 152928 239148 153208
rect 800 150488 239148 152928
rect 800 150208 239068 150488
rect 800 149128 239148 150208
rect 880 148848 239148 149128
rect 800 146408 239148 148848
rect 800 146128 239068 146408
rect 800 145048 239148 146128
rect 880 144768 239148 145048
rect 800 142328 239148 144768
rect 800 142048 239068 142328
rect 800 140968 239148 142048
rect 880 140688 239148 140968
rect 800 138248 239148 140688
rect 800 137968 239068 138248
rect 800 136888 239148 137968
rect 880 136608 239148 136888
rect 800 134168 239148 136608
rect 800 133888 239068 134168
rect 800 132808 239148 133888
rect 880 132528 239148 132808
rect 800 130088 239148 132528
rect 800 129808 239068 130088
rect 800 128728 239148 129808
rect 880 128448 239148 128728
rect 800 126008 239148 128448
rect 800 125728 239068 126008
rect 800 124648 239148 125728
rect 880 124368 239148 124648
rect 800 121248 239148 124368
rect 800 120968 239068 121248
rect 800 120568 239148 120968
rect 880 120288 239148 120568
rect 800 117168 239148 120288
rect 800 116888 239068 117168
rect 800 115808 239148 116888
rect 880 115528 239148 115808
rect 800 113088 239148 115528
rect 800 112808 239068 113088
rect 800 111728 239148 112808
rect 880 111448 239148 111728
rect 800 109008 239148 111448
rect 800 108728 239068 109008
rect 800 107648 239148 108728
rect 880 107368 239148 107648
rect 800 104928 239148 107368
rect 800 104648 239068 104928
rect 800 103568 239148 104648
rect 880 103288 239148 103568
rect 800 100848 239148 103288
rect 800 100568 239068 100848
rect 800 99488 239148 100568
rect 880 99208 239148 99488
rect 800 96768 239148 99208
rect 800 96488 239068 96768
rect 800 95408 239148 96488
rect 880 95128 239148 95408
rect 800 92688 239148 95128
rect 800 92408 239068 92688
rect 800 91328 239148 92408
rect 880 91048 239148 91328
rect 800 88608 239148 91048
rect 800 88328 239068 88608
rect 800 87248 239148 88328
rect 880 86968 239148 87248
rect 800 84528 239148 86968
rect 800 84248 239068 84528
rect 800 83168 239148 84248
rect 880 82888 239148 83168
rect 800 80448 239148 82888
rect 800 80168 239068 80448
rect 800 79088 239148 80168
rect 880 78808 239148 79088
rect 800 76368 239148 78808
rect 800 76088 239068 76368
rect 800 75008 239148 76088
rect 880 74728 239148 75008
rect 800 72288 239148 74728
rect 800 72008 239068 72288
rect 800 70928 239148 72008
rect 880 70648 239148 70928
rect 800 68208 239148 70648
rect 800 67928 239068 68208
rect 800 66848 239148 67928
rect 880 66568 239148 66848
rect 800 64128 239148 66568
rect 800 63848 239068 64128
rect 800 62768 239148 63848
rect 880 62488 239148 62768
rect 800 59368 239148 62488
rect 800 59088 239068 59368
rect 800 58008 239148 59088
rect 880 57728 239148 58008
rect 800 55288 239148 57728
rect 800 55008 239068 55288
rect 800 53928 239148 55008
rect 880 53648 239148 53928
rect 800 51208 239148 53648
rect 800 50928 239068 51208
rect 800 49848 239148 50928
rect 880 49568 239148 49848
rect 800 47128 239148 49568
rect 800 46848 239068 47128
rect 800 45768 239148 46848
rect 880 45488 239148 45768
rect 800 43048 239148 45488
rect 800 42768 239068 43048
rect 800 41688 239148 42768
rect 880 41408 239148 41688
rect 800 38968 239148 41408
rect 800 38688 239068 38968
rect 800 37608 239148 38688
rect 880 37328 239148 37608
rect 800 34888 239148 37328
rect 800 34608 239068 34888
rect 800 33528 239148 34608
rect 880 33248 239148 33528
rect 800 30808 239148 33248
rect 800 30528 239068 30808
rect 800 29448 239148 30528
rect 880 29168 239148 29448
rect 800 26728 239148 29168
rect 800 26448 239068 26728
rect 800 25368 239148 26448
rect 880 25088 239148 25368
rect 800 22648 239148 25088
rect 800 22368 239068 22648
rect 800 21288 239148 22368
rect 880 21008 239148 21288
rect 800 18568 239148 21008
rect 800 18288 239068 18568
rect 800 17208 239148 18288
rect 880 16928 239148 17208
rect 800 14488 239148 16928
rect 800 14208 239068 14488
rect 800 13128 239148 14208
rect 880 12848 239148 13128
rect 800 10408 239148 12848
rect 800 10128 239068 10408
rect 800 9048 239148 10128
rect 880 8768 239148 9048
rect 800 6328 239148 8768
rect 800 6048 239068 6328
rect 800 4968 239148 6048
rect 880 4688 239148 4968
rect 800 1568 239148 4688
rect 800 1395 239068 1568
<< metal4 >>
rect 4208 2128 4528 239952
rect 9208 2128 9528 239952
rect 14208 2128 14528 239952
rect 19208 100452 19528 239952
rect 24208 100452 24528 239952
rect 29208 100452 29528 239952
rect 34208 100452 34528 239952
rect 39208 100452 39528 239952
rect 44208 100452 44528 239952
rect 49208 100452 49528 239952
rect 54208 100452 54528 239952
rect 59208 100452 59528 239952
rect 64208 100452 64528 239952
rect 69208 100452 69528 239952
rect 74208 100452 74528 239952
rect 79208 100452 79528 239952
rect 84208 100452 84528 239952
rect 89208 100452 89528 239952
rect 94208 100452 94528 239952
rect 99208 100452 99528 239952
rect 104208 100452 104528 239952
rect 109208 100452 109528 239952
rect 114208 100452 114528 239952
rect 19208 2128 19528 19048
rect 24208 2128 24528 19048
rect 29208 2128 29528 19048
rect 34208 2128 34528 19048
rect 39208 2128 39528 19048
rect 44208 2128 44528 19048
rect 49208 2128 49528 19048
rect 54208 2128 54528 19048
rect 59208 2128 59528 19048
rect 64208 2128 64528 19048
rect 69208 2128 69528 19048
rect 74208 2128 74528 19048
rect 79208 2128 79528 19048
rect 84208 2128 84528 19048
rect 89208 2128 89528 19048
rect 94208 2128 94528 19048
rect 99208 2128 99528 19048
rect 104208 2128 104528 19048
rect 109208 2128 109528 19048
rect 114208 2128 114528 19048
rect 119208 2128 119528 239952
rect 124208 2128 124528 239952
rect 129208 2128 129528 239952
rect 134208 2128 134528 239952
rect 139208 2128 139528 239952
rect 144208 2128 144528 239952
rect 149208 2128 149528 239952
rect 154208 2128 154528 239952
rect 159208 2128 159528 239952
rect 164208 2128 164528 239952
rect 169208 2128 169528 239952
rect 174208 2128 174528 239952
rect 179208 2128 179528 239952
rect 184208 2128 184528 239952
rect 189208 2128 189528 239952
rect 194208 2128 194528 239952
rect 199208 2128 199528 239952
rect 204208 2128 204528 239952
rect 209208 2128 209528 239952
rect 214208 2128 214528 239952
rect 219208 2128 219528 239952
rect 224208 2128 224528 239952
rect 229208 2128 229528 239952
rect 234208 2128 234528 239952
<< obsm4 >>
rect 19011 240032 215221 240549
rect 19011 100372 19128 240032
rect 19608 100372 24128 240032
rect 24608 100372 29128 240032
rect 29608 100372 34128 240032
rect 34608 100372 39128 240032
rect 39608 100372 44128 240032
rect 44608 100372 49128 240032
rect 49608 100372 54128 240032
rect 54608 100372 59128 240032
rect 59608 100372 64128 240032
rect 64608 100372 69128 240032
rect 69608 100372 74128 240032
rect 74608 100372 79128 240032
rect 79608 100372 84128 240032
rect 84608 100372 89128 240032
rect 89608 100372 94128 240032
rect 94608 100372 99128 240032
rect 99608 100372 104128 240032
rect 104608 100372 109128 240032
rect 109608 100372 114128 240032
rect 114608 100372 119128 240032
rect 19011 19128 119128 100372
rect 19011 2048 19128 19128
rect 19608 2048 24128 19128
rect 24608 2048 29128 19128
rect 29608 2048 34128 19128
rect 34608 2048 39128 19128
rect 39608 2048 44128 19128
rect 44608 2048 49128 19128
rect 49608 2048 54128 19128
rect 54608 2048 59128 19128
rect 59608 2048 64128 19128
rect 64608 2048 69128 19128
rect 69608 2048 74128 19128
rect 74608 2048 79128 19128
rect 79608 2048 84128 19128
rect 84608 2048 89128 19128
rect 89608 2048 94128 19128
rect 94608 2048 99128 19128
rect 99608 2048 104128 19128
rect 104608 2048 109128 19128
rect 109608 2048 114128 19128
rect 114608 2048 119128 19128
rect 119608 2048 124128 240032
rect 124608 2048 129128 240032
rect 129608 2048 134128 240032
rect 134608 2048 139128 240032
rect 139608 2048 144128 240032
rect 144608 2048 149128 240032
rect 149608 2048 154128 240032
rect 154608 2048 159128 240032
rect 159608 2048 164128 240032
rect 164608 2048 169128 240032
rect 169608 2048 174128 240032
rect 174608 2048 179128 240032
rect 179608 2048 184128 240032
rect 184608 2048 189128 240032
rect 189608 2048 194128 240032
rect 194608 2048 199128 240032
rect 199608 2048 204128 240032
rect 204608 2048 209128 240032
rect 209608 2048 214128 240032
rect 214608 2048 215221 240032
rect 19011 1803 215221 2048
<< metal5 >>
rect 1104 235068 238832 235388
rect 1104 219750 238832 220070
rect 1104 204432 238832 204752
rect 1104 189114 238832 189434
rect 1104 173796 238832 174116
rect 1104 158478 238832 158798
rect 1104 143160 238832 143480
rect 1104 127842 238832 128162
rect 1104 112524 238832 112844
rect 1104 97206 238832 97526
rect 1104 81888 238832 82208
rect 1104 66570 238832 66890
rect 1104 51252 238832 51572
rect 1104 35934 238832 36254
rect 1104 20616 238832 20936
rect 1104 5298 238832 5618
<< labels >>
rlabel metal3 s 0 29248 800 29368 6 clk_i
port 1 nsew signal input
rlabel metal3 s 239148 183608 239948 183728 6 debug_req_i
port 2 nsew signal input
rlabel metal2 s 233698 241292 233754 242092 6 eFPGA_delay_o[0]
port 3 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 eFPGA_delay_o[1]
port 4 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 eFPGA_delay_o[2]
port 5 nsew signal output
rlabel metal2 s 172518 241292 172574 242092 6 eFPGA_delay_o[3]
port 6 nsew signal output
rlabel metal2 s 88798 241292 88854 242092 6 eFPGA_en_o
port 7 nsew signal output
rlabel metal2 s 103518 0 103574 800 6 eFPGA_fpga_done_i
port 8 nsew signal input
rlabel metal3 s 239148 174768 239948 174888 6 eFPGA_operand_a_o[0]
port 9 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 eFPGA_operand_a_o[10]
port 10 nsew signal output
rlabel metal3 s 0 231208 800 231328 6 eFPGA_operand_a_o[11]
port 11 nsew signal output
rlabel metal2 s 234618 0 234674 800 6 eFPGA_operand_a_o[12]
port 12 nsew signal output
rlabel metal2 s 72698 0 72754 800 6 eFPGA_operand_a_o[13]
port 13 nsew signal output
rlabel metal2 s 148138 0 148194 800 6 eFPGA_operand_a_o[14]
port 14 nsew signal output
rlabel metal2 s 228178 241292 228234 242092 6 eFPGA_operand_a_o[15]
port 15 nsew signal output
rlabel metal3 s 239148 104728 239948 104848 6 eFPGA_operand_a_o[16]
port 16 nsew signal output
rlabel metal2 s 203338 241292 203394 242092 6 eFPGA_operand_a_o[17]
port 17 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 eFPGA_operand_a_o[18]
port 18 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 eFPGA_operand_a_o[19]
port 19 nsew signal output
rlabel metal2 s 16118 241292 16174 242092 6 eFPGA_operand_a_o[1]
port 20 nsew signal output
rlabel metal3 s 0 66648 800 66768 6 eFPGA_operand_a_o[20]
port 21 nsew signal output
rlabel metal3 s 239148 158448 239948 158568 6 eFPGA_operand_a_o[21]
port 22 nsew signal output
rlabel metal3 s 239148 34688 239948 34808 6 eFPGA_operand_a_o[22]
port 23 nsew signal output
rlabel metal3 s 239148 46928 239948 47048 6 eFPGA_operand_a_o[23]
port 24 nsew signal output
rlabel metal3 s 0 210808 800 210928 6 eFPGA_operand_a_o[24]
port 25 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 eFPGA_operand_a_o[25]
port 26 nsew signal output
rlabel metal3 s 239148 204008 239948 204128 6 eFPGA_operand_a_o[26]
port 27 nsew signal output
rlabel metal3 s 239148 195848 239948 195968 6 eFPGA_operand_a_o[27]
port 28 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 eFPGA_operand_a_o[28]
port 29 nsew signal output
rlabel metal2 s 166998 241292 167054 242092 6 eFPGA_operand_a_o[29]
port 30 nsew signal output
rlabel metal3 s 239148 63928 239948 64048 6 eFPGA_operand_a_o[2]
port 31 nsew signal output
rlabel metal2 s 201498 0 201554 800 6 eFPGA_operand_a_o[30]
port 32 nsew signal output
rlabel metal2 s 144458 241292 144514 242092 6 eFPGA_operand_a_o[31]
port 33 nsew signal output
rlabel metal2 s 229098 0 229154 800 6 eFPGA_operand_a_o[3]
port 34 nsew signal output
rlabel metal2 s 222658 241292 222714 242092 6 eFPGA_operand_a_o[4]
port 35 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 eFPGA_operand_a_o[5]
port 36 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 eFPGA_operand_a_o[6]
port 37 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 eFPGA_operand_a_o[7]
port 38 nsew signal output
rlabel metal2 s 173438 0 173494 800 6 eFPGA_operand_a_o[8]
port 39 nsew signal output
rlabel metal2 s 110878 241292 110934 242092 6 eFPGA_operand_a_o[9]
port 40 nsew signal output
rlabel metal3 s 239148 212168 239948 212288 6 eFPGA_operand_b_o[0]
port 41 nsew signal output
rlabel metal3 s 239148 220328 239948 220448 6 eFPGA_operand_b_o[10]
port 42 nsew signal output
rlabel metal2 s 130658 241292 130714 242092 6 eFPGA_operand_b_o[11]
port 43 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 eFPGA_operand_b_o[12]
port 44 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 eFPGA_operand_b_o[13]
port 45 nsew signal output
rlabel metal2 s 149978 241292 150034 242092 6 eFPGA_operand_b_o[14]
port 46 nsew signal output
rlabel metal2 s 86038 241292 86094 242092 6 eFPGA_operand_b_o[15]
port 47 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 eFPGA_operand_b_o[16]
port 48 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 eFPGA_operand_b_o[17]
port 49 nsew signal output
rlabel metal2 s 223578 0 223634 800 6 eFPGA_operand_b_o[18]
port 50 nsew signal output
rlabel metal2 s 41418 241292 41474 242092 6 eFPGA_operand_b_o[19]
port 51 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 eFPGA_operand_b_o[1]
port 52 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 eFPGA_operand_b_o[20]
port 53 nsew signal output
rlabel metal3 s 239148 116968 239948 117088 6 eFPGA_operand_b_o[21]
port 54 nsew signal output
rlabel metal2 s 158258 241292 158314 242092 6 eFPGA_operand_b_o[22]
port 55 nsew signal output
rlabel metal2 s 113638 241292 113694 242092 6 eFPGA_operand_b_o[23]
port 56 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 eFPGA_operand_b_o[24]
port 57 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 eFPGA_operand_b_o[25]
port 58 nsew signal output
rlabel metal2 s 162398 0 162454 800 6 eFPGA_operand_b_o[26]
port 59 nsew signal output
rlabel metal2 s 11518 0 11574 800 6 eFPGA_operand_b_o[27]
port 60 nsew signal output
rlabel metal2 s 29918 241292 29974 242092 6 eFPGA_operand_b_o[28]
port 61 nsew signal output
rlabel metal2 s 167918 0 167974 800 6 eFPGA_operand_b_o[29]
port 62 nsew signal output
rlabel metal3 s 239148 146208 239948 146328 6 eFPGA_operand_b_o[2]
port 63 nsew signal output
rlabel metal3 s 239148 68008 239948 68128 6 eFPGA_operand_b_o[30]
port 64 nsew signal output
rlabel metal2 s 89718 0 89774 800 6 eFPGA_operand_b_o[31]
port 65 nsew signal output
rlabel metal3 s 0 144848 800 144968 6 eFPGA_operand_b_o[3]
port 66 nsew signal output
rlabel metal3 s 0 182248 800 182368 6 eFPGA_operand_b_o[4]
port 67 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 eFPGA_operand_b_o[5]
port 68 nsew signal output
rlabel metal2 s 155498 241292 155554 242092 6 eFPGA_operand_b_o[6]
port 69 nsew signal output
rlabel metal3 s 0 153008 800 153128 6 eFPGA_operand_b_o[7]
port 70 nsew signal output
rlabel metal2 s 186318 241292 186374 242092 6 eFPGA_operand_b_o[8]
port 71 nsew signal output
rlabel metal2 s 189998 0 190054 800 6 eFPGA_operand_b_o[9]
port 72 nsew signal output
rlabel metal3 s 0 107448 800 107568 6 eFPGA_operator_o[0]
port 73 nsew signal output
rlabel metal3 s 239148 142128 239948 142248 6 eFPGA_operator_o[1]
port 74 nsew signal output
rlabel metal2 s 57978 241292 58034 242092 6 eFPGA_result_a_i[0]
port 75 nsew signal input
rlabel metal3 s 0 169328 800 169448 6 eFPGA_result_a_i[10]
port 76 nsew signal input
rlabel metal2 s 152738 241292 152794 242092 6 eFPGA_result_a_i[11]
port 77 nsew signal input
rlabel metal3 s 0 214888 800 215008 6 eFPGA_result_a_i[12]
port 78 nsew signal input
rlabel metal3 s 239148 216248 239948 216368 6 eFPGA_result_a_i[13]
port 79 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 eFPGA_result_a_i[14]
port 80 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 eFPGA_result_a_i[15]
port 81 nsew signal input
rlabel metal2 s 183558 241292 183614 242092 6 eFPGA_result_a_i[16]
port 82 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 eFPGA_result_a_i[17]
port 83 nsew signal input
rlabel metal2 s 55218 241292 55274 242092 6 eFPGA_result_a_i[18]
port 84 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 eFPGA_result_a_i[19]
port 85 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 eFPGA_result_a_i[1]
port 86 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 eFPGA_result_a_i[20]
port 87 nsew signal input
rlabel metal2 s 95238 0 95294 800 6 eFPGA_result_a_i[21]
port 88 nsew signal input
rlabel metal3 s 239148 18368 239948 18488 6 eFPGA_result_a_i[22]
port 89 nsew signal input
rlabel metal3 s 0 161168 800 161288 6 eFPGA_result_a_i[23]
port 90 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 eFPGA_result_a_i[24]
port 91 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 eFPGA_result_a_i[25]
port 92 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 eFPGA_result_a_i[26]
port 93 nsew signal input
rlabel metal3 s 0 198568 800 198688 6 eFPGA_result_a_i[27]
port 94 nsew signal input
rlabel metal2 s 119618 241292 119674 242092 6 eFPGA_result_a_i[28]
port 95 nsew signal input
rlabel metal2 s 156418 0 156474 800 6 eFPGA_result_a_i[29]
port 96 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 eFPGA_result_a_i[2]
port 97 nsew signal input
rlabel metal3 s 239148 187688 239948 187808 6 eFPGA_result_a_i[30]
port 98 nsew signal input
rlabel metal2 s 116398 241292 116454 242092 6 eFPGA_result_a_i[31]
port 99 nsew signal input
rlabel metal2 s 189078 241292 189134 242092 6 eFPGA_result_a_i[3]
port 100 nsew signal input
rlabel metal2 s 102598 241292 102654 242092 6 eFPGA_result_a_i[4]
port 101 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 eFPGA_result_a_i[5]
port 102 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 eFPGA_result_a_i[6]
port 103 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 eFPGA_result_a_i[7]
port 104 nsew signal input
rlabel metal2 s 217138 241292 217194 242092 6 eFPGA_result_a_i[8]
port 105 nsew signal input
rlabel metal2 s 105358 241292 105414 242092 6 eFPGA_result_a_i[9]
port 106 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 eFPGA_result_b_i[0]
port 107 nsew signal input
rlabel metal3 s 239148 112888 239948 113008 6 eFPGA_result_b_i[10]
port 108 nsew signal input
rlabel metal2 s 200578 241292 200634 242092 6 eFPGA_result_b_i[11]
port 109 nsew signal input
rlabel metal3 s 239148 100648 239948 100768 6 eFPGA_result_b_i[12]
port 110 nsew signal input
rlabel metal2 s 99838 241292 99894 242092 6 eFPGA_result_b_i[13]
port 111 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 eFPGA_result_b_i[14]
port 112 nsew signal input
rlabel metal2 s 7838 241292 7894 242092 6 eFPGA_result_b_i[15]
port 113 nsew signal input
rlabel metal3 s 239148 224408 239948 224528 6 eFPGA_result_b_i[16]
port 114 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 eFPGA_result_b_i[17]
port 115 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 eFPGA_result_b_i[18]
port 116 nsew signal input
rlabel metal2 s 180798 241292 180854 242092 6 eFPGA_result_b_i[19]
port 117 nsew signal input
rlabel metal2 s 181718 0 181774 800 6 eFPGA_result_b_i[1]
port 118 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 eFPGA_result_b_i[20]
port 119 nsew signal input
rlabel metal2 s 138938 241292 138994 242092 6 eFPGA_result_b_i[21]
port 120 nsew signal input
rlabel metal3 s 0 240048 800 240168 6 eFPGA_result_b_i[22]
port 121 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 eFPGA_result_b_i[23]
port 122 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 eFPGA_result_b_i[24]
port 123 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 eFPGA_result_b_i[25]
port 124 nsew signal input
rlabel metal2 s 125138 241292 125194 242092 6 eFPGA_result_b_i[26]
port 125 nsew signal input
rlabel metal3 s 0 227128 800 227248 6 eFPGA_result_b_i[27]
port 126 nsew signal input
rlabel metal3 s 239148 191768 239948 191888 6 eFPGA_result_b_i[28]
port 127 nsew signal input
rlabel metal3 s 239148 199928 239948 200048 6 eFPGA_result_b_i[29]
port 128 nsew signal input
rlabel metal2 s 46938 241292 46994 242092 6 eFPGA_result_b_i[2]
port 129 nsew signal input
rlabel metal2 s 10598 241292 10654 242092 6 eFPGA_result_b_i[30]
port 130 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 eFPGA_result_b_i[31]
port 131 nsew signal input
rlabel metal2 s 219898 241292 219954 242092 6 eFPGA_result_b_i[3]
port 132 nsew signal input
rlabel metal3 s 239148 208088 239948 208208 6 eFPGA_result_b_i[4]
port 133 nsew signal input
rlabel metal3 s 0 173408 800 173528 6 eFPGA_result_b_i[5]
port 134 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 eFPGA_result_b_i[6]
port 135 nsew signal input
rlabel metal3 s 239148 10208 239948 10328 6 eFPGA_result_b_i[7]
port 136 nsew signal input
rlabel metal2 s 176198 0 176254 800 6 eFPGA_result_b_i[8]
port 137 nsew signal input
rlabel metal2 s 97078 241292 97134 242092 6 eFPGA_result_b_i[9]
port 138 nsew signal input
rlabel metal2 s 133418 241292 133474 242092 6 eFPGA_result_c_i[0]
port 139 nsew signal input
rlabel metal2 s 178038 241292 178094 242092 6 eFPGA_result_c_i[10]
port 140 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 eFPGA_result_c_i[11]
port 141 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 eFPGA_result_c_i[12]
port 142 nsew signal input
rlabel metal2 s 209778 0 209834 800 6 eFPGA_result_c_i[13]
port 143 nsew signal input
rlabel metal2 s 147218 241292 147274 242092 6 eFPGA_result_c_i[14]
port 144 nsew signal input
rlabel metal3 s 239148 42848 239948 42968 6 eFPGA_result_c_i[15]
port 145 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 eFPGA_result_c_i[16]
port 146 nsew signal input
rlabel metal3 s 0 186328 800 186448 6 eFPGA_result_c_i[17]
port 147 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 eFPGA_result_c_i[18]
port 148 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 eFPGA_result_c_i[19]
port 149 nsew signal input
rlabel metal2 s 215298 0 215354 800 6 eFPGA_result_c_i[1]
port 150 nsew signal input
rlabel metal3 s 239148 26528 239948 26648 6 eFPGA_result_c_i[20]
port 151 nsew signal input
rlabel metal3 s 239148 55088 239948 55208 6 eFPGA_result_c_i[21]
port 152 nsew signal input
rlabel metal2 s 478 0 534 800 6 eFPGA_result_c_i[22]
port 153 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 eFPGA_result_c_i[23]
port 154 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 eFPGA_result_c_i[24]
port 155 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 eFPGA_result_c_i[25]
port 156 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 eFPGA_result_c_i[26]
port 157 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 eFPGA_result_c_i[27]
port 158 nsew signal input
rlabel metal2 s 71778 241292 71834 242092 6 eFPGA_result_c_i[28]
port 159 nsew signal input
rlabel metal2 s 32678 241292 32734 242092 6 eFPGA_result_c_i[29]
port 160 nsew signal input
rlabel metal2 s 178958 0 179014 800 6 eFPGA_result_c_i[2]
port 161 nsew signal input
rlabel metal2 s 214378 241292 214434 242092 6 eFPGA_result_c_i[30]
port 162 nsew signal input
rlabel metal3 s 0 194488 800 194608 6 eFPGA_result_c_i[31]
port 163 nsew signal input
rlabel metal2 s 24398 241292 24454 242092 6 eFPGA_result_c_i[3]
port 164 nsew signal input
rlabel metal2 s 142618 0 142674 800 6 eFPGA_result_c_i[4]
port 165 nsew signal input
rlabel metal3 s 239148 96568 239948 96688 6 eFPGA_result_c_i[5]
port 166 nsew signal input
rlabel metal2 s 136178 241292 136234 242092 6 eFPGA_result_c_i[6]
port 167 nsew signal input
rlabel metal2 s 236458 241292 236514 242092 6 eFPGA_result_c_i[7]
port 168 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 eFPGA_result_c_i[8]
port 169 nsew signal input
rlabel metal3 s 239148 84328 239948 84448 6 eFPGA_result_c_i[9]
port 170 nsew signal input
rlabel metal2 s 77298 241292 77354 242092 6 eFPGA_write_strobe_o
port 171 nsew signal output
rlabel metal2 s 231858 0 231914 800 6 ext_data_addr_i[0]
port 172 nsew signal input
rlabel metal3 s 239148 236648 239948 236768 6 ext_data_addr_i[10]
port 173 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 ext_data_addr_i[11]
port 174 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 ext_data_addr_i[12]
port 175 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 ext_data_addr_i[13]
port 176 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 ext_data_addr_i[14]
port 177 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 ext_data_addr_i[15]
port 178 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 ext_data_addr_i[16]
port 179 nsew signal input
rlabel metal2 s 80518 241292 80574 242092 6 ext_data_addr_i[17]
port 180 nsew signal input
rlabel metal2 s 204258 0 204314 800 6 ext_data_addr_i[18]
port 181 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 ext_data_addr_i[19]
port 182 nsew signal input
rlabel metal3 s 239148 121048 239948 121168 6 ext_data_addr_i[1]
port 183 nsew signal input
rlabel metal2 s 18878 241292 18934 242092 6 ext_data_addr_i[20]
port 184 nsew signal input
rlabel metal3 s 239148 166608 239948 166728 6 ext_data_addr_i[21]
port 185 nsew signal input
rlabel metal2 s 69018 241292 69074 242092 6 ext_data_addr_i[22]
port 186 nsew signal input
rlabel metal3 s 239148 59168 239948 59288 6 ext_data_addr_i[23]
port 187 nsew signal input
rlabel metal2 s 212538 0 212594 800 6 ext_data_addr_i[24]
port 188 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 ext_data_addr_i[25]
port 189 nsew signal input
rlabel metal3 s 239148 232568 239948 232688 6 ext_data_addr_i[26]
port 190 nsew signal input
rlabel metal2 s 49698 241292 49754 242092 6 ext_data_addr_i[27]
port 191 nsew signal input
rlabel metal2 s 169758 241292 169814 242092 6 ext_data_addr_i[28]
port 192 nsew signal input
rlabel metal2 s 191838 241292 191894 242092 6 ext_data_addr_i[29]
port 193 nsew signal input
rlabel metal2 s 198278 0 198334 800 6 ext_data_addr_i[2]
port 194 nsew signal input
rlabel metal2 s 83278 241292 83334 242092 6 ext_data_addr_i[30]
port 195 nsew signal input
rlabel metal2 s 108118 241292 108174 242092 6 ext_data_addr_i[31]
port 196 nsew signal input
rlabel metal2 s 60738 241292 60794 242092 6 ext_data_addr_i[3]
port 197 nsew signal input
rlabel metal2 s 225418 241292 225474 242092 6 ext_data_addr_i[4]
port 198 nsew signal input
rlabel metal3 s 239148 30608 239948 30728 6 ext_data_addr_i[5]
port 199 nsew signal input
rlabel metal2 s 44178 241292 44234 242092 6 ext_data_addr_i[6]
port 200 nsew signal input
rlabel metal2 s 74538 241292 74594 242092 6 ext_data_addr_i[7]
port 201 nsew signal input
rlabel metal3 s 0 206728 800 206848 6 ext_data_addr_i[8]
port 202 nsew signal input
rlabel metal3 s 0 202648 800 202768 6 ext_data_addr_i[9]
port 203 nsew signal input
rlabel metal2 s 27158 241292 27214 242092 6 ext_data_be_i[0]
port 204 nsew signal input
rlabel metal3 s 239148 22448 239948 22568 6 ext_data_be_i[1]
port 205 nsew signal input
rlabel metal2 s 13358 241292 13414 242092 6 ext_data_be_i[2]
port 206 nsew signal input
rlabel metal3 s 0 165248 800 165368 6 ext_data_be_i[3]
port 207 nsew signal input
rlabel metal3 s 0 218968 800 219088 6 ext_data_rdata_o[0]
port 208 nsew signal output
rlabel metal2 s 220818 0 220874 800 6 ext_data_rdata_o[10]
port 209 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 ext_data_rdata_o[11]
port 210 nsew signal output
rlabel metal3 s 239148 150288 239948 150408 6 ext_data_rdata_o[12]
port 211 nsew signal output
rlabel metal2 s 122378 241292 122434 242092 6 ext_data_rdata_o[13]
port 212 nsew signal output
rlabel metal3 s 239148 162528 239948 162648 6 ext_data_rdata_o[14]
port 213 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 ext_data_rdata_o[15]
port 214 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 ext_data_rdata_o[16]
port 215 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 ext_data_rdata_o[17]
port 216 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 ext_data_rdata_o[18]
port 217 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 ext_data_rdata_o[19]
port 218 nsew signal output
rlabel metal3 s 239148 133968 239948 134088 6 ext_data_rdata_o[1]
port 219 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 ext_data_rdata_o[20]
port 220 nsew signal output
rlabel metal3 s 239148 6128 239948 6248 6 ext_data_rdata_o[21]
port 221 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 ext_data_rdata_o[22]
port 222 nsew signal output
rlabel metal3 s 239148 72088 239948 72208 6 ext_data_rdata_o[23]
port 223 nsew signal output
rlabel metal2 s 61658 0 61714 800 6 ext_data_rdata_o[24]
port 224 nsew signal output
rlabel metal2 s 194598 241292 194654 242092 6 ext_data_rdata_o[25]
port 225 nsew signal output
rlabel metal3 s 0 223048 800 223168 6 ext_data_rdata_o[26]
port 226 nsew signal output
rlabel metal2 s 38198 241292 38254 242092 6 ext_data_rdata_o[27]
port 227 nsew signal output
rlabel metal2 s 187238 0 187294 800 6 ext_data_rdata_o[28]
port 228 nsew signal output
rlabel metal2 s 239218 241292 239274 242092 6 ext_data_rdata_o[29]
port 229 nsew signal output
rlabel metal2 s 126058 0 126114 800 6 ext_data_rdata_o[2]
port 230 nsew signal output
rlabel metal2 s 237378 0 237434 800 6 ext_data_rdata_o[30]
port 231 nsew signal output
rlabel metal2 s 21638 241292 21694 242092 6 ext_data_rdata_o[31]
port 232 nsew signal output
rlabel metal3 s 239148 38768 239948 38888 6 ext_data_rdata_o[3]
port 233 nsew signal output
rlabel metal3 s 239148 138048 239948 138168 6 ext_data_rdata_o[4]
port 234 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 ext_data_rdata_o[5]
port 235 nsew signal output
rlabel metal3 s 239148 76168 239948 76288 6 ext_data_rdata_o[6]
port 236 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 ext_data_rdata_o[7]
port 237 nsew signal output
rlabel metal2 s 175278 241292 175334 242092 6 ext_data_rdata_o[8]
port 238 nsew signal output
rlabel metal2 s 164238 241292 164294 242092 6 ext_data_rdata_o[9]
port 239 nsew signal output
rlabel metal2 s 2318 241292 2374 242092 6 ext_data_req_i
port 240 nsew signal input
rlabel metal2 s 66258 241292 66314 242092 6 ext_data_rvalid_o
port 241 nsew signal output
rlabel metal2 s 35438 241292 35494 242092 6 ext_data_wdata_i[0]
port 242 nsew signal input
rlabel metal3 s 239148 228488 239948 228608 6 ext_data_wdata_i[10]
port 243 nsew signal input
rlabel metal2 s 153658 0 153714 800 6 ext_data_wdata_i[11]
port 244 nsew signal input
rlabel metal3 s 239148 108808 239948 108928 6 ext_data_wdata_i[12]
port 245 nsew signal input
rlabel metal3 s 239148 80248 239948 80368 6 ext_data_wdata_i[13]
port 246 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 ext_data_wdata_i[14]
port 247 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 ext_data_wdata_i[15]
port 248 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 ext_data_wdata_i[16]
port 249 nsew signal input
rlabel metal2 s 195518 0 195574 800 6 ext_data_wdata_i[17]
port 250 nsew signal input
rlabel metal3 s 239148 129888 239948 130008 6 ext_data_wdata_i[18]
port 251 nsew signal input
rlabel metal2 s 206098 241292 206154 242092 6 ext_data_wdata_i[19]
port 252 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 ext_data_wdata_i[1]
port 253 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 ext_data_wdata_i[20]
port 254 nsew signal input
rlabel metal3 s 239148 170688 239948 170808 6 ext_data_wdata_i[21]
port 255 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 ext_data_wdata_i[22]
port 256 nsew signal input
rlabel metal3 s 0 235288 800 235408 6 ext_data_wdata_i[23]
port 257 nsew signal input
rlabel metal2 s 230938 241292 230994 242092 6 ext_data_wdata_i[24]
port 258 nsew signal input
rlabel metal2 s 161478 241292 161534 242092 6 ext_data_wdata_i[25]
port 259 nsew signal input
rlabel metal2 s 127898 241292 127954 242092 6 ext_data_wdata_i[26]
port 260 nsew signal input
rlabel metal2 s 218058 0 218114 800 6 ext_data_wdata_i[27]
port 261 nsew signal input
rlabel metal3 s 239148 125808 239948 125928 6 ext_data_wdata_i[28]
port 262 nsew signal input
rlabel metal3 s 0 132608 800 132728 6 ext_data_wdata_i[29]
port 263 nsew signal input
rlabel metal3 s 239148 92488 239948 92608 6 ext_data_wdata_i[2]
port 264 nsew signal input
rlabel metal2 s 211618 241292 211674 242092 6 ext_data_wdata_i[30]
port 265 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 ext_data_wdata_i[31]
port 266 nsew signal input
rlabel metal2 s 52458 241292 52514 242092 6 ext_data_wdata_i[3]
port 267 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 ext_data_wdata_i[4]
port 268 nsew signal input
rlabel metal3 s 239148 178848 239948 178968 6 ext_data_wdata_i[5]
port 269 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 ext_data_wdata_i[6]
port 270 nsew signal input
rlabel metal2 s 5078 241292 5134 242092 6 ext_data_wdata_i[7]
port 271 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 ext_data_wdata_i[8]
port 272 nsew signal input
rlabel metal2 s 63498 241292 63554 242092 6 ext_data_wdata_i[9]
port 273 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 ext_data_we_i
port 274 nsew signal input
rlabel metal3 s 239148 1368 239948 1488 6 fetch_enable_i
port 275 nsew signal input
rlabel metal2 s 91558 241292 91614 242092 6 irq_ack_o
port 276 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 irq_i
port 277 nsew signal input
rlabel metal2 s 197358 241292 197414 242092 6 irq_id_i[0]
port 278 nsew signal input
rlabel metal3 s 0 177488 800 177608 6 irq_id_i[1]
port 279 nsew signal input
rlabel metal2 s 94318 241292 94374 242092 6 irq_id_i[2]
port 280 nsew signal input
rlabel metal3 s 239148 88408 239948 88528 6 irq_id_i[3]
port 281 nsew signal input
rlabel metal3 s 239148 14288 239948 14408 6 irq_id_i[4]
port 282 nsew signal input
rlabel metal2 s 141698 241292 141754 242092 6 irq_id_o[0]
port 283 nsew signal output
rlabel metal3 s 239148 51008 239948 51128 6 irq_id_o[1]
port 284 nsew signal output
rlabel metal2 s 208858 241292 208914 242092 6 irq_id_o[2]
port 285 nsew signal output
rlabel metal3 s 0 190408 800 190528 6 irq_id_o[3]
port 286 nsew signal output
rlabel metal3 s 239148 154368 239948 154488 6 irq_id_o[4]
port 287 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 reset
port 288 nsew signal input
rlabel metal4 s 234208 2128 234528 239952 6 VPWR
port 289 nsew power bidirectional
rlabel metal4 s 224208 2128 224528 239952 6 VPWR
port 290 nsew power bidirectional
rlabel metal4 s 214208 2128 214528 239952 6 VPWR
port 291 nsew power bidirectional
rlabel metal4 s 204208 2128 204528 239952 6 VPWR
port 292 nsew power bidirectional
rlabel metal4 s 194208 2128 194528 239952 6 VPWR
port 293 nsew power bidirectional
rlabel metal4 s 184208 2128 184528 239952 6 VPWR
port 294 nsew power bidirectional
rlabel metal4 s 174208 2128 174528 239952 6 VPWR
port 295 nsew power bidirectional
rlabel metal4 s 164208 2128 164528 239952 6 VPWR
port 296 nsew power bidirectional
rlabel metal4 s 154208 2128 154528 239952 6 VPWR
port 297 nsew power bidirectional
rlabel metal4 s 144208 2128 144528 239952 6 VPWR
port 298 nsew power bidirectional
rlabel metal4 s 134208 2128 134528 239952 6 VPWR
port 299 nsew power bidirectional
rlabel metal4 s 124208 2128 124528 239952 6 VPWR
port 300 nsew power bidirectional
rlabel metal4 s 114208 100452 114528 239952 6 VPWR
port 301 nsew power bidirectional
rlabel metal4 s 104208 100452 104528 239952 6 VPWR
port 302 nsew power bidirectional
rlabel metal4 s 94208 100452 94528 239952 6 VPWR
port 303 nsew power bidirectional
rlabel metal4 s 84208 100452 84528 239952 6 VPWR
port 304 nsew power bidirectional
rlabel metal4 s 74208 100452 74528 239952 6 VPWR
port 305 nsew power bidirectional
rlabel metal4 s 64208 100452 64528 239952 6 VPWR
port 306 nsew power bidirectional
rlabel metal4 s 54208 100452 54528 239952 6 VPWR
port 307 nsew power bidirectional
rlabel metal4 s 44208 100452 44528 239952 6 VPWR
port 308 nsew power bidirectional
rlabel metal4 s 34208 100452 34528 239952 6 VPWR
port 309 nsew power bidirectional
rlabel metal4 s 24208 100452 24528 239952 6 VPWR
port 310 nsew power bidirectional
rlabel metal4 s 14208 2128 14528 239952 6 VPWR
port 311 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 239952 6 VPWR
port 312 nsew power bidirectional
rlabel metal4 s 114208 2128 114528 19048 6 VPWR
port 313 nsew power bidirectional
rlabel metal4 s 104208 2128 104528 19048 6 VPWR
port 314 nsew power bidirectional
rlabel metal4 s 94208 2128 94528 19048 6 VPWR
port 315 nsew power bidirectional
rlabel metal4 s 84208 2128 84528 19048 6 VPWR
port 316 nsew power bidirectional
rlabel metal4 s 74208 2128 74528 19048 6 VPWR
port 317 nsew power bidirectional
rlabel metal4 s 64208 2128 64528 19048 6 VPWR
port 318 nsew power bidirectional
rlabel metal4 s 54208 2128 54528 19048 6 VPWR
port 319 nsew power bidirectional
rlabel metal4 s 44208 2128 44528 19048 6 VPWR
port 320 nsew power bidirectional
rlabel metal4 s 34208 2128 34528 19048 6 VPWR
port 321 nsew power bidirectional
rlabel metal4 s 24208 2128 24528 19048 6 VPWR
port 322 nsew power bidirectional
rlabel metal5 s 1104 219750 238832 220070 6 VPWR
port 323 nsew power bidirectional
rlabel metal5 s 1104 189114 238832 189434 6 VPWR
port 324 nsew power bidirectional
rlabel metal5 s 1104 158478 238832 158798 6 VPWR
port 325 nsew power bidirectional
rlabel metal5 s 1104 127842 238832 128162 6 VPWR
port 326 nsew power bidirectional
rlabel metal5 s 1104 97206 238832 97526 6 VPWR
port 327 nsew power bidirectional
rlabel metal5 s 1104 66570 238832 66890 6 VPWR
port 328 nsew power bidirectional
rlabel metal5 s 1104 35934 238832 36254 6 VPWR
port 329 nsew power bidirectional
rlabel metal5 s 1104 5298 238832 5618 6 VPWR
port 330 nsew power bidirectional
rlabel metal4 s 229208 2128 229528 239952 6 VGND
port 331 nsew ground bidirectional
rlabel metal4 s 219208 2128 219528 239952 6 VGND
port 332 nsew ground bidirectional
rlabel metal4 s 209208 2128 209528 239952 6 VGND
port 333 nsew ground bidirectional
rlabel metal4 s 199208 2128 199528 239952 6 VGND
port 334 nsew ground bidirectional
rlabel metal4 s 189208 2128 189528 239952 6 VGND
port 335 nsew ground bidirectional
rlabel metal4 s 179208 2128 179528 239952 6 VGND
port 336 nsew ground bidirectional
rlabel metal4 s 169208 2128 169528 239952 6 VGND
port 337 nsew ground bidirectional
rlabel metal4 s 159208 2128 159528 239952 6 VGND
port 338 nsew ground bidirectional
rlabel metal4 s 149208 2128 149528 239952 6 VGND
port 339 nsew ground bidirectional
rlabel metal4 s 139208 2128 139528 239952 6 VGND
port 340 nsew ground bidirectional
rlabel metal4 s 129208 2128 129528 239952 6 VGND
port 341 nsew ground bidirectional
rlabel metal4 s 119208 2128 119528 239952 6 VGND
port 342 nsew ground bidirectional
rlabel metal4 s 109208 100452 109528 239952 6 VGND
port 343 nsew ground bidirectional
rlabel metal4 s 99208 100452 99528 239952 6 VGND
port 344 nsew ground bidirectional
rlabel metal4 s 89208 100452 89528 239952 6 VGND
port 345 nsew ground bidirectional
rlabel metal4 s 79208 100452 79528 239952 6 VGND
port 346 nsew ground bidirectional
rlabel metal4 s 69208 100452 69528 239952 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 59208 100452 59528 239952 6 VGND
port 348 nsew ground bidirectional
rlabel metal4 s 49208 100452 49528 239952 6 VGND
port 349 nsew ground bidirectional
rlabel metal4 s 39208 100452 39528 239952 6 VGND
port 350 nsew ground bidirectional
rlabel metal4 s 29208 100452 29528 239952 6 VGND
port 351 nsew ground bidirectional
rlabel metal4 s 19208 100452 19528 239952 6 VGND
port 352 nsew ground bidirectional
rlabel metal4 s 9208 2128 9528 239952 6 VGND
port 353 nsew ground bidirectional
rlabel metal4 s 109208 2128 109528 19048 6 VGND
port 354 nsew ground bidirectional
rlabel metal4 s 99208 2128 99528 19048 6 VGND
port 355 nsew ground bidirectional
rlabel metal4 s 89208 2128 89528 19048 6 VGND
port 356 nsew ground bidirectional
rlabel metal4 s 79208 2128 79528 19048 6 VGND
port 357 nsew ground bidirectional
rlabel metal4 s 69208 2128 69528 19048 6 VGND
port 358 nsew ground bidirectional
rlabel metal4 s 59208 2128 59528 19048 6 VGND
port 359 nsew ground bidirectional
rlabel metal4 s 49208 2128 49528 19048 6 VGND
port 360 nsew ground bidirectional
rlabel metal4 s 39208 2128 39528 19048 6 VGND
port 361 nsew ground bidirectional
rlabel metal4 s 29208 2128 29528 19048 6 VGND
port 362 nsew ground bidirectional
rlabel metal4 s 19208 2128 19528 19048 6 VGND
port 363 nsew ground bidirectional
rlabel metal5 s 1104 235068 238832 235388 6 VGND
port 364 nsew ground bidirectional
rlabel metal5 s 1104 204432 238832 204752 6 VGND
port 365 nsew ground bidirectional
rlabel metal5 s 1104 173796 238832 174116 6 VGND
port 366 nsew ground bidirectional
rlabel metal5 s 1104 143160 238832 143480 6 VGND
port 367 nsew ground bidirectional
rlabel metal5 s 1104 112524 238832 112844 6 VGND
port 368 nsew ground bidirectional
rlabel metal5 s 1104 81888 238832 82208 6 VGND
port 369 nsew ground bidirectional
rlabel metal5 s 1104 51252 238832 51572 6 VGND
port 370 nsew ground bidirectional
rlabel metal5 s 1104 20616 238832 20936 6 VGND
port 371 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 239948 242092
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 77548278
string GDS_START 10615672
<< end >>

