magic
tech sky130A
magscale 1 2
timestamp 1624482375
<< obsli1 >>
rect 1104 2159 428812 177361
<< obsm1 >>
rect 474 1300 428812 178084
<< metal2 >>
rect 2778 179200 2834 180000
rect 5538 179200 5594 180000
rect 8298 179200 8354 180000
rect 11058 179200 11114 180000
rect 13818 179200 13874 180000
rect 16578 179200 16634 180000
rect 19338 179200 19394 180000
rect 22098 179200 22154 180000
rect 24858 179200 24914 180000
rect 27618 179200 27674 180000
rect 30378 179200 30434 180000
rect 33138 179200 33194 180000
rect 35898 179200 35954 180000
rect 38198 179200 38254 180000
rect 40958 179200 41014 180000
rect 43718 179200 43774 180000
rect 46478 179200 46534 180000
rect 49238 179200 49294 180000
rect 51998 179200 52054 180000
rect 54758 179200 54814 180000
rect 57518 179200 57574 180000
rect 60278 179200 60334 180000
rect 63038 179200 63094 180000
rect 65798 179200 65854 180000
rect 68558 179200 68614 180000
rect 71318 179200 71374 180000
rect 74078 179200 74134 180000
rect 76838 179200 76894 180000
rect 79598 179200 79654 180000
rect 82358 179200 82414 180000
rect 85118 179200 85174 180000
rect 87878 179200 87934 180000
rect 90638 179200 90694 180000
rect 93398 179200 93454 180000
rect 96158 179200 96214 180000
rect 98918 179200 98974 180000
rect 101678 179200 101734 180000
rect 104438 179200 104494 180000
rect 107198 179200 107254 180000
rect 109958 179200 110014 180000
rect 112718 179200 112774 180000
rect 115018 179200 115074 180000
rect 117778 179200 117834 180000
rect 120538 179200 120594 180000
rect 123298 179200 123354 180000
rect 126058 179200 126114 180000
rect 128818 179200 128874 180000
rect 131578 179200 131634 180000
rect 134338 179200 134394 180000
rect 137098 179200 137154 180000
rect 139858 179200 139914 180000
rect 142618 179200 142674 180000
rect 145378 179200 145434 180000
rect 148138 179200 148194 180000
rect 150898 179200 150954 180000
rect 153658 179200 153714 180000
rect 156418 179200 156474 180000
rect 159178 179200 159234 180000
rect 161938 179200 161994 180000
rect 164698 179200 164754 180000
rect 167458 179200 167514 180000
rect 170218 179200 170274 180000
rect 172978 179200 173034 180000
rect 175738 179200 175794 180000
rect 178498 179200 178554 180000
rect 181258 179200 181314 180000
rect 184018 179200 184074 180000
rect 186778 179200 186834 180000
rect 189538 179200 189594 180000
rect 192298 179200 192354 180000
rect 194598 179200 194654 180000
rect 197358 179200 197414 180000
rect 200118 179200 200174 180000
rect 202878 179200 202934 180000
rect 205638 179200 205694 180000
rect 208398 179200 208454 180000
rect 211158 179200 211214 180000
rect 213918 179200 213974 180000
rect 216678 179200 216734 180000
rect 219438 179200 219494 180000
rect 222198 179200 222254 180000
rect 224958 179200 225014 180000
rect 227718 179200 227774 180000
rect 230478 179200 230534 180000
rect 233238 179200 233294 180000
rect 235998 179200 236054 180000
rect 238758 179200 238814 180000
rect 241518 179200 241574 180000
rect 244278 179200 244334 180000
rect 247038 179200 247094 180000
rect 249798 179200 249854 180000
rect 252558 179200 252614 180000
rect 255318 179200 255374 180000
rect 258078 179200 258134 180000
rect 260838 179200 260894 180000
rect 263598 179200 263654 180000
rect 266358 179200 266414 180000
rect 269118 179200 269174 180000
rect 271878 179200 271934 180000
rect 274178 179200 274234 180000
rect 276938 179200 276994 180000
rect 279698 179200 279754 180000
rect 282458 179200 282514 180000
rect 285218 179200 285274 180000
rect 287978 179200 288034 180000
rect 290738 179200 290794 180000
rect 293498 179200 293554 180000
rect 296258 179200 296314 180000
rect 299018 179200 299074 180000
rect 301778 179200 301834 180000
rect 304538 179200 304594 180000
rect 307298 179200 307354 180000
rect 310058 179200 310114 180000
rect 312818 179200 312874 180000
rect 315578 179200 315634 180000
rect 318338 179200 318394 180000
rect 321098 179200 321154 180000
rect 323858 179200 323914 180000
rect 326618 179200 326674 180000
rect 329378 179200 329434 180000
rect 332138 179200 332194 180000
rect 334898 179200 334954 180000
rect 337658 179200 337714 180000
rect 340418 179200 340474 180000
rect 343178 179200 343234 180000
rect 345938 179200 345994 180000
rect 348698 179200 348754 180000
rect 350998 179200 351054 180000
rect 353758 179200 353814 180000
rect 356518 179200 356574 180000
rect 359278 179200 359334 180000
rect 362038 179200 362094 180000
rect 364798 179200 364854 180000
rect 367558 179200 367614 180000
rect 370318 179200 370374 180000
rect 373078 179200 373134 180000
rect 375838 179200 375894 180000
rect 378598 179200 378654 180000
rect 381358 179200 381414 180000
rect 384118 179200 384174 180000
rect 386878 179200 386934 180000
rect 389638 179200 389694 180000
rect 392398 179200 392454 180000
rect 395158 179200 395214 180000
rect 397918 179200 397974 180000
rect 400678 179200 400734 180000
rect 403438 179200 403494 180000
rect 406198 179200 406254 180000
rect 408958 179200 409014 180000
rect 411718 179200 411774 180000
rect 414478 179200 414534 180000
rect 417238 179200 417294 180000
rect 419998 179200 420054 180000
rect 422758 179200 422814 180000
rect 425518 179200 425574 180000
rect 428278 179200 428334 180000
rect 478 0 534 800
rect 2778 0 2834 800
rect 5538 0 5594 800
rect 8298 0 8354 800
rect 11058 0 11114 800
rect 13818 0 13874 800
rect 16578 0 16634 800
rect 19338 0 19394 800
rect 22098 0 22154 800
rect 24858 0 24914 800
rect 27618 0 27674 800
rect 30378 0 30434 800
rect 33138 0 33194 800
rect 35898 0 35954 800
rect 38658 0 38714 800
rect 41418 0 41474 800
rect 44178 0 44234 800
rect 46938 0 46994 800
rect 49698 0 49754 800
rect 52458 0 52514 800
rect 55218 0 55274 800
rect 57978 0 58034 800
rect 60738 0 60794 800
rect 63498 0 63554 800
rect 66258 0 66314 800
rect 69018 0 69074 800
rect 71778 0 71834 800
rect 74538 0 74594 800
rect 77298 0 77354 800
rect 79598 0 79654 800
rect 82358 0 82414 800
rect 85118 0 85174 800
rect 87878 0 87934 800
rect 90638 0 90694 800
rect 93398 0 93454 800
rect 96158 0 96214 800
rect 98918 0 98974 800
rect 101678 0 101734 800
rect 104438 0 104494 800
rect 107198 0 107254 800
rect 109958 0 110014 800
rect 112718 0 112774 800
rect 115478 0 115534 800
rect 118238 0 118294 800
rect 120998 0 121054 800
rect 123758 0 123814 800
rect 126518 0 126574 800
rect 129278 0 129334 800
rect 132038 0 132094 800
rect 134798 0 134854 800
rect 137558 0 137614 800
rect 140318 0 140374 800
rect 143078 0 143134 800
rect 145838 0 145894 800
rect 148598 0 148654 800
rect 151358 0 151414 800
rect 154118 0 154174 800
rect 156878 0 156934 800
rect 159178 0 159234 800
rect 161938 0 161994 800
rect 164698 0 164754 800
rect 167458 0 167514 800
rect 170218 0 170274 800
rect 172978 0 173034 800
rect 175738 0 175794 800
rect 178498 0 178554 800
rect 181258 0 181314 800
rect 184018 0 184074 800
rect 186778 0 186834 800
rect 189538 0 189594 800
rect 192298 0 192354 800
rect 195058 0 195114 800
rect 197818 0 197874 800
rect 200578 0 200634 800
rect 203338 0 203394 800
rect 206098 0 206154 800
rect 208858 0 208914 800
rect 211618 0 211674 800
rect 214378 0 214434 800
rect 217138 0 217194 800
rect 219898 0 219954 800
rect 222658 0 222714 800
rect 225418 0 225474 800
rect 228178 0 228234 800
rect 230938 0 230994 800
rect 233698 0 233754 800
rect 235998 0 236054 800
rect 238758 0 238814 800
rect 241518 0 241574 800
rect 244278 0 244334 800
rect 247038 0 247094 800
rect 249798 0 249854 800
rect 252558 0 252614 800
rect 255318 0 255374 800
rect 258078 0 258134 800
rect 260838 0 260894 800
rect 263598 0 263654 800
rect 266358 0 266414 800
rect 269118 0 269174 800
rect 271878 0 271934 800
rect 274638 0 274694 800
rect 277398 0 277454 800
rect 280158 0 280214 800
rect 282918 0 282974 800
rect 285678 0 285734 800
rect 288438 0 288494 800
rect 291198 0 291254 800
rect 293958 0 294014 800
rect 296718 0 296774 800
rect 299478 0 299534 800
rect 302238 0 302294 800
rect 304998 0 305054 800
rect 307758 0 307814 800
rect 310518 0 310574 800
rect 313278 0 313334 800
rect 315578 0 315634 800
rect 318338 0 318394 800
rect 321098 0 321154 800
rect 323858 0 323914 800
rect 326618 0 326674 800
rect 329378 0 329434 800
rect 332138 0 332194 800
rect 334898 0 334954 800
rect 337658 0 337714 800
rect 340418 0 340474 800
rect 343178 0 343234 800
rect 345938 0 345994 800
rect 348698 0 348754 800
rect 351458 0 351514 800
rect 354218 0 354274 800
rect 356978 0 357034 800
rect 359738 0 359794 800
rect 362498 0 362554 800
rect 365258 0 365314 800
rect 368018 0 368074 800
rect 370778 0 370834 800
rect 373538 0 373594 800
rect 376298 0 376354 800
rect 379058 0 379114 800
rect 381818 0 381874 800
rect 384578 0 384634 800
rect 387338 0 387394 800
rect 390098 0 390154 800
rect 392858 0 392914 800
rect 395158 0 395214 800
rect 397918 0 397974 800
rect 400678 0 400734 800
rect 403438 0 403494 800
rect 406198 0 406254 800
rect 408958 0 409014 800
rect 411718 0 411774 800
rect 414478 0 414534 800
rect 417238 0 417294 800
rect 419998 0 420054 800
rect 422758 0 422814 800
rect 425518 0 425574 800
rect 428278 0 428334 800
<< obsm2 >>
rect 480 179144 2722 179200
rect 2890 179144 5482 179200
rect 5650 179144 8242 179200
rect 8410 179144 11002 179200
rect 11170 179144 13762 179200
rect 13930 179144 16522 179200
rect 16690 179144 19282 179200
rect 19450 179144 22042 179200
rect 22210 179144 24802 179200
rect 24970 179144 27562 179200
rect 27730 179144 30322 179200
rect 30490 179144 33082 179200
rect 33250 179144 35842 179200
rect 36010 179144 38142 179200
rect 38310 179144 40902 179200
rect 41070 179144 43662 179200
rect 43830 179144 46422 179200
rect 46590 179144 49182 179200
rect 49350 179144 51942 179200
rect 52110 179144 54702 179200
rect 54870 179144 57462 179200
rect 57630 179144 60222 179200
rect 60390 179144 62982 179200
rect 63150 179144 65742 179200
rect 65910 179144 68502 179200
rect 68670 179144 71262 179200
rect 71430 179144 74022 179200
rect 74190 179144 76782 179200
rect 76950 179144 79542 179200
rect 79710 179144 82302 179200
rect 82470 179144 85062 179200
rect 85230 179144 87822 179200
rect 87990 179144 90582 179200
rect 90750 179144 93342 179200
rect 93510 179144 96102 179200
rect 96270 179144 98862 179200
rect 99030 179144 101622 179200
rect 101790 179144 104382 179200
rect 104550 179144 107142 179200
rect 107310 179144 109902 179200
rect 110070 179144 112662 179200
rect 112830 179144 114962 179200
rect 115130 179144 117722 179200
rect 117890 179144 120482 179200
rect 120650 179144 123242 179200
rect 123410 179144 126002 179200
rect 126170 179144 128762 179200
rect 128930 179144 131522 179200
rect 131690 179144 134282 179200
rect 134450 179144 137042 179200
rect 137210 179144 139802 179200
rect 139970 179144 142562 179200
rect 142730 179144 145322 179200
rect 145490 179144 148082 179200
rect 148250 179144 150842 179200
rect 151010 179144 153602 179200
rect 153770 179144 156362 179200
rect 156530 179144 159122 179200
rect 159290 179144 161882 179200
rect 162050 179144 164642 179200
rect 164810 179144 167402 179200
rect 167570 179144 170162 179200
rect 170330 179144 172922 179200
rect 173090 179144 175682 179200
rect 175850 179144 178442 179200
rect 178610 179144 181202 179200
rect 181370 179144 183962 179200
rect 184130 179144 186722 179200
rect 186890 179144 189482 179200
rect 189650 179144 192242 179200
rect 192410 179144 194542 179200
rect 194710 179144 197302 179200
rect 197470 179144 200062 179200
rect 200230 179144 202822 179200
rect 202990 179144 205582 179200
rect 205750 179144 208342 179200
rect 208510 179144 211102 179200
rect 211270 179144 213862 179200
rect 214030 179144 216622 179200
rect 216790 179144 219382 179200
rect 219550 179144 222142 179200
rect 222310 179144 224902 179200
rect 225070 179144 227662 179200
rect 227830 179144 230422 179200
rect 230590 179144 233182 179200
rect 233350 179144 235942 179200
rect 236110 179144 238702 179200
rect 238870 179144 241462 179200
rect 241630 179144 244222 179200
rect 244390 179144 246982 179200
rect 247150 179144 249742 179200
rect 249910 179144 252502 179200
rect 252670 179144 255262 179200
rect 255430 179144 258022 179200
rect 258190 179144 260782 179200
rect 260950 179144 263542 179200
rect 263710 179144 266302 179200
rect 266470 179144 269062 179200
rect 269230 179144 271822 179200
rect 271990 179144 274122 179200
rect 274290 179144 276882 179200
rect 277050 179144 279642 179200
rect 279810 179144 282402 179200
rect 282570 179144 285162 179200
rect 285330 179144 287922 179200
rect 288090 179144 290682 179200
rect 290850 179144 293442 179200
rect 293610 179144 296202 179200
rect 296370 179144 298962 179200
rect 299130 179144 301722 179200
rect 301890 179144 304482 179200
rect 304650 179144 307242 179200
rect 307410 179144 310002 179200
rect 310170 179144 312762 179200
rect 312930 179144 315522 179200
rect 315690 179144 318282 179200
rect 318450 179144 321042 179200
rect 321210 179144 323802 179200
rect 323970 179144 326562 179200
rect 326730 179144 329322 179200
rect 329490 179144 332082 179200
rect 332250 179144 334842 179200
rect 335010 179144 337602 179200
rect 337770 179144 340362 179200
rect 340530 179144 343122 179200
rect 343290 179144 345882 179200
rect 346050 179144 348642 179200
rect 348810 179144 350942 179200
rect 351110 179144 353702 179200
rect 353870 179144 356462 179200
rect 356630 179144 359222 179200
rect 359390 179144 361982 179200
rect 362150 179144 364742 179200
rect 364910 179144 367502 179200
rect 367670 179144 370262 179200
rect 370430 179144 373022 179200
rect 373190 179144 375782 179200
rect 375950 179144 378542 179200
rect 378710 179144 381302 179200
rect 381470 179144 384062 179200
rect 384230 179144 386822 179200
rect 386990 179144 389582 179200
rect 389750 179144 392342 179200
rect 392510 179144 395102 179200
rect 395270 179144 397862 179200
rect 398030 179144 400622 179200
rect 400790 179144 403382 179200
rect 403550 179144 406142 179200
rect 406310 179144 408902 179200
rect 409070 179144 411662 179200
rect 411830 179144 414422 179200
rect 414590 179144 417182 179200
rect 417350 179144 419942 179200
rect 420110 179144 422702 179200
rect 422870 179144 425462 179200
rect 425630 179144 428222 179200
rect 480 856 428332 179144
rect 590 800 2722 856
rect 2890 800 5482 856
rect 5650 800 8242 856
rect 8410 800 11002 856
rect 11170 800 13762 856
rect 13930 800 16522 856
rect 16690 800 19282 856
rect 19450 800 22042 856
rect 22210 800 24802 856
rect 24970 800 27562 856
rect 27730 800 30322 856
rect 30490 800 33082 856
rect 33250 800 35842 856
rect 36010 800 38602 856
rect 38770 800 41362 856
rect 41530 800 44122 856
rect 44290 800 46882 856
rect 47050 800 49642 856
rect 49810 800 52402 856
rect 52570 800 55162 856
rect 55330 800 57922 856
rect 58090 800 60682 856
rect 60850 800 63442 856
rect 63610 800 66202 856
rect 66370 800 68962 856
rect 69130 800 71722 856
rect 71890 800 74482 856
rect 74650 800 77242 856
rect 77410 800 79542 856
rect 79710 800 82302 856
rect 82470 800 85062 856
rect 85230 800 87822 856
rect 87990 800 90582 856
rect 90750 800 93342 856
rect 93510 800 96102 856
rect 96270 800 98862 856
rect 99030 800 101622 856
rect 101790 800 104382 856
rect 104550 800 107142 856
rect 107310 800 109902 856
rect 110070 800 112662 856
rect 112830 800 115422 856
rect 115590 800 118182 856
rect 118350 800 120942 856
rect 121110 800 123702 856
rect 123870 800 126462 856
rect 126630 800 129222 856
rect 129390 800 131982 856
rect 132150 800 134742 856
rect 134910 800 137502 856
rect 137670 800 140262 856
rect 140430 800 143022 856
rect 143190 800 145782 856
rect 145950 800 148542 856
rect 148710 800 151302 856
rect 151470 800 154062 856
rect 154230 800 156822 856
rect 156990 800 159122 856
rect 159290 800 161882 856
rect 162050 800 164642 856
rect 164810 800 167402 856
rect 167570 800 170162 856
rect 170330 800 172922 856
rect 173090 800 175682 856
rect 175850 800 178442 856
rect 178610 800 181202 856
rect 181370 800 183962 856
rect 184130 800 186722 856
rect 186890 800 189482 856
rect 189650 800 192242 856
rect 192410 800 195002 856
rect 195170 800 197762 856
rect 197930 800 200522 856
rect 200690 800 203282 856
rect 203450 800 206042 856
rect 206210 800 208802 856
rect 208970 800 211562 856
rect 211730 800 214322 856
rect 214490 800 217082 856
rect 217250 800 219842 856
rect 220010 800 222602 856
rect 222770 800 225362 856
rect 225530 800 228122 856
rect 228290 800 230882 856
rect 231050 800 233642 856
rect 233810 800 235942 856
rect 236110 800 238702 856
rect 238870 800 241462 856
rect 241630 800 244222 856
rect 244390 800 246982 856
rect 247150 800 249742 856
rect 249910 800 252502 856
rect 252670 800 255262 856
rect 255430 800 258022 856
rect 258190 800 260782 856
rect 260950 800 263542 856
rect 263710 800 266302 856
rect 266470 800 269062 856
rect 269230 800 271822 856
rect 271990 800 274582 856
rect 274750 800 277342 856
rect 277510 800 280102 856
rect 280270 800 282862 856
rect 283030 800 285622 856
rect 285790 800 288382 856
rect 288550 800 291142 856
rect 291310 800 293902 856
rect 294070 800 296662 856
rect 296830 800 299422 856
rect 299590 800 302182 856
rect 302350 800 304942 856
rect 305110 800 307702 856
rect 307870 800 310462 856
rect 310630 800 313222 856
rect 313390 800 315522 856
rect 315690 800 318282 856
rect 318450 800 321042 856
rect 321210 800 323802 856
rect 323970 800 326562 856
rect 326730 800 329322 856
rect 329490 800 332082 856
rect 332250 800 334842 856
rect 335010 800 337602 856
rect 337770 800 340362 856
rect 340530 800 343122 856
rect 343290 800 345882 856
rect 346050 800 348642 856
rect 348810 800 351402 856
rect 351570 800 354162 856
rect 354330 800 356922 856
rect 357090 800 359682 856
rect 359850 800 362442 856
rect 362610 800 365202 856
rect 365370 800 367962 856
rect 368130 800 370722 856
rect 370890 800 373482 856
rect 373650 800 376242 856
rect 376410 800 379002 856
rect 379170 800 381762 856
rect 381930 800 384522 856
rect 384690 800 387282 856
rect 387450 800 390042 856
rect 390210 800 392802 856
rect 392970 800 395102 856
rect 395270 800 397862 856
rect 398030 800 400622 856
rect 400790 800 403382 856
rect 403550 800 406142 856
rect 406310 800 408902 856
rect 409070 800 411662 856
rect 411830 800 414422 856
rect 414590 800 417182 856
rect 417350 800 419942 856
rect 420110 800 422702 856
rect 422870 800 425462 856
rect 425630 800 428222 856
<< metal3 >>
rect 0 178848 800 178968
rect 429200 177488 430000 177608
rect 0 174768 800 174888
rect 429200 173408 430000 173528
rect 0 170688 800 170808
rect 429200 169328 430000 169448
rect 0 166608 800 166728
rect 429200 165248 430000 165368
rect 0 162528 800 162648
rect 429200 161168 430000 161288
rect 0 158448 800 158568
rect 429200 157088 430000 157208
rect 0 154368 800 154488
rect 429200 153008 430000 153128
rect 0 150288 800 150408
rect 429200 148928 430000 149048
rect 0 146208 800 146328
rect 429200 144848 430000 144968
rect 0 142128 800 142248
rect 429200 140768 430000 140888
rect 0 138048 800 138168
rect 429200 136688 430000 136808
rect 0 133968 800 134088
rect 429200 132608 430000 132728
rect 0 129888 800 130008
rect 429200 128528 430000 128648
rect 0 125808 800 125928
rect 429200 124448 430000 124568
rect 0 121728 800 121848
rect 429200 120368 430000 120488
rect 0 117648 800 117768
rect 429200 116288 430000 116408
rect 0 114248 800 114368
rect 429200 112208 430000 112328
rect 0 110168 800 110288
rect 429200 108128 430000 108248
rect 0 106088 800 106208
rect 429200 104048 430000 104168
rect 0 102008 800 102128
rect 429200 99968 430000 100088
rect 0 97928 800 98048
rect 429200 95888 430000 96008
rect 0 93848 800 93968
rect 429200 91808 430000 91928
rect 0 89768 800 89888
rect 429200 87728 430000 87848
rect 0 85688 800 85808
rect 429200 83648 430000 83768
rect 0 81608 800 81728
rect 429200 79568 430000 79688
rect 0 77528 800 77648
rect 429200 75488 430000 75608
rect 0 73448 800 73568
rect 429200 71408 430000 71528
rect 0 69368 800 69488
rect 429200 67328 430000 67448
rect 0 65288 800 65408
rect 429200 63248 430000 63368
rect 0 61208 800 61328
rect 429200 59848 430000 59968
rect 0 57128 800 57248
rect 429200 55768 430000 55888
rect 0 53048 800 53168
rect 429200 51688 430000 51808
rect 0 48968 800 49088
rect 429200 47608 430000 47728
rect 0 44888 800 45008
rect 429200 43528 430000 43648
rect 0 40808 800 40928
rect 429200 39448 430000 39568
rect 0 36728 800 36848
rect 429200 35368 430000 35488
rect 0 32648 800 32768
rect 429200 31288 430000 31408
rect 0 28568 800 28688
rect 429200 27208 430000 27328
rect 0 24488 800 24608
rect 429200 23128 430000 23248
rect 0 20408 800 20528
rect 429200 19048 430000 19168
rect 0 16328 800 16448
rect 429200 14968 430000 15088
rect 0 12248 800 12368
rect 429200 10888 430000 11008
rect 0 8168 800 8288
rect 429200 6808 430000 6928
rect 0 4088 800 4208
rect 429200 2728 430000 2848
<< obsm3 >>
rect 880 178768 429200 178941
rect 800 177688 429200 178768
rect 800 177408 429120 177688
rect 800 174968 429200 177408
rect 880 174688 429200 174968
rect 800 173608 429200 174688
rect 800 173328 429120 173608
rect 800 170888 429200 173328
rect 880 170608 429200 170888
rect 800 169528 429200 170608
rect 800 169248 429120 169528
rect 800 166808 429200 169248
rect 880 166528 429200 166808
rect 800 165448 429200 166528
rect 800 165168 429120 165448
rect 800 162728 429200 165168
rect 880 162448 429200 162728
rect 800 161368 429200 162448
rect 800 161088 429120 161368
rect 800 158648 429200 161088
rect 880 158368 429200 158648
rect 800 157288 429200 158368
rect 800 157008 429120 157288
rect 800 154568 429200 157008
rect 880 154288 429200 154568
rect 800 153208 429200 154288
rect 800 152928 429120 153208
rect 800 150488 429200 152928
rect 880 150208 429200 150488
rect 800 149128 429200 150208
rect 800 148848 429120 149128
rect 800 146408 429200 148848
rect 880 146128 429200 146408
rect 800 145048 429200 146128
rect 800 144768 429120 145048
rect 800 142328 429200 144768
rect 880 142048 429200 142328
rect 800 140968 429200 142048
rect 800 140688 429120 140968
rect 800 138248 429200 140688
rect 880 137968 429200 138248
rect 800 136888 429200 137968
rect 800 136608 429120 136888
rect 800 134168 429200 136608
rect 880 133888 429200 134168
rect 800 132808 429200 133888
rect 800 132528 429120 132808
rect 800 130088 429200 132528
rect 880 129808 429200 130088
rect 800 128728 429200 129808
rect 800 128448 429120 128728
rect 800 126008 429200 128448
rect 880 125728 429200 126008
rect 800 124648 429200 125728
rect 800 124368 429120 124648
rect 800 121928 429200 124368
rect 880 121648 429200 121928
rect 800 120568 429200 121648
rect 800 120288 429120 120568
rect 800 117848 429200 120288
rect 880 117568 429200 117848
rect 800 116488 429200 117568
rect 800 116208 429120 116488
rect 800 114448 429200 116208
rect 880 114168 429200 114448
rect 800 112408 429200 114168
rect 800 112128 429120 112408
rect 800 110368 429200 112128
rect 880 110088 429200 110368
rect 800 108328 429200 110088
rect 800 108048 429120 108328
rect 800 106288 429200 108048
rect 880 106008 429200 106288
rect 800 104248 429200 106008
rect 800 103968 429120 104248
rect 800 102208 429200 103968
rect 880 101928 429200 102208
rect 800 100168 429200 101928
rect 800 99888 429120 100168
rect 800 98128 429200 99888
rect 880 97848 429200 98128
rect 800 96088 429200 97848
rect 800 95808 429120 96088
rect 800 94048 429200 95808
rect 880 93768 429200 94048
rect 800 92008 429200 93768
rect 800 91728 429120 92008
rect 800 89968 429200 91728
rect 880 89688 429200 89968
rect 800 87928 429200 89688
rect 800 87648 429120 87928
rect 800 85888 429200 87648
rect 880 85608 429200 85888
rect 800 83848 429200 85608
rect 800 83568 429120 83848
rect 800 81808 429200 83568
rect 880 81528 429200 81808
rect 800 79768 429200 81528
rect 800 79488 429120 79768
rect 800 77728 429200 79488
rect 880 77448 429200 77728
rect 800 75688 429200 77448
rect 800 75408 429120 75688
rect 800 73648 429200 75408
rect 880 73368 429200 73648
rect 800 71608 429200 73368
rect 800 71328 429120 71608
rect 800 69568 429200 71328
rect 880 69288 429200 69568
rect 800 67528 429200 69288
rect 800 67248 429120 67528
rect 800 65488 429200 67248
rect 880 65208 429200 65488
rect 800 63448 429200 65208
rect 800 63168 429120 63448
rect 800 61408 429200 63168
rect 880 61128 429200 61408
rect 800 60048 429200 61128
rect 800 59768 429120 60048
rect 800 57328 429200 59768
rect 880 57048 429200 57328
rect 800 55968 429200 57048
rect 800 55688 429120 55968
rect 800 53248 429200 55688
rect 880 52968 429200 53248
rect 800 51888 429200 52968
rect 800 51608 429120 51888
rect 800 49168 429200 51608
rect 880 48888 429200 49168
rect 800 47808 429200 48888
rect 800 47528 429120 47808
rect 800 45088 429200 47528
rect 880 44808 429200 45088
rect 800 43728 429200 44808
rect 800 43448 429120 43728
rect 800 41008 429200 43448
rect 880 40728 429200 41008
rect 800 39648 429200 40728
rect 800 39368 429120 39648
rect 800 36928 429200 39368
rect 880 36648 429200 36928
rect 800 35568 429200 36648
rect 800 35288 429120 35568
rect 800 32848 429200 35288
rect 880 32568 429200 32848
rect 800 31488 429200 32568
rect 800 31208 429120 31488
rect 800 28768 429200 31208
rect 880 28488 429200 28768
rect 800 27408 429200 28488
rect 800 27128 429120 27408
rect 800 24688 429200 27128
rect 880 24408 429200 24688
rect 800 23328 429200 24408
rect 800 23048 429120 23328
rect 800 20608 429200 23048
rect 880 20328 429200 20608
rect 800 19248 429200 20328
rect 800 18968 429120 19248
rect 800 16528 429200 18968
rect 880 16248 429200 16528
rect 800 15168 429200 16248
rect 800 14888 429120 15168
rect 800 12448 429200 14888
rect 880 12168 429200 12448
rect 800 11088 429200 12168
rect 800 10808 429120 11088
rect 800 8368 429200 10808
rect 880 8088 429200 8368
rect 800 7008 429200 8088
rect 800 6728 429120 7008
rect 800 4288 429200 6728
rect 880 4008 429200 4288
rect 800 2928 429200 4008
rect 800 2648 429120 2928
rect 800 1939 429200 2648
<< metal4 >>
rect 4208 2128 4528 177392
rect 19568 2128 19888 177392
rect 34928 2128 35248 177392
rect 50288 2128 50608 177392
rect 65648 2128 65968 177392
rect 81008 2128 81328 177392
rect 96368 2128 96688 177392
rect 111728 2128 112048 177392
rect 127088 2128 127408 177392
rect 142448 2128 142768 177392
rect 157808 2128 158128 177392
rect 173168 2128 173488 177392
rect 188528 2128 188848 177392
rect 203888 2128 204208 177392
rect 219248 2128 219568 177392
rect 234608 2128 234928 177392
rect 249968 2128 250288 177392
rect 265328 2128 265648 177392
rect 280688 2128 281008 177392
rect 296048 2128 296368 177392
rect 311408 2128 311728 177392
rect 326768 2128 327088 177392
rect 342128 2128 342448 177392
rect 357488 2128 357808 177392
rect 372848 2128 373168 177392
rect 388208 2128 388528 177392
rect 403568 2128 403888 177392
rect 418928 2128 419248 177392
<< obsm4 >>
rect 18091 2048 19488 177173
rect 19968 2048 34848 177173
rect 35328 2048 50208 177173
rect 50688 2048 65568 177173
rect 66048 2048 80928 177173
rect 81408 2048 96288 177173
rect 96768 2048 111648 177173
rect 112128 2048 127008 177173
rect 127488 2048 142368 177173
rect 142848 2048 157728 177173
rect 158208 2048 173088 177173
rect 173568 2048 188448 177173
rect 188928 2048 203808 177173
rect 204288 2048 219168 177173
rect 219648 2048 234528 177173
rect 235008 2048 249888 177173
rect 250368 2048 265248 177173
rect 265728 2048 280608 177173
rect 281088 2048 295968 177173
rect 296448 2048 311328 177173
rect 311808 2048 326688 177173
rect 327168 2048 342048 177173
rect 342528 2048 357408 177173
rect 357888 2048 372768 177173
rect 373248 2048 387997 177173
rect 18091 1939 387997 2048
<< metal5 >>
rect 1104 173796 428812 174116
rect 1104 158478 428812 158798
rect 1104 143160 428812 143480
rect 1104 127842 428812 128162
rect 1104 112524 428812 112844
rect 1104 97206 428812 97526
rect 1104 81888 428812 82208
rect 1104 66570 428812 66890
rect 1104 51252 428812 51572
rect 1104 35934 428812 36254
rect 1104 20616 428812 20936
rect 1104 5298 428812 5618
<< obsm5 >>
rect 45932 113164 359604 126300
rect 45932 97846 359604 112204
rect 45932 82528 359604 96886
rect 45932 67210 359604 81568
rect 45932 60700 359604 66250
<< labels >>
rlabel metal2 s 375838 179200 375894 180000 6 boot_addr_i[0]
port 1 nsew signal input
rlabel metal2 s 186778 179200 186834 180000 6 boot_addr_i[10]
port 2 nsew signal input
rlabel metal2 s 403438 0 403494 800 6 boot_addr_i[11]
port 3 nsew signal input
rlabel metal2 s 123298 179200 123354 180000 6 boot_addr_i[12]
port 4 nsew signal input
rlabel metal2 s 181258 179200 181314 180000 6 boot_addr_i[13]
port 5 nsew signal input
rlabel metal3 s 429200 51688 430000 51808 6 boot_addr_i[14]
port 6 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 boot_addr_i[15]
port 7 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 boot_addr_i[16]
port 8 nsew signal input
rlabel metal2 s 354218 0 354274 800 6 boot_addr_i[17]
port 9 nsew signal input
rlabel metal2 s 280158 0 280214 800 6 boot_addr_i[18]
port 10 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 boot_addr_i[19]
port 11 nsew signal input
rlabel metal3 s 429200 87728 430000 87848 6 boot_addr_i[1]
port 12 nsew signal input
rlabel metal3 s 429200 153008 430000 153128 6 boot_addr_i[20]
port 13 nsew signal input
rlabel metal2 s 307758 0 307814 800 6 boot_addr_i[21]
port 14 nsew signal input
rlabel metal2 s 315578 179200 315634 180000 6 boot_addr_i[22]
port 15 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 boot_addr_i[23]
port 16 nsew signal input
rlabel metal2 s 318338 0 318394 800 6 boot_addr_i[24]
port 17 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 boot_addr_i[25]
port 18 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 boot_addr_i[26]
port 19 nsew signal input
rlabel metal3 s 0 174768 800 174888 6 boot_addr_i[27]
port 20 nsew signal input
rlabel metal2 s 230478 179200 230534 180000 6 boot_addr_i[28]
port 21 nsew signal input
rlabel metal2 s 65798 179200 65854 180000 6 boot_addr_i[29]
port 22 nsew signal input
rlabel metal2 s 131578 179200 131634 180000 6 boot_addr_i[2]
port 23 nsew signal input
rlabel metal2 s 329378 0 329434 800 6 boot_addr_i[30]
port 24 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 boot_addr_i[31]
port 25 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 boot_addr_i[3]
port 26 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 boot_addr_i[4]
port 27 nsew signal input
rlabel metal2 s 8298 179200 8354 180000 6 boot_addr_i[5]
port 28 nsew signal input
rlabel metal2 s 276938 179200 276994 180000 6 boot_addr_i[6]
port 29 nsew signal input
rlabel metal3 s 429200 59848 430000 59968 6 boot_addr_i[7]
port 30 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 boot_addr_i[8]
port 31 nsew signal input
rlabel metal2 s 71318 179200 71374 180000 6 boot_addr_i[9]
port 32 nsew signal input
rlabel metal2 s 178498 179200 178554 180000 6 clk_i
port 33 nsew signal input
rlabel metal3 s 429200 39448 430000 39568 6 cluster_id_i[0]
port 34 nsew signal input
rlabel metal2 s 386878 179200 386934 180000 6 cluster_id_i[1]
port 35 nsew signal input
rlabel metal2 s 414478 0 414534 800 6 cluster_id_i[2]
port 36 nsew signal input
rlabel metal2 s 109958 179200 110014 180000 6 cluster_id_i[3]
port 37 nsew signal input
rlabel metal2 s 252558 179200 252614 180000 6 cluster_id_i[4]
port 38 nsew signal input
rlabel metal2 s 51998 179200 52054 180000 6 cluster_id_i[5]
port 39 nsew signal input
rlabel metal3 s 429200 140768 430000 140888 6 core_id_i[0]
port 40 nsew signal input
rlabel metal2 s 186778 0 186834 800 6 core_id_i[1]
port 41 nsew signal input
rlabel metal2 s 293958 0 294014 800 6 core_id_i[2]
port 42 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 core_id_i[3]
port 43 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 data_addr_o[0]
port 44 nsew signal output
rlabel metal2 s 235998 179200 236054 180000 6 data_addr_o[10]
port 45 nsew signal output
rlabel metal2 s 350998 179200 351054 180000 6 data_addr_o[11]
port 46 nsew signal output
rlabel metal2 s 293498 179200 293554 180000 6 data_addr_o[12]
port 47 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 data_addr_o[13]
port 48 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 data_addr_o[14]
port 49 nsew signal output
rlabel metal2 s 150898 179200 150954 180000 6 data_addr_o[15]
port 50 nsew signal output
rlabel metal2 s 230938 0 230994 800 6 data_addr_o[16]
port 51 nsew signal output
rlabel metal2 s 19338 179200 19394 180000 6 data_addr_o[17]
port 52 nsew signal output
rlabel metal3 s 429200 177488 430000 177608 6 data_addr_o[18]
port 53 nsew signal output
rlabel metal3 s 429200 161168 430000 161288 6 data_addr_o[19]
port 54 nsew signal output
rlabel metal2 s 406198 0 406254 800 6 data_addr_o[1]
port 55 nsew signal output
rlabel metal2 s 392858 0 392914 800 6 data_addr_o[20]
port 56 nsew signal output
rlabel metal2 s 197358 179200 197414 180000 6 data_addr_o[21]
port 57 nsew signal output
rlabel metal3 s 429200 116288 430000 116408 6 data_addr_o[22]
port 58 nsew signal output
rlabel metal2 s 170218 179200 170274 180000 6 data_addr_o[23]
port 59 nsew signal output
rlabel metal2 s 356978 0 357034 800 6 data_addr_o[24]
port 60 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 data_addr_o[25]
port 61 nsew signal output
rlabel metal2 s 345938 0 345994 800 6 data_addr_o[26]
port 62 nsew signal output
rlabel metal2 s 403438 179200 403494 180000 6 data_addr_o[27]
port 63 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 data_addr_o[28]
port 64 nsew signal output
rlabel metal2 s 282918 0 282974 800 6 data_addr_o[29]
port 65 nsew signal output
rlabel metal2 s 74078 179200 74134 180000 6 data_addr_o[2]
port 66 nsew signal output
rlabel metal2 s 145378 179200 145434 180000 6 data_addr_o[30]
port 67 nsew signal output
rlabel metal2 s 310518 0 310574 800 6 data_addr_o[31]
port 68 nsew signal output
rlabel metal3 s 429200 75488 430000 75608 6 data_addr_o[3]
port 69 nsew signal output
rlabel metal3 s 429200 2728 430000 2848 6 data_addr_o[4]
port 70 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 data_addr_o[5]
port 71 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 data_addr_o[6]
port 72 nsew signal output
rlabel metal2 s 258078 179200 258134 180000 6 data_addr_o[7]
port 73 nsew signal output
rlabel metal2 s 40958 179200 41014 180000 6 data_addr_o[8]
port 74 nsew signal output
rlabel metal2 s 381358 179200 381414 180000 6 data_addr_o[9]
port 75 nsew signal output
rlabel metal2 s 109958 0 110014 800 6 data_be_o[0]
port 76 nsew signal output
rlabel metal2 s 63038 179200 63094 180000 6 data_be_o[1]
port 77 nsew signal output
rlabel metal2 s 329378 179200 329434 180000 6 data_be_o[2]
port 78 nsew signal output
rlabel metal2 s 381818 0 381874 800 6 data_be_o[3]
port 79 nsew signal output
rlabel metal2 s 247038 179200 247094 180000 6 data_err_i
port 80 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 data_gnt_i
port 81 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 data_rdata_i[0]
port 82 nsew signal input
rlabel metal3 s 429200 35368 430000 35488 6 data_rdata_i[10]
port 83 nsew signal input
rlabel metal2 s 400678 179200 400734 180000 6 data_rdata_i[11]
port 84 nsew signal input
rlabel metal2 s 192298 179200 192354 180000 6 data_rdata_i[12]
port 85 nsew signal input
rlabel metal2 s 351458 0 351514 800 6 data_rdata_i[13]
port 86 nsew signal input
rlabel metal3 s 429200 6808 430000 6928 6 data_rdata_i[14]
port 87 nsew signal input
rlabel metal2 s 222198 179200 222254 180000 6 data_rdata_i[15]
port 88 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 data_rdata_i[16]
port 89 nsew signal input
rlabel metal2 s 249798 0 249854 800 6 data_rdata_i[17]
port 90 nsew signal input
rlabel metal2 s 285218 179200 285274 180000 6 data_rdata_i[18]
port 91 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 data_rdata_i[19]
port 92 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 data_rdata_i[1]
port 93 nsew signal input
rlabel metal2 s 411718 179200 411774 180000 6 data_rdata_i[20]
port 94 nsew signal input
rlabel metal2 s 318338 179200 318394 180000 6 data_rdata_i[21]
port 95 nsew signal input
rlabel metal2 s 211618 0 211674 800 6 data_rdata_i[22]
port 96 nsew signal input
rlabel metal2 s 16578 179200 16634 180000 6 data_rdata_i[23]
port 97 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 data_rdata_i[24]
port 98 nsew signal input
rlabel metal3 s 429200 132608 430000 132728 6 data_rdata_i[25]
port 99 nsew signal input
rlabel metal2 s 216678 179200 216734 180000 6 data_rdata_i[26]
port 100 nsew signal input
rlabel metal3 s 429200 27208 430000 27328 6 data_rdata_i[27]
port 101 nsew signal input
rlabel metal2 s 184018 0 184074 800 6 data_rdata_i[28]
port 102 nsew signal input
rlabel metal2 s 326618 179200 326674 180000 6 data_rdata_i[29]
port 103 nsew signal input
rlabel metal2 s 326618 0 326674 800 6 data_rdata_i[2]
port 104 nsew signal input
rlabel metal2 s 164698 0 164754 800 6 data_rdata_i[30]
port 105 nsew signal input
rlabel metal2 s 54758 179200 54814 180000 6 data_rdata_i[31]
port 106 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 data_rdata_i[3]
port 107 nsew signal input
rlabel metal2 s 258078 0 258134 800 6 data_rdata_i[4]
port 108 nsew signal input
rlabel metal2 s 244278 179200 244334 180000 6 data_rdata_i[5]
port 109 nsew signal input
rlabel metal2 s 76838 179200 76894 180000 6 data_rdata_i[6]
port 110 nsew signal input
rlabel metal2 s 304998 0 305054 800 6 data_rdata_i[7]
port 111 nsew signal input
rlabel metal2 s 43718 179200 43774 180000 6 data_rdata_i[8]
port 112 nsew signal input
rlabel metal2 s 120538 179200 120594 180000 6 data_rdata_i[9]
port 113 nsew signal input
rlabel metal2 s 390098 0 390154 800 6 data_req_o
port 114 nsew signal output
rlabel metal2 s 408958 179200 409014 180000 6 data_rvalid_i
port 115 nsew signal input
rlabel metal2 s 252558 0 252614 800 6 data_wdata_o[0]
port 116 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 data_wdata_o[10]
port 117 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 data_wdata_o[11]
port 118 nsew signal output
rlabel metal2 s 213918 179200 213974 180000 6 data_wdata_o[12]
port 119 nsew signal output
rlabel metal3 s 429200 169328 430000 169448 6 data_wdata_o[13]
port 120 nsew signal output
rlabel metal2 s 345938 179200 345994 180000 6 data_wdata_o[14]
port 121 nsew signal output
rlabel metal2 s 156418 179200 156474 180000 6 data_wdata_o[15]
port 122 nsew signal output
rlabel metal2 s 225418 0 225474 800 6 data_wdata_o[16]
port 123 nsew signal output
rlabel metal2 s 222658 0 222714 800 6 data_wdata_o[17]
port 124 nsew signal output
rlabel metal2 s 60278 179200 60334 180000 6 data_wdata_o[18]
port 125 nsew signal output
rlabel metal3 s 429200 23128 430000 23248 6 data_wdata_o[19]
port 126 nsew signal output
rlabel metal2 s 313278 0 313334 800 6 data_wdata_o[1]
port 127 nsew signal output
rlabel metal2 s 365258 0 365314 800 6 data_wdata_o[20]
port 128 nsew signal output
rlabel metal2 s 370778 0 370834 800 6 data_wdata_o[21]
port 129 nsew signal output
rlabel metal2 s 249798 179200 249854 180000 6 data_wdata_o[22]
port 130 nsew signal output
rlabel metal2 s 356518 179200 356574 180000 6 data_wdata_o[23]
port 131 nsew signal output
rlabel metal2 s 206098 0 206154 800 6 data_wdata_o[24]
port 132 nsew signal output
rlabel metal2 s 241518 0 241574 800 6 data_wdata_o[25]
port 133 nsew signal output
rlabel metal2 s 301778 179200 301834 180000 6 data_wdata_o[26]
port 134 nsew signal output
rlabel metal2 s 178498 0 178554 800 6 data_wdata_o[27]
port 135 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 data_wdata_o[28]
port 136 nsew signal output
rlabel metal2 s 90638 179200 90694 180000 6 data_wdata_o[29]
port 137 nsew signal output
rlabel metal3 s 0 170688 800 170808 6 data_wdata_o[2]
port 138 nsew signal output
rlabel metal2 s 79598 179200 79654 180000 6 data_wdata_o[30]
port 139 nsew signal output
rlabel metal3 s 429200 43528 430000 43648 6 data_wdata_o[31]
port 140 nsew signal output
rlabel metal2 s 46478 179200 46534 180000 6 data_wdata_o[3]
port 141 nsew signal output
rlabel metal3 s 429200 63248 430000 63368 6 data_wdata_o[4]
port 142 nsew signal output
rlabel metal2 s 263598 179200 263654 180000 6 data_wdata_o[5]
port 143 nsew signal output
rlabel metal2 s 112718 0 112774 800 6 data_wdata_o[6]
port 144 nsew signal output
rlabel metal3 s 429200 55768 430000 55888 6 data_wdata_o[7]
port 145 nsew signal output
rlabel metal3 s 429200 95888 430000 96008 6 data_wdata_o[8]
port 146 nsew signal output
rlabel metal2 s 370318 179200 370374 180000 6 data_wdata_o[9]
port 147 nsew signal output
rlabel metal3 s 0 133968 800 134088 6 data_we_o
port 148 nsew signal output
rlabel metal2 s 315578 0 315634 800 6 debug_req_i
port 149 nsew signal input
rlabel metal2 s 334898 0 334954 800 6 eFPGA_delay_o[0]
port 150 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 eFPGA_delay_o[1]
port 151 nsew signal output
rlabel metal2 s 189538 179200 189594 180000 6 eFPGA_delay_o[2]
port 152 nsew signal output
rlabel metal2 s 408958 0 409014 800 6 eFPGA_delay_o[3]
port 153 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 eFPGA_en_o
port 154 nsew signal output
rlabel metal2 s 348698 0 348754 800 6 eFPGA_fpga_done_i
port 155 nsew signal input
rlabel metal2 s 211158 179200 211214 180000 6 eFPGA_operand_a_o[0]
port 156 nsew signal output
rlabel metal2 s 30378 179200 30434 180000 6 eFPGA_operand_a_o[10]
port 157 nsew signal output
rlabel metal2 s 269118 179200 269174 180000 6 eFPGA_operand_a_o[11]
port 158 nsew signal output
rlabel metal3 s 429200 67328 430000 67448 6 eFPGA_operand_a_o[12]
port 159 nsew signal output
rlabel metal2 s 417238 179200 417294 180000 6 eFPGA_operand_a_o[13]
port 160 nsew signal output
rlabel metal2 s 378598 179200 378654 180000 6 eFPGA_operand_a_o[14]
port 161 nsew signal output
rlabel metal2 s 238758 179200 238814 180000 6 eFPGA_operand_a_o[15]
port 162 nsew signal output
rlabel metal2 s 288438 0 288494 800 6 eFPGA_operand_a_o[16]
port 163 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 eFPGA_operand_a_o[17]
port 164 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 eFPGA_operand_a_o[18]
port 165 nsew signal output
rlabel metal2 s 321098 179200 321154 180000 6 eFPGA_operand_a_o[19]
port 166 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 eFPGA_operand_a_o[1]
port 167 nsew signal output
rlabel metal2 s 118238 0 118294 800 6 eFPGA_operand_a_o[20]
port 168 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 eFPGA_operand_a_o[21]
port 169 nsew signal output
rlabel metal3 s 0 178848 800 178968 6 eFPGA_operand_a_o[22]
port 170 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 eFPGA_operand_a_o[23]
port 171 nsew signal output
rlabel metal2 s 422758 179200 422814 180000 6 eFPGA_operand_a_o[24]
port 172 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 eFPGA_operand_a_o[25]
port 173 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 eFPGA_operand_a_o[26]
port 174 nsew signal output
rlabel metal2 s 425518 179200 425574 180000 6 eFPGA_operand_a_o[27]
port 175 nsew signal output
rlabel metal2 s 184018 179200 184074 180000 6 eFPGA_operand_a_o[28]
port 176 nsew signal output
rlabel metal2 s 117778 179200 117834 180000 6 eFPGA_operand_a_o[29]
port 177 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 eFPGA_operand_a_o[2]
port 178 nsew signal output
rlabel metal3 s 429200 144848 430000 144968 6 eFPGA_operand_a_o[30]
port 179 nsew signal output
rlabel metal2 s 285678 0 285734 800 6 eFPGA_operand_a_o[31]
port 180 nsew signal output
rlabel metal2 s 340418 0 340474 800 6 eFPGA_operand_a_o[3]
port 181 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 eFPGA_operand_a_o[4]
port 182 nsew signal output
rlabel metal2 s 312818 179200 312874 180000 6 eFPGA_operand_a_o[5]
port 183 nsew signal output
rlabel metal3 s 0 125808 800 125928 6 eFPGA_operand_a_o[6]
port 184 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 eFPGA_operand_a_o[7]
port 185 nsew signal output
rlabel metal2 s 304538 179200 304594 180000 6 eFPGA_operand_a_o[8]
port 186 nsew signal output
rlabel metal2 s 137098 179200 137154 180000 6 eFPGA_operand_a_o[9]
port 187 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 eFPGA_operand_b_o[0]
port 188 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 eFPGA_operand_b_o[10]
port 189 nsew signal output
rlabel metal2 s 411718 0 411774 800 6 eFPGA_operand_b_o[11]
port 190 nsew signal output
rlabel metal2 s 197818 0 197874 800 6 eFPGA_operand_b_o[12]
port 191 nsew signal output
rlabel metal2 s 395158 179200 395214 180000 6 eFPGA_operand_b_o[13]
port 192 nsew signal output
rlabel metal2 s 233698 0 233754 800 6 eFPGA_operand_b_o[14]
port 193 nsew signal output
rlabel metal2 s 161938 179200 161994 180000 6 eFPGA_operand_b_o[15]
port 194 nsew signal output
rlabel metal2 s 343178 179200 343234 180000 6 eFPGA_operand_b_o[16]
port 195 nsew signal output
rlabel metal2 s 428278 179200 428334 180000 6 eFPGA_operand_b_o[17]
port 196 nsew signal output
rlabel metal2 s 478 0 534 800 6 eFPGA_operand_b_o[18]
port 197 nsew signal output
rlabel metal2 s 134338 179200 134394 180000 6 eFPGA_operand_b_o[19]
port 198 nsew signal output
rlabel metal2 s 332138 179200 332194 180000 6 eFPGA_operand_b_o[1]
port 199 nsew signal output
rlabel metal2 s 5538 179200 5594 180000 6 eFPGA_operand_b_o[20]
port 200 nsew signal output
rlabel metal2 s 389638 179200 389694 180000 6 eFPGA_operand_b_o[21]
port 201 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 eFPGA_operand_b_o[22]
port 202 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 eFPGA_operand_b_o[23]
port 203 nsew signal output
rlabel metal2 s 87878 179200 87934 180000 6 eFPGA_operand_b_o[24]
port 204 nsew signal output
rlabel metal2 s 373078 179200 373134 180000 6 eFPGA_operand_b_o[25]
port 205 nsew signal output
rlabel metal2 s 27618 179200 27674 180000 6 eFPGA_operand_b_o[26]
port 206 nsew signal output
rlabel metal2 s 115478 0 115534 800 6 eFPGA_operand_b_o[27]
port 207 nsew signal output
rlabel metal2 s 296258 179200 296314 180000 6 eFPGA_operand_b_o[28]
port 208 nsew signal output
rlabel metal2 s 387338 0 387394 800 6 eFPGA_operand_b_o[29]
port 209 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 eFPGA_operand_b_o[2]
port 210 nsew signal output
rlabel metal2 s 164698 179200 164754 180000 6 eFPGA_operand_b_o[30]
port 211 nsew signal output
rlabel metal2 s 175738 0 175794 800 6 eFPGA_operand_b_o[31]
port 212 nsew signal output
rlabel metal2 s 274638 0 274694 800 6 eFPGA_operand_b_o[3]
port 213 nsew signal output
rlabel metal2 s 159178 179200 159234 180000 6 eFPGA_operand_b_o[4]
port 214 nsew signal output
rlabel metal3 s 429200 148928 430000 149048 6 eFPGA_operand_b_o[5]
port 215 nsew signal output
rlabel metal2 s 192298 0 192354 800 6 eFPGA_operand_b_o[6]
port 216 nsew signal output
rlabel metal2 s 241518 179200 241574 180000 6 eFPGA_operand_b_o[7]
port 217 nsew signal output
rlabel metal2 s 208398 179200 208454 180000 6 eFPGA_operand_b_o[8]
port 218 nsew signal output
rlabel metal2 s 287978 179200 288034 180000 6 eFPGA_operand_b_o[9]
port 219 nsew signal output
rlabel metal2 s 205638 179200 205694 180000 6 eFPGA_operator_o[0]
port 220 nsew signal output
rlabel metal2 s 153658 179200 153714 180000 6 eFPGA_operator_o[1]
port 221 nsew signal output
rlabel metal2 s 321098 0 321154 800 6 eFPGA_result_a_i[0]
port 222 nsew signal input
rlabel metal3 s 429200 79568 430000 79688 6 eFPGA_result_a_i[10]
port 223 nsew signal input
rlabel metal2 s 22098 179200 22154 180000 6 eFPGA_result_a_i[11]
port 224 nsew signal input
rlabel metal3 s 429200 91808 430000 91928 6 eFPGA_result_a_i[12]
port 225 nsew signal input
rlabel metal2 s 68558 179200 68614 180000 6 eFPGA_result_a_i[13]
port 226 nsew signal input
rlabel metal2 s 334898 179200 334954 180000 6 eFPGA_result_a_i[14]
port 227 nsew signal input
rlabel metal2 s 49238 179200 49294 180000 6 eFPGA_result_a_i[15]
port 228 nsew signal input
rlabel metal2 s 417238 0 417294 800 6 eFPGA_result_a_i[16]
port 229 nsew signal input
rlabel metal2 s 38198 179200 38254 180000 6 eFPGA_result_a_i[17]
port 230 nsew signal input
rlabel metal2 s 291198 0 291254 800 6 eFPGA_result_a_i[18]
port 231 nsew signal input
rlabel metal3 s 429200 99968 430000 100088 6 eFPGA_result_a_i[19]
port 232 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 eFPGA_result_a_i[1]
port 233 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 eFPGA_result_a_i[20]
port 234 nsew signal input
rlabel metal2 s 323858 0 323914 800 6 eFPGA_result_a_i[21]
port 235 nsew signal input
rlabel metal2 s 359278 179200 359334 180000 6 eFPGA_result_a_i[22]
port 236 nsew signal input
rlabel metal2 s 112718 179200 112774 180000 6 eFPGA_result_a_i[23]
port 237 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 eFPGA_result_a_i[24]
port 238 nsew signal input
rlabel metal2 s 271878 0 271934 800 6 eFPGA_result_a_i[25]
port 239 nsew signal input
rlabel metal2 s 175738 179200 175794 180000 6 eFPGA_result_a_i[26]
port 240 nsew signal input
rlabel metal2 s 148138 179200 148194 180000 6 eFPGA_result_a_i[27]
port 241 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 eFPGA_result_a_i[28]
port 242 nsew signal input
rlabel metal2 s 353758 179200 353814 180000 6 eFPGA_result_a_i[29]
port 243 nsew signal input
rlabel metal3 s 429200 120368 430000 120488 6 eFPGA_result_a_i[2]
port 244 nsew signal input
rlabel metal2 s 337658 0 337714 800 6 eFPGA_result_a_i[30]
port 245 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 eFPGA_result_a_i[31]
port 246 nsew signal input
rlabel metal2 s 422758 0 422814 800 6 eFPGA_result_a_i[3]
port 247 nsew signal input
rlabel metal2 s 279698 179200 279754 180000 6 eFPGA_result_a_i[4]
port 248 nsew signal input
rlabel metal2 s 13818 179200 13874 180000 6 eFPGA_result_a_i[5]
port 249 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 eFPGA_result_a_i[6]
port 250 nsew signal input
rlabel metal3 s 429200 83648 430000 83768 6 eFPGA_result_a_i[7]
port 251 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 eFPGA_result_a_i[8]
port 252 nsew signal input
rlabel metal2 s 33138 179200 33194 180000 6 eFPGA_result_a_i[9]
port 253 nsew signal input
rlabel metal2 s 101678 179200 101734 180000 6 eFPGA_result_b_i[0]
port 254 nsew signal input
rlabel metal2 s 167458 179200 167514 180000 6 eFPGA_result_b_i[10]
port 255 nsew signal input
rlabel metal2 s 376298 0 376354 800 6 eFPGA_result_b_i[11]
port 256 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 eFPGA_result_b_i[12]
port 257 nsew signal input
rlabel metal2 s 395158 0 395214 800 6 eFPGA_result_b_i[13]
port 258 nsew signal input
rlabel metal2 s 266358 0 266414 800 6 eFPGA_result_b_i[14]
port 259 nsew signal input
rlabel metal2 s 400678 0 400734 800 6 eFPGA_result_b_i[15]
port 260 nsew signal input
rlabel metal2 s 233238 179200 233294 180000 6 eFPGA_result_b_i[16]
port 261 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 eFPGA_result_b_i[17]
port 262 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 eFPGA_result_b_i[18]
port 263 nsew signal input
rlabel metal2 s 274178 179200 274234 180000 6 eFPGA_result_b_i[19]
port 264 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 eFPGA_result_b_i[1]
port 265 nsew signal input
rlabel metal2 s 425518 0 425574 800 6 eFPGA_result_b_i[20]
port 266 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 eFPGA_result_b_i[21]
port 267 nsew signal input
rlabel metal3 s 429200 124448 430000 124568 6 eFPGA_result_b_i[22]
port 268 nsew signal input
rlabel metal3 s 0 121728 800 121848 6 eFPGA_result_b_i[23]
port 269 nsew signal input
rlabel metal2 s 266358 179200 266414 180000 6 eFPGA_result_b_i[24]
port 270 nsew signal input
rlabel metal2 s 24858 179200 24914 180000 6 eFPGA_result_b_i[25]
port 271 nsew signal input
rlabel metal2 s 397918 0 397974 800 6 eFPGA_result_b_i[26]
port 272 nsew signal input
rlabel metal2 s 255318 0 255374 800 6 eFPGA_result_b_i[27]
port 273 nsew signal input
rlabel metal2 s 368018 0 368074 800 6 eFPGA_result_b_i[28]
port 274 nsew signal input
rlabel metal2 s 219438 179200 219494 180000 6 eFPGA_result_b_i[29]
port 275 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 eFPGA_result_b_i[2]
port 276 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 eFPGA_result_b_i[30]
port 277 nsew signal input
rlabel metal2 s 98918 179200 98974 180000 6 eFPGA_result_b_i[31]
port 278 nsew signal input
rlabel metal2 s 362498 0 362554 800 6 eFPGA_result_b_i[3]
port 279 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 eFPGA_result_b_i[4]
port 280 nsew signal input
rlabel metal3 s 429200 136688 430000 136808 6 eFPGA_result_b_i[5]
port 281 nsew signal input
rlabel metal3 s 0 129888 800 130008 6 eFPGA_result_b_i[6]
port 282 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 eFPGA_result_b_i[7]
port 283 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 eFPGA_result_b_i[8]
port 284 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 eFPGA_result_b_i[9]
port 285 nsew signal input
rlabel metal2 s 299478 0 299534 800 6 eFPGA_result_c_i[0]
port 286 nsew signal input
rlabel metal2 s 2778 179200 2834 180000 6 eFPGA_result_c_i[10]
port 287 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 eFPGA_result_c_i[11]
port 288 nsew signal input
rlabel metal2 s 379058 0 379114 800 6 eFPGA_result_c_i[12]
port 289 nsew signal input
rlabel metal2 s 126058 179200 126114 180000 6 eFPGA_result_c_i[13]
port 290 nsew signal input
rlabel metal3 s 429200 128528 430000 128648 6 eFPGA_result_c_i[14]
port 291 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 eFPGA_result_c_i[15]
port 292 nsew signal input
rlabel metal2 s 104438 179200 104494 180000 6 eFPGA_result_c_i[16]
port 293 nsew signal input
rlabel metal2 s 194598 179200 194654 180000 6 eFPGA_result_c_i[17]
port 294 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 eFPGA_result_c_i[18]
port 295 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 eFPGA_result_c_i[19]
port 296 nsew signal input
rlabel metal2 s 128818 179200 128874 180000 6 eFPGA_result_c_i[1]
port 297 nsew signal input
rlabel metal2 s 96158 179200 96214 180000 6 eFPGA_result_c_i[20]
port 298 nsew signal input
rlabel metal3 s 429200 104048 430000 104168 6 eFPGA_result_c_i[21]
port 299 nsew signal input
rlabel metal2 s 172978 0 173034 800 6 eFPGA_result_c_i[22]
port 300 nsew signal input
rlabel metal2 s 384578 0 384634 800 6 eFPGA_result_c_i[23]
port 301 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 eFPGA_result_c_i[24]
port 302 nsew signal input
rlabel metal2 s 260838 179200 260894 180000 6 eFPGA_result_c_i[25]
port 303 nsew signal input
rlabel metal3 s 429200 47608 430000 47728 6 eFPGA_result_c_i[26]
port 304 nsew signal input
rlabel metal2 s 307298 179200 307354 180000 6 eFPGA_result_c_i[27]
port 305 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 eFPGA_result_c_i[28]
port 306 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 eFPGA_result_c_i[29]
port 307 nsew signal input
rlabel metal3 s 429200 112208 430000 112328 6 eFPGA_result_c_i[2]
port 308 nsew signal input
rlabel metal3 s 0 166608 800 166728 6 eFPGA_result_c_i[30]
port 309 nsew signal input
rlabel metal2 s 260838 0 260894 800 6 eFPGA_result_c_i[31]
port 310 nsew signal input
rlabel metal2 s 217138 0 217194 800 6 eFPGA_result_c_i[3]
port 311 nsew signal input
rlabel metal2 s 359738 0 359794 800 6 eFPGA_result_c_i[4]
port 312 nsew signal input
rlabel metal3 s 0 138048 800 138168 6 eFPGA_result_c_i[5]
port 313 nsew signal input
rlabel metal2 s 202878 179200 202934 180000 6 eFPGA_result_c_i[6]
port 314 nsew signal input
rlabel metal2 s 11058 179200 11114 180000 6 eFPGA_result_c_i[7]
port 315 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 eFPGA_result_c_i[8]
port 316 nsew signal input
rlabel metal2 s 142618 179200 142674 180000 6 eFPGA_result_c_i[9]
port 317 nsew signal input
rlabel metal3 s 429200 165248 430000 165368 6 eFPGA_write_strobe_o
port 318 nsew signal output
rlabel metal2 s 373538 0 373594 800 6 ext_perf_counters_i
port 319 nsew signal input
rlabel metal2 s 364798 179200 364854 180000 6 fetch_enable_i
port 320 nsew signal input
rlabel metal2 s 244278 0 244334 800 6 instr_addr_o[0]
port 321 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 instr_addr_o[10]
port 322 nsew signal output
rlabel metal2 s 299018 179200 299074 180000 6 instr_addr_o[11]
port 323 nsew signal output
rlabel metal2 s 238758 0 238814 800 6 instr_addr_o[12]
port 324 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 instr_addr_o[13]
port 325 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 instr_addr_o[14]
port 326 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 instr_addr_o[15]
port 327 nsew signal output
rlabel metal2 s 290738 179200 290794 180000 6 instr_addr_o[16]
port 328 nsew signal output
rlabel metal3 s 429200 108128 430000 108248 6 instr_addr_o[17]
port 329 nsew signal output
rlabel metal3 s 429200 10888 430000 11008 6 instr_addr_o[18]
port 330 nsew signal output
rlabel metal2 s 85118 179200 85174 180000 6 instr_addr_o[19]
port 331 nsew signal output
rlabel metal2 s 200578 0 200634 800 6 instr_addr_o[1]
port 332 nsew signal output
rlabel metal3 s 429200 19048 430000 19168 6 instr_addr_o[20]
port 333 nsew signal output
rlabel metal2 s 343178 0 343234 800 6 instr_addr_o[21]
port 334 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 instr_addr_o[22]
port 335 nsew signal output
rlabel metal2 s 271878 179200 271934 180000 6 instr_addr_o[23]
port 336 nsew signal output
rlabel metal2 s 46938 0 46994 800 6 instr_addr_o[24]
port 337 nsew signal output
rlabel metal2 s 419998 0 420054 800 6 instr_addr_o[25]
port 338 nsew signal output
rlabel metal3 s 429200 71408 430000 71528 6 instr_addr_o[26]
port 339 nsew signal output
rlabel metal2 s 384118 179200 384174 180000 6 instr_addr_o[27]
port 340 nsew signal output
rlabel metal2 s 414478 179200 414534 180000 6 instr_addr_o[28]
port 341 nsew signal output
rlabel metal3 s 429200 157088 430000 157208 6 instr_addr_o[29]
port 342 nsew signal output
rlabel metal2 s 367558 179200 367614 180000 6 instr_addr_o[2]
port 343 nsew signal output
rlabel metal2 s 255318 179200 255374 180000 6 instr_addr_o[30]
port 344 nsew signal output
rlabel metal2 s 22098 0 22154 800 6 instr_addr_o[31]
port 345 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 instr_addr_o[3]
port 346 nsew signal output
rlabel metal2 s 282458 179200 282514 180000 6 instr_addr_o[4]
port 347 nsew signal output
rlabel metal2 s 115018 179200 115074 180000 6 instr_addr_o[5]
port 348 nsew signal output
rlabel metal2 s 107198 179200 107254 180000 6 instr_addr_o[6]
port 349 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 instr_addr_o[7]
port 350 nsew signal output
rlabel metal3 s 429200 14968 430000 15088 6 instr_addr_o[8]
port 351 nsew signal output
rlabel metal2 s 228178 0 228234 800 6 instr_addr_o[9]
port 352 nsew signal output
rlabel metal2 s 302238 0 302294 800 6 instr_gnt_i
port 353 nsew signal input
rlabel metal3 s 0 154368 800 154488 6 instr_rdata_i[0]
port 354 nsew signal input
rlabel metal2 s 35898 179200 35954 180000 6 instr_rdata_i[10]
port 355 nsew signal input
rlabel metal3 s 429200 31288 430000 31408 6 instr_rdata_i[11]
port 356 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 instr_rdata_i[12]
port 357 nsew signal input
rlabel metal2 s 419998 179200 420054 180000 6 instr_rdata_i[13]
port 358 nsew signal input
rlabel metal2 s 362038 179200 362094 180000 6 instr_rdata_i[14]
port 359 nsew signal input
rlabel metal2 s 337658 179200 337714 180000 6 instr_rdata_i[15]
port 360 nsew signal input
rlabel metal2 s 406198 179200 406254 180000 6 instr_rdata_i[16]
port 361 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 instr_rdata_i[17]
port 362 nsew signal input
rlabel metal2 s 392398 179200 392454 180000 6 instr_rdata_i[18]
port 363 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 instr_rdata_i[19]
port 364 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 instr_rdata_i[1]
port 365 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 instr_rdata_i[20]
port 366 nsew signal input
rlabel metal2 s 348698 179200 348754 180000 6 instr_rdata_i[21]
port 367 nsew signal input
rlabel metal2 s 139858 179200 139914 180000 6 instr_rdata_i[22]
port 368 nsew signal input
rlabel metal2 s 82358 179200 82414 180000 6 instr_rdata_i[23]
port 369 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 instr_rdata_i[24]
port 370 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 instr_rdata_i[25]
port 371 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 instr_rdata_i[26]
port 372 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 instr_rdata_i[27]
port 373 nsew signal input
rlabel metal2 s 189538 0 189594 800 6 instr_rdata_i[28]
port 374 nsew signal input
rlabel metal2 s 332138 0 332194 800 6 instr_rdata_i[29]
port 375 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 instr_rdata_i[2]
port 376 nsew signal input
rlabel metal2 s 93398 179200 93454 180000 6 instr_rdata_i[30]
port 377 nsew signal input
rlabel metal2 s 224958 179200 225014 180000 6 instr_rdata_i[31]
port 378 nsew signal input
rlabel metal2 s 397918 179200 397974 180000 6 instr_rdata_i[3]
port 379 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 instr_rdata_i[4]
port 380 nsew signal input
rlabel metal2 s 227718 179200 227774 180000 6 instr_rdata_i[5]
port 381 nsew signal input
rlabel metal2 s 269118 0 269174 800 6 instr_rdata_i[6]
port 382 nsew signal input
rlabel metal2 s 428278 0 428334 800 6 instr_rdata_i[7]
port 383 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 instr_rdata_i[8]
port 384 nsew signal input
rlabel metal2 s 323858 179200 323914 180000 6 instr_rdata_i[9]
port 385 nsew signal input
rlabel metal2 s 57518 179200 57574 180000 6 instr_req_o
port 386 nsew signal output
rlabel metal2 s 172978 179200 173034 180000 6 instr_rvalid_i
port 387 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 irq_ack_o
port 388 nsew signal output
rlabel metal2 s 310058 179200 310114 180000 6 irq_i
port 389 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 irq_id_i[0]
port 390 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 irq_id_i[1]
port 391 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 irq_id_i[2]
port 392 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 irq_id_i[3]
port 393 nsew signal input
rlabel metal2 s 340418 179200 340474 180000 6 irq_id_i[4]
port 394 nsew signal input
rlabel metal3 s 429200 173408 430000 173528 6 irq_id_o[0]
port 395 nsew signal output
rlabel metal2 s 235998 0 236054 800 6 irq_id_o[1]
port 396 nsew signal output
rlabel metal2 s 296718 0 296774 800 6 irq_id_o[2]
port 397 nsew signal output
rlabel metal2 s 200118 179200 200174 180000 6 irq_id_o[3]
port 398 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 irq_id_o[4]
port 399 nsew signal output
rlabel metal2 s 277398 0 277454 800 6 rst_ni
port 400 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 test_en_i
port 401 nsew signal input
rlabel metal4 s 403568 2128 403888 177392 6 VPWR
port 402 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 177392 6 VPWR
port 403 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 177392 6 VPWR
port 404 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 177392 6 VPWR
port 405 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 177392 6 VPWR
port 406 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 177392 6 VPWR
port 407 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 177392 6 VPWR
port 408 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 177392 6 VPWR
port 409 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 177392 6 VPWR
port 410 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 177392 6 VPWR
port 411 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 177392 6 VPWR
port 412 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 177392 6 VPWR
port 413 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 177392 6 VPWR
port 414 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 177392 6 VPWR
port 415 nsew power bidirectional
rlabel metal5 s 1104 158478 428812 158798 6 VPWR
port 416 nsew power bidirectional
rlabel metal5 s 1104 127842 428812 128162 6 VPWR
port 417 nsew power bidirectional
rlabel metal5 s 1104 97206 428812 97526 6 VPWR
port 418 nsew power bidirectional
rlabel metal5 s 1104 66570 428812 66890 6 VPWR
port 419 nsew power bidirectional
rlabel metal5 s 1104 35934 428812 36254 6 VPWR
port 420 nsew power bidirectional
rlabel metal5 s 1104 5298 428812 5618 6 VPWR
port 421 nsew power bidirectional
rlabel metal4 s 418928 2128 419248 177392 6 VGND
port 422 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 177392 6 VGND
port 423 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 177392 6 VGND
port 424 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 177392 6 VGND
port 425 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 177392 6 VGND
port 426 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 177392 6 VGND
port 427 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 177392 6 VGND
port 428 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 177392 6 VGND
port 429 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 177392 6 VGND
port 430 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 177392 6 VGND
port 431 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 177392 6 VGND
port 432 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 177392 6 VGND
port 433 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 177392 6 VGND
port 434 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 177392 6 VGND
port 435 nsew ground bidirectional
rlabel metal5 s 1104 173796 428812 174116 6 VGND
port 436 nsew ground bidirectional
rlabel metal5 s 1104 143160 428812 143480 6 VGND
port 437 nsew ground bidirectional
rlabel metal5 s 1104 112524 428812 112844 6 VGND
port 438 nsew ground bidirectional
rlabel metal5 s 1104 81888 428812 82208 6 VGND
port 439 nsew ground bidirectional
rlabel metal5 s 1104 51252 428812 51572 6 VGND
port 440 nsew ground bidirectional
rlabel metal5 s 1104 20616 428812 20936 6 VGND
port 441 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 430000 180000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 71523502
string GDS_START 1211584
<< end >>

