VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core_sram
  CLASS BLOCK ;
  FOREIGN core_sram ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 800.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.590 0.000 1161.870 4.000 ;
    END
  END clk_i
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 737.840 1200.000 738.440 ;
    END
  END debug_req_i
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.190 796.000 1028.470 800.000 ;
    END
  END eFPGA_delay_o[0]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.490 0.000 1122.770 4.000 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 796.000 740.970 800.000 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 796.000 349.970 800.000 ;
    END
  END eFPGA_en_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 700.440 1200.000 701.040 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 0.000 1097.470 4.000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.590 796.000 1000.870 800.000 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 374.040 1200.000 374.640 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 796.000 883.570 800.000 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 796.000 11.870 800.000 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 796.000 232.670 800.000 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 622.240 1200.000 622.840 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 44.240 1200.000 44.840 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 102.040 1200.000 102.640 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1170.790 796.000 1171.070 800.000 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 796.000 1196.370 800.000 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 796.000 715.670 800.000 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 180.240 1200.000 180.840 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 0.000 941.070 4.000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 796.000 609.870 800.000 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 796.000 975.570 800.000 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 796.000 375.270 800.000 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 796.000 453.470 800.000 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 796.000 1145.770 800.000 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 796.000 1118.170 800.000 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 796.000 545.470 800.000 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.090 0.000 575.370 4.000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 796.000 637.470 800.000 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 796.000 336.170 800.000 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 0.000 1044.570 4.000 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 796.000 129.170 800.000 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 431.840 1200.000 432.440 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 796.000 676.570 800.000 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 796.000 467.270 800.000 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.890 796.000 911.170 800.000 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 796.000 76.270 800.000 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 0.000 784.670 4.000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 564.440 1200.000 565.040 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 200.640 1200.000 201.240 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 796.000 662.770 800.000 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 796.000 805.370 800.000 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.890 0.000 888.170 4.000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 547.440 1200.000 548.040 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 796.000 207.370 800.000 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 796.000 648.970 800.000 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 796.000 1131.970 800.000 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 796.000 179.770 800.000 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 796.000 793.870 800.000 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 796.000 363.770 800.000 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 796.000 193.570 800.000 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 605.240 1200.000 605.840 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 0.000 67.070 4.000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 0.000 1175.670 4.000 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 796.000 492.570 800.000 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 758.240 1200.000 758.840 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 796.000 481.070 800.000 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.890 796.000 819.170 800.000 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 796.000 414.370 800.000 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.990 796.000 858.270 800.000 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 796.000 950.270 800.000 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 796.000 428.170 800.000 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 411.440 1200.000 412.040 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.790 796.000 872.070 800.000 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 353.640 1200.000 354.240 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 796.000 402.870 800.000 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 796.000 598.370 800.000 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.390 796.000 1106.670 800.000 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 796.000 780.070 800.000 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 0.000 849.070 4.000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 796.000 584.570 800.000 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 796.000 520.170 800.000 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 778.640 1200.000 779.240 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.590 796.000 1184.870 800.000 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 796.000 154.470 800.000 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 771.840 4.000 772.440 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.490 796.000 961.770 800.000 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 796.000 1157.270 800.000 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.790 0.000 1148.070 4.000 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.490 0.000 823.770 4.000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 796.000 389.070 800.000 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 796.000 559.270 800.000 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 796.000 766.270 800.000 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 979.890 0.000 980.170 4.000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 796.000 623.670 800.000 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 85.040 1200.000 85.640 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.690 0.000 901.970 4.000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 6.840 1200.000 7.440 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 142.840 1200.000 143.440 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 796.000 271.770 800.000 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 796.000 90.070 800.000 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 0.000 835.270 4.000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 796.000 936.470 800.000 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 796.000 50.970 800.000 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 333.240 1200.000 333.840 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 796.000 570.770 800.000 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.690 796.000 1039.970 800.000 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 275.440 1200.000 276.040 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 796.000 297.070 800.000 ;
    END
  END eFPGA_write_strobe_o
  PIN ext_data_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.390 0.000 1083.670 4.000 ;
    END
  END ext_data_addr_i[0]
  PIN ext_data_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 796.000 1067.570 800.000 ;
    END
  END ext_data_addr_i[1]
  PIN ext_data_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END ext_data_addr_i[2]
  PIN ext_data_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END ext_data_addr_i[3]
  PIN ext_data_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END ext_data_addr_i[4]
  PIN ext_data_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 0.000 1058.370 4.000 ;
    END
  END ext_data_addr_i[5]
  PIN ext_data_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END ext_data_addr_i[6]
  PIN ext_data_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 0.000 770.870 4.000 ;
    END
  END ext_data_addr_i[7]
  PIN ext_data_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 796.000 310.870 800.000 ;
    END
  END ext_data_addr_i[8]
  PIN ext_data_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 952.290 0.000 952.570 4.000 ;
    END
  END ext_data_addr_i[9]
  PIN ext_data_be_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END ext_data_be_i[0]
  PIN ext_data_be_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 448.840 1200.000 449.440 ;
    END
  END ext_data_be_i[1]
  PIN ext_data_be_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 796.000 23.370 800.000 ;
    END
  END ext_data_be_i[2]
  PIN ext_data_be_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 663.040 1200.000 663.640 ;
    END
  END ext_data_be_i[3]
  PIN ext_data_rdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 796.000 257.970 800.000 ;
    END
  END ext_data_rdata_o[0]
  PIN ext_data_rdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 159.840 1200.000 160.440 ;
    END
  END ext_data_rdata_o[10]
  PIN ext_data_rdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END ext_data_rdata_o[11]
  PIN ext_data_rdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END ext_data_rdata_o[12]
  PIN ext_data_rdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.790 796.000 1079.070 800.000 ;
    END
  END ext_data_rdata_o[13]
  PIN ext_data_rdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 796.000 168.270 800.000 ;
    END
  END ext_data_rdata_o[14]
  PIN ext_data_rdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 796.000 727.170 800.000 ;
    END
  END ext_data_rdata_o[15]
  PIN ext_data_rdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 796.000 832.970 800.000 ;
    END
  END ext_data_rdata_o[16]
  PIN ext_data_rdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.990 0.000 927.270 4.000 ;
    END
  END ext_data_rdata_o[17]
  PIN ext_data_rdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 796.000 324.670 800.000 ;
    END
  END ext_data_rdata_o[18]
  PIN ext_data_rdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 796.000 441.970 800.000 ;
    END
  END ext_data_rdata_o[19]
  PIN ext_data_rdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 796.000 218.870 800.000 ;
    END
  END ext_data_rdata_o[1]
  PIN ext_data_rdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.090 796.000 989.370 800.000 ;
    END
  END ext_data_rdata_o[20]
  PIN ext_data_rdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 27.240 1200.000 27.840 ;
    END
  END ext_data_rdata_o[21]
  PIN ext_data_rdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 796.000 140.670 800.000 ;
    END
  END ext_data_rdata_o[22]
  PIN ext_data_rdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.290 796.000 285.570 800.000 ;
    END
  END ext_data_rdata_o[23]
  PIN ext_data_rdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END ext_data_rdata_o[24]
  PIN ext_data_rdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END ext_data_rdata_o[25]
  PIN ext_data_rdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 796.000 62.470 800.000 ;
    END
  END ext_data_rdata_o[26]
  PIN ext_data_rdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END ext_data_rdata_o[27]
  PIN ext_data_rdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END ext_data_rdata_o[28]
  PIN ext_data_rdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END ext_data_rdata_o[29]
  PIN ext_data_rdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END ext_data_rdata_o[2]
  PIN ext_data_rdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 0.000 1030.770 4.000 ;
    END
  END ext_data_rdata_o[30]
  PIN ext_data_rdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END ext_data_rdata_o[31]
  PIN ext_data_rdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 584.840 1200.000 585.440 ;
    END
  END ext_data_rdata_o[3]
  PIN ext_data_rdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 796.000 506.370 800.000 ;
    END
  END ext_data_rdata_o[4]
  PIN ext_data_rdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 642.640 1200.000 643.240 ;
    END
  END ext_data_rdata_o[5]
  PIN ext_data_rdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 122.440 1200.000 123.040 ;
    END
  END ext_data_rdata_o[6]
  PIN ext_data_rdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END ext_data_rdata_o[7]
  PIN ext_data_rdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 720.840 1200.000 721.440 ;
    END
  END ext_data_rdata_o[8]
  PIN ext_data_rdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END ext_data_rdata_o[9]
  PIN ext_data_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 295.840 1200.000 296.440 ;
    END
  END ext_data_req_i
  PIN ext_data_rvalid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 506.640 1200.000 507.240 ;
    END
  END ext_data_rvalid_o
  PIN ext_data_wdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END ext_data_wdata_i[0]
  PIN ext_data_wdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.290 0.000 1136.570 4.000 ;
    END
  END ext_data_wdata_i[10]
  PIN ext_data_wdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END ext_data_wdata_i[11]
  PIN ext_data_wdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 217.640 1200.000 218.240 ;
    END
  END ext_data_wdata_i[12]
  PIN ext_data_wdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END ext_data_wdata_i[13]
  PIN ext_data_wdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.190 796.000 844.470 800.000 ;
    END
  END ext_data_wdata_i[14]
  PIN ext_data_wdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END ext_data_wdata_i[15]
  PIN ext_data_wdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 796.000 115.370 800.000 ;
    END
  END ext_data_wdata_i[16]
  PIN ext_data_wdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.090 0.000 874.370 4.000 ;
    END
  END ext_data_wdata_i[17]
  PIN ext_data_wdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.490 796.000 1053.770 800.000 ;
    END
  END ext_data_wdata_i[18]
  PIN ext_data_wdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END ext_data_wdata_i[19]
  PIN ext_data_wdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 0.000 1108.970 4.000 ;
    END
  END ext_data_wdata_i[1]
  PIN ext_data_wdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 796.000 37.170 800.000 ;
    END
  END ext_data_wdata_i[20]
  PIN ext_data_wdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 64.640 1200.000 65.240 ;
    END
  END ext_data_wdata_i[21]
  PIN ext_data_wdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 527.040 1200.000 527.640 ;
    END
  END ext_data_wdata_i[22]
  PIN ext_data_wdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END ext_data_wdata_i[23]
  PIN ext_data_wdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 238.040 1200.000 238.640 ;
    END
  END ext_data_wdata_i[24]
  PIN ext_data_wdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END ext_data_wdata_i[25]
  PIN ext_data_wdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 796.000 754.770 800.000 ;
    END
  END ext_data_wdata_i[26]
  PIN ext_data_wdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 796.000 701.870 800.000 ;
    END
  END ext_data_wdata_i[27]
  PIN ext_data_wdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END ext_data_wdata_i[28]
  PIN ext_data_wdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 796.000 246.470 800.000 ;
    END
  END ext_data_wdata_i[29]
  PIN ext_data_wdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 796.000 101.570 800.000 ;
    END
  END ext_data_wdata_i[2]
  PIN ext_data_wdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 796.000 1092.870 800.000 ;
    END
  END ext_data_wdata_i[30]
  PIN ext_data_wdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END ext_data_wdata_i[31]
  PIN ext_data_wdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 391.040 1200.000 391.640 ;
    END
  END ext_data_wdata_i[3]
  PIN ext_data_wdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 258.440 1200.000 259.040 ;
    END
  END ext_data_wdata_i[4]
  PIN ext_data_wdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END ext_data_wdata_i[5]
  PIN ext_data_wdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 4.000 ;
    END
  END ext_data_wdata_i[6]
  PIN ext_data_wdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END ext_data_wdata_i[7]
  PIN ext_data_wdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 4.000 ;
    END
  END ext_data_wdata_i[8]
  PIN ext_data_wdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 489.640 1200.000 490.240 ;
    END
  END ext_data_wdata_i[9]
  PIN ext_data_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 796.000 897.370 800.000 ;
    END
  END ext_data_we_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END fetch_enable_i
  PIN irq_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END irq_ack_o
  PIN irq_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 680.040 1200.000 680.640 ;
    END
  END irq_i
  PIN irq_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END irq_id_i[0]
  PIN irq_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END irq_id_i[1]
  PIN irq_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 796.000 1014.670 800.000 ;
    END
  END irq_id_i[2]
  PIN irq_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 796.000 688.070 800.000 ;
    END
  END irq_id_i[3]
  PIN irq_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 796.000 531.670 800.000 ;
    END
  END irq_id_i[4]
  PIN irq_id_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 0.000 1019.270 4.000 ;
    END
  END irq_id_o[0]
  PIN irq_id_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 469.240 1200.000 469.840 ;
    END
  END irq_id_o[1]
  PIN irq_id_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END irq_id_o[2]
  PIN irq_id_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1196.000 316.240 1200.000 316.840 ;
    END
  END irq_id_o[3]
  PIN irq_id_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 796.000 922.670 800.000 ;
    END
  END irq_id_o[4]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END reset
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 477.260 522.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 477.260 472.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 477.260 422.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 477.260 372.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 477.260 322.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 477.260 272.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 477.260 222.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 477.260 172.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 477.260 122.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 477.260 72.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 70.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 1194.160 640.810 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 1194.160 487.630 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 1194.160 334.450 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 1194.160 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 1194.160 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 477.260 547.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 477.260 497.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 477.260 447.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 477.260 397.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 477.260 347.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 477.260 297.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 477.260 247.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 477.260 197.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 477.260 147.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 477.260 97.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 789.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 70.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 715.800 1194.160 717.400 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 1194.160 564.220 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 1194.160 411.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 1194.160 257.860 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 1194.160 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.935 794.155 ;
      LAYER met1 ;
        RECT 2.370 9.220 1196.390 794.200 ;
      LAYER met2 ;
        RECT 2.400 795.720 11.310 796.000 ;
        RECT 12.150 795.720 22.810 796.000 ;
        RECT 23.650 795.720 36.610 796.000 ;
        RECT 37.450 795.720 50.410 796.000 ;
        RECT 51.250 795.720 61.910 796.000 ;
        RECT 62.750 795.720 75.710 796.000 ;
        RECT 76.550 795.720 89.510 796.000 ;
        RECT 90.350 795.720 101.010 796.000 ;
        RECT 101.850 795.720 114.810 796.000 ;
        RECT 115.650 795.720 128.610 796.000 ;
        RECT 129.450 795.720 140.110 796.000 ;
        RECT 140.950 795.720 153.910 796.000 ;
        RECT 154.750 795.720 167.710 796.000 ;
        RECT 168.550 795.720 179.210 796.000 ;
        RECT 180.050 795.720 193.010 796.000 ;
        RECT 193.850 795.720 206.810 796.000 ;
        RECT 207.650 795.720 218.310 796.000 ;
        RECT 219.150 795.720 232.110 796.000 ;
        RECT 232.950 795.720 245.910 796.000 ;
        RECT 246.750 795.720 257.410 796.000 ;
        RECT 258.250 795.720 271.210 796.000 ;
        RECT 272.050 795.720 285.010 796.000 ;
        RECT 285.850 795.720 296.510 796.000 ;
        RECT 297.350 795.720 310.310 796.000 ;
        RECT 311.150 795.720 324.110 796.000 ;
        RECT 324.950 795.720 335.610 796.000 ;
        RECT 336.450 795.720 349.410 796.000 ;
        RECT 350.250 795.720 363.210 796.000 ;
        RECT 364.050 795.720 374.710 796.000 ;
        RECT 375.550 795.720 388.510 796.000 ;
        RECT 389.350 795.720 402.310 796.000 ;
        RECT 403.150 795.720 413.810 796.000 ;
        RECT 414.650 795.720 427.610 796.000 ;
        RECT 428.450 795.720 441.410 796.000 ;
        RECT 442.250 795.720 452.910 796.000 ;
        RECT 453.750 795.720 466.710 796.000 ;
        RECT 467.550 795.720 480.510 796.000 ;
        RECT 481.350 795.720 492.010 796.000 ;
        RECT 492.850 795.720 505.810 796.000 ;
        RECT 506.650 795.720 519.610 796.000 ;
        RECT 520.450 795.720 531.110 796.000 ;
        RECT 531.950 795.720 544.910 796.000 ;
        RECT 545.750 795.720 558.710 796.000 ;
        RECT 559.550 795.720 570.210 796.000 ;
        RECT 571.050 795.720 584.010 796.000 ;
        RECT 584.850 795.720 597.810 796.000 ;
        RECT 598.650 795.720 609.310 796.000 ;
        RECT 610.150 795.720 623.110 796.000 ;
        RECT 623.950 795.720 636.910 796.000 ;
        RECT 637.750 795.720 648.410 796.000 ;
        RECT 649.250 795.720 662.210 796.000 ;
        RECT 663.050 795.720 676.010 796.000 ;
        RECT 676.850 795.720 687.510 796.000 ;
        RECT 688.350 795.720 701.310 796.000 ;
        RECT 702.150 795.720 715.110 796.000 ;
        RECT 715.950 795.720 726.610 796.000 ;
        RECT 727.450 795.720 740.410 796.000 ;
        RECT 741.250 795.720 754.210 796.000 ;
        RECT 755.050 795.720 765.710 796.000 ;
        RECT 766.550 795.720 779.510 796.000 ;
        RECT 780.350 795.720 793.310 796.000 ;
        RECT 794.150 795.720 804.810 796.000 ;
        RECT 805.650 795.720 818.610 796.000 ;
        RECT 819.450 795.720 832.410 796.000 ;
        RECT 833.250 795.720 843.910 796.000 ;
        RECT 844.750 795.720 857.710 796.000 ;
        RECT 858.550 795.720 871.510 796.000 ;
        RECT 872.350 795.720 883.010 796.000 ;
        RECT 883.850 795.720 896.810 796.000 ;
        RECT 897.650 795.720 910.610 796.000 ;
        RECT 911.450 795.720 922.110 796.000 ;
        RECT 922.950 795.720 935.910 796.000 ;
        RECT 936.750 795.720 949.710 796.000 ;
        RECT 950.550 795.720 961.210 796.000 ;
        RECT 962.050 795.720 975.010 796.000 ;
        RECT 975.850 795.720 988.810 796.000 ;
        RECT 989.650 795.720 1000.310 796.000 ;
        RECT 1001.150 795.720 1014.110 796.000 ;
        RECT 1014.950 795.720 1027.910 796.000 ;
        RECT 1028.750 795.720 1039.410 796.000 ;
        RECT 1040.250 795.720 1053.210 796.000 ;
        RECT 1054.050 795.720 1067.010 796.000 ;
        RECT 1067.850 795.720 1078.510 796.000 ;
        RECT 1079.350 795.720 1092.310 796.000 ;
        RECT 1093.150 795.720 1106.110 796.000 ;
        RECT 1106.950 795.720 1117.610 796.000 ;
        RECT 1118.450 795.720 1131.410 796.000 ;
        RECT 1132.250 795.720 1145.210 796.000 ;
        RECT 1146.050 795.720 1156.710 796.000 ;
        RECT 1157.550 795.720 1170.510 796.000 ;
        RECT 1171.350 795.720 1184.310 796.000 ;
        RECT 1185.150 795.720 1195.810 796.000 ;
        RECT 2.400 4.280 1196.360 795.720 ;
        RECT 2.950 4.000 13.610 4.280 ;
        RECT 14.450 4.000 27.410 4.280 ;
        RECT 28.250 4.000 41.210 4.280 ;
        RECT 42.050 4.000 52.710 4.280 ;
        RECT 53.550 4.000 66.510 4.280 ;
        RECT 67.350 4.000 80.310 4.280 ;
        RECT 81.150 4.000 91.810 4.280 ;
        RECT 92.650 4.000 105.610 4.280 ;
        RECT 106.450 4.000 119.410 4.280 ;
        RECT 120.250 4.000 130.910 4.280 ;
        RECT 131.750 4.000 144.710 4.280 ;
        RECT 145.550 4.000 158.510 4.280 ;
        RECT 159.350 4.000 170.010 4.280 ;
        RECT 170.850 4.000 183.810 4.280 ;
        RECT 184.650 4.000 197.610 4.280 ;
        RECT 198.450 4.000 209.110 4.280 ;
        RECT 209.950 4.000 222.910 4.280 ;
        RECT 223.750 4.000 236.710 4.280 ;
        RECT 237.550 4.000 248.210 4.280 ;
        RECT 249.050 4.000 262.010 4.280 ;
        RECT 262.850 4.000 275.810 4.280 ;
        RECT 276.650 4.000 287.310 4.280 ;
        RECT 288.150 4.000 301.110 4.280 ;
        RECT 301.950 4.000 314.910 4.280 ;
        RECT 315.750 4.000 326.410 4.280 ;
        RECT 327.250 4.000 340.210 4.280 ;
        RECT 341.050 4.000 354.010 4.280 ;
        RECT 354.850 4.000 365.510 4.280 ;
        RECT 366.350 4.000 379.310 4.280 ;
        RECT 380.150 4.000 393.110 4.280 ;
        RECT 393.950 4.000 404.610 4.280 ;
        RECT 405.450 4.000 418.410 4.280 ;
        RECT 419.250 4.000 432.210 4.280 ;
        RECT 433.050 4.000 443.710 4.280 ;
        RECT 444.550 4.000 457.510 4.280 ;
        RECT 458.350 4.000 471.310 4.280 ;
        RECT 472.150 4.000 482.810 4.280 ;
        RECT 483.650 4.000 496.610 4.280 ;
        RECT 497.450 4.000 510.410 4.280 ;
        RECT 511.250 4.000 521.910 4.280 ;
        RECT 522.750 4.000 535.710 4.280 ;
        RECT 536.550 4.000 549.510 4.280 ;
        RECT 550.350 4.000 561.010 4.280 ;
        RECT 561.850 4.000 574.810 4.280 ;
        RECT 575.650 4.000 588.610 4.280 ;
        RECT 589.450 4.000 600.110 4.280 ;
        RECT 600.950 4.000 613.910 4.280 ;
        RECT 614.750 4.000 627.710 4.280 ;
        RECT 628.550 4.000 639.210 4.280 ;
        RECT 640.050 4.000 653.010 4.280 ;
        RECT 653.850 4.000 666.810 4.280 ;
        RECT 667.650 4.000 678.310 4.280 ;
        RECT 679.150 4.000 692.110 4.280 ;
        RECT 692.950 4.000 705.910 4.280 ;
        RECT 706.750 4.000 717.410 4.280 ;
        RECT 718.250 4.000 731.210 4.280 ;
        RECT 732.050 4.000 745.010 4.280 ;
        RECT 745.850 4.000 756.510 4.280 ;
        RECT 757.350 4.000 770.310 4.280 ;
        RECT 771.150 4.000 784.110 4.280 ;
        RECT 784.950 4.000 795.610 4.280 ;
        RECT 796.450 4.000 809.410 4.280 ;
        RECT 810.250 4.000 823.210 4.280 ;
        RECT 824.050 4.000 834.710 4.280 ;
        RECT 835.550 4.000 848.510 4.280 ;
        RECT 849.350 4.000 862.310 4.280 ;
        RECT 863.150 4.000 873.810 4.280 ;
        RECT 874.650 4.000 887.610 4.280 ;
        RECT 888.450 4.000 901.410 4.280 ;
        RECT 902.250 4.000 912.910 4.280 ;
        RECT 913.750 4.000 926.710 4.280 ;
        RECT 927.550 4.000 940.510 4.280 ;
        RECT 941.350 4.000 952.010 4.280 ;
        RECT 952.850 4.000 965.810 4.280 ;
        RECT 966.650 4.000 979.610 4.280 ;
        RECT 980.450 4.000 991.110 4.280 ;
        RECT 991.950 4.000 1004.910 4.280 ;
        RECT 1005.750 4.000 1018.710 4.280 ;
        RECT 1019.550 4.000 1030.210 4.280 ;
        RECT 1031.050 4.000 1044.010 4.280 ;
        RECT 1044.850 4.000 1057.810 4.280 ;
        RECT 1058.650 4.000 1069.310 4.280 ;
        RECT 1070.150 4.000 1083.110 4.280 ;
        RECT 1083.950 4.000 1096.910 4.280 ;
        RECT 1097.750 4.000 1108.410 4.280 ;
        RECT 1109.250 4.000 1122.210 4.280 ;
        RECT 1123.050 4.000 1136.010 4.280 ;
        RECT 1136.850 4.000 1147.510 4.280 ;
        RECT 1148.350 4.000 1161.310 4.280 ;
        RECT 1162.150 4.000 1175.110 4.280 ;
        RECT 1175.950 4.000 1186.610 4.280 ;
        RECT 1187.450 4.000 1196.360 4.280 ;
      LAYER met3 ;
        RECT 4.400 791.840 1196.000 792.705 ;
        RECT 4.000 779.640 1196.000 791.840 ;
        RECT 4.000 778.240 1195.600 779.640 ;
        RECT 4.000 772.840 1196.000 778.240 ;
        RECT 4.400 771.440 1196.000 772.840 ;
        RECT 4.000 759.240 1196.000 771.440 ;
        RECT 4.000 757.840 1195.600 759.240 ;
        RECT 4.000 755.840 1196.000 757.840 ;
        RECT 4.400 754.440 1196.000 755.840 ;
        RECT 4.000 738.840 1196.000 754.440 ;
        RECT 4.000 737.440 1195.600 738.840 ;
        RECT 4.000 735.440 1196.000 737.440 ;
        RECT 4.400 734.040 1196.000 735.440 ;
        RECT 4.000 721.840 1196.000 734.040 ;
        RECT 4.000 720.440 1195.600 721.840 ;
        RECT 4.000 715.040 1196.000 720.440 ;
        RECT 4.400 713.640 1196.000 715.040 ;
        RECT 4.000 701.440 1196.000 713.640 ;
        RECT 4.000 700.040 1195.600 701.440 ;
        RECT 4.000 698.040 1196.000 700.040 ;
        RECT 4.400 696.640 1196.000 698.040 ;
        RECT 4.000 681.040 1196.000 696.640 ;
        RECT 4.000 679.640 1195.600 681.040 ;
        RECT 4.000 677.640 1196.000 679.640 ;
        RECT 4.400 676.240 1196.000 677.640 ;
        RECT 4.000 664.040 1196.000 676.240 ;
        RECT 4.000 662.640 1195.600 664.040 ;
        RECT 4.000 657.240 1196.000 662.640 ;
        RECT 4.400 655.840 1196.000 657.240 ;
        RECT 4.000 643.640 1196.000 655.840 ;
        RECT 4.000 642.240 1195.600 643.640 ;
        RECT 4.000 640.240 1196.000 642.240 ;
        RECT 4.400 638.840 1196.000 640.240 ;
        RECT 4.000 623.240 1196.000 638.840 ;
        RECT 4.000 621.840 1195.600 623.240 ;
        RECT 4.000 619.840 1196.000 621.840 ;
        RECT 4.400 618.440 1196.000 619.840 ;
        RECT 4.000 606.240 1196.000 618.440 ;
        RECT 4.000 604.840 1195.600 606.240 ;
        RECT 4.000 599.440 1196.000 604.840 ;
        RECT 4.400 598.040 1196.000 599.440 ;
        RECT 4.000 585.840 1196.000 598.040 ;
        RECT 4.000 584.440 1195.600 585.840 ;
        RECT 4.000 582.440 1196.000 584.440 ;
        RECT 4.400 581.040 1196.000 582.440 ;
        RECT 4.000 565.440 1196.000 581.040 ;
        RECT 4.000 564.040 1195.600 565.440 ;
        RECT 4.000 562.040 1196.000 564.040 ;
        RECT 4.400 560.640 1196.000 562.040 ;
        RECT 4.000 548.440 1196.000 560.640 ;
        RECT 4.000 547.040 1195.600 548.440 ;
        RECT 4.000 541.640 1196.000 547.040 ;
        RECT 4.400 540.240 1196.000 541.640 ;
        RECT 4.000 528.040 1196.000 540.240 ;
        RECT 4.000 526.640 1195.600 528.040 ;
        RECT 4.000 524.640 1196.000 526.640 ;
        RECT 4.400 523.240 1196.000 524.640 ;
        RECT 4.000 507.640 1196.000 523.240 ;
        RECT 4.000 506.240 1195.600 507.640 ;
        RECT 4.000 504.240 1196.000 506.240 ;
        RECT 4.400 502.840 1196.000 504.240 ;
        RECT 4.000 490.640 1196.000 502.840 ;
        RECT 4.000 489.240 1195.600 490.640 ;
        RECT 4.000 483.840 1196.000 489.240 ;
        RECT 4.400 482.440 1196.000 483.840 ;
        RECT 4.000 470.240 1196.000 482.440 ;
        RECT 4.000 468.840 1195.600 470.240 ;
        RECT 4.000 466.840 1196.000 468.840 ;
        RECT 4.400 465.440 1196.000 466.840 ;
        RECT 4.000 449.840 1196.000 465.440 ;
        RECT 4.000 448.440 1195.600 449.840 ;
        RECT 4.000 446.440 1196.000 448.440 ;
        RECT 4.400 445.040 1196.000 446.440 ;
        RECT 4.000 432.840 1196.000 445.040 ;
        RECT 4.000 431.440 1195.600 432.840 ;
        RECT 4.000 426.040 1196.000 431.440 ;
        RECT 4.400 424.640 1196.000 426.040 ;
        RECT 4.000 412.440 1196.000 424.640 ;
        RECT 4.000 411.040 1195.600 412.440 ;
        RECT 4.000 409.040 1196.000 411.040 ;
        RECT 4.400 407.640 1196.000 409.040 ;
        RECT 4.000 392.040 1196.000 407.640 ;
        RECT 4.000 390.640 1195.600 392.040 ;
        RECT 4.000 388.640 1196.000 390.640 ;
        RECT 4.400 387.240 1196.000 388.640 ;
        RECT 4.000 375.040 1196.000 387.240 ;
        RECT 4.000 373.640 1195.600 375.040 ;
        RECT 4.000 368.240 1196.000 373.640 ;
        RECT 4.400 366.840 1196.000 368.240 ;
        RECT 4.000 354.640 1196.000 366.840 ;
        RECT 4.000 353.240 1195.600 354.640 ;
        RECT 4.000 351.240 1196.000 353.240 ;
        RECT 4.400 349.840 1196.000 351.240 ;
        RECT 4.000 334.240 1196.000 349.840 ;
        RECT 4.000 332.840 1195.600 334.240 ;
        RECT 4.000 330.840 1196.000 332.840 ;
        RECT 4.400 329.440 1196.000 330.840 ;
        RECT 4.000 317.240 1196.000 329.440 ;
        RECT 4.000 315.840 1195.600 317.240 ;
        RECT 4.000 310.440 1196.000 315.840 ;
        RECT 4.400 309.040 1196.000 310.440 ;
        RECT 4.000 296.840 1196.000 309.040 ;
        RECT 4.000 295.440 1195.600 296.840 ;
        RECT 4.000 293.440 1196.000 295.440 ;
        RECT 4.400 292.040 1196.000 293.440 ;
        RECT 4.000 276.440 1196.000 292.040 ;
        RECT 4.000 275.040 1195.600 276.440 ;
        RECT 4.000 273.040 1196.000 275.040 ;
        RECT 4.400 271.640 1196.000 273.040 ;
        RECT 4.000 259.440 1196.000 271.640 ;
        RECT 4.000 258.040 1195.600 259.440 ;
        RECT 4.000 252.640 1196.000 258.040 ;
        RECT 4.400 251.240 1196.000 252.640 ;
        RECT 4.000 239.040 1196.000 251.240 ;
        RECT 4.000 237.640 1195.600 239.040 ;
        RECT 4.000 235.640 1196.000 237.640 ;
        RECT 4.400 234.240 1196.000 235.640 ;
        RECT 4.000 218.640 1196.000 234.240 ;
        RECT 4.000 217.240 1195.600 218.640 ;
        RECT 4.000 215.240 1196.000 217.240 ;
        RECT 4.400 213.840 1196.000 215.240 ;
        RECT 4.000 201.640 1196.000 213.840 ;
        RECT 4.000 200.240 1195.600 201.640 ;
        RECT 4.000 194.840 1196.000 200.240 ;
        RECT 4.400 193.440 1196.000 194.840 ;
        RECT 4.000 181.240 1196.000 193.440 ;
        RECT 4.000 179.840 1195.600 181.240 ;
        RECT 4.000 177.840 1196.000 179.840 ;
        RECT 4.400 176.440 1196.000 177.840 ;
        RECT 4.000 160.840 1196.000 176.440 ;
        RECT 4.000 159.440 1195.600 160.840 ;
        RECT 4.000 157.440 1196.000 159.440 ;
        RECT 4.400 156.040 1196.000 157.440 ;
        RECT 4.000 143.840 1196.000 156.040 ;
        RECT 4.000 142.440 1195.600 143.840 ;
        RECT 4.000 137.040 1196.000 142.440 ;
        RECT 4.400 135.640 1196.000 137.040 ;
        RECT 4.000 123.440 1196.000 135.640 ;
        RECT 4.000 122.040 1195.600 123.440 ;
        RECT 4.000 120.040 1196.000 122.040 ;
        RECT 4.400 118.640 1196.000 120.040 ;
        RECT 4.000 103.040 1196.000 118.640 ;
        RECT 4.000 101.640 1195.600 103.040 ;
        RECT 4.000 99.640 1196.000 101.640 ;
        RECT 4.400 98.240 1196.000 99.640 ;
        RECT 4.000 86.040 1196.000 98.240 ;
        RECT 4.000 84.640 1195.600 86.040 ;
        RECT 4.000 79.240 1196.000 84.640 ;
        RECT 4.400 77.840 1196.000 79.240 ;
        RECT 4.000 65.640 1196.000 77.840 ;
        RECT 4.000 64.240 1195.600 65.640 ;
        RECT 4.000 62.240 1196.000 64.240 ;
        RECT 4.400 60.840 1196.000 62.240 ;
        RECT 4.000 45.240 1196.000 60.840 ;
        RECT 4.000 43.840 1195.600 45.240 ;
        RECT 4.000 41.840 1196.000 43.840 ;
        RECT 4.400 40.440 1196.000 41.840 ;
        RECT 4.000 28.240 1196.000 40.440 ;
        RECT 4.000 26.840 1195.600 28.240 ;
        RECT 4.000 21.440 1196.000 26.840 ;
        RECT 4.400 20.040 1196.000 21.440 ;
        RECT 4.000 7.840 1196.000 20.040 ;
        RECT 4.000 6.975 1195.600 7.840 ;
      LAYER met4 ;
        RECT 9.990 11.735 20.640 787.945 ;
        RECT 23.040 11.735 45.640 787.945 ;
        RECT 48.040 476.860 70.640 787.945 ;
        RECT 73.040 476.860 95.640 787.945 ;
        RECT 98.040 476.860 120.640 787.945 ;
        RECT 123.040 476.860 145.640 787.945 ;
        RECT 148.040 476.860 170.640 787.945 ;
        RECT 173.040 476.860 195.640 787.945 ;
        RECT 198.040 476.860 220.640 787.945 ;
        RECT 223.040 476.860 245.640 787.945 ;
        RECT 248.040 476.860 270.640 787.945 ;
        RECT 273.040 476.860 295.640 787.945 ;
        RECT 298.040 476.860 320.640 787.945 ;
        RECT 323.040 476.860 345.640 787.945 ;
        RECT 348.040 476.860 370.640 787.945 ;
        RECT 373.040 476.860 395.640 787.945 ;
        RECT 398.040 476.860 420.640 787.945 ;
        RECT 423.040 476.860 445.640 787.945 ;
        RECT 448.040 476.860 470.640 787.945 ;
        RECT 473.040 476.860 495.640 787.945 ;
        RECT 498.040 476.860 520.640 787.945 ;
        RECT 523.040 476.860 545.640 787.945 ;
        RECT 548.040 476.860 570.640 787.945 ;
        RECT 48.040 70.640 570.640 476.860 ;
        RECT 48.040 11.735 70.640 70.640 ;
        RECT 73.040 11.735 95.640 70.640 ;
        RECT 98.040 11.735 120.640 70.640 ;
        RECT 123.040 11.735 145.640 70.640 ;
        RECT 148.040 11.735 170.640 70.640 ;
        RECT 173.040 11.735 195.640 70.640 ;
        RECT 198.040 11.735 220.640 70.640 ;
        RECT 223.040 11.735 245.640 70.640 ;
        RECT 248.040 11.735 270.640 70.640 ;
        RECT 273.040 11.735 295.640 70.640 ;
        RECT 298.040 11.735 320.640 70.640 ;
        RECT 323.040 11.735 345.640 70.640 ;
        RECT 348.040 11.735 370.640 70.640 ;
        RECT 373.040 11.735 395.640 70.640 ;
        RECT 398.040 11.735 420.640 70.640 ;
        RECT 423.040 11.735 445.640 70.640 ;
        RECT 448.040 11.735 470.640 70.640 ;
        RECT 473.040 11.735 495.640 70.640 ;
        RECT 498.040 11.735 520.640 70.640 ;
        RECT 523.040 11.735 545.640 70.640 ;
        RECT 548.040 11.735 570.640 70.640 ;
        RECT 573.040 11.735 595.640 787.945 ;
        RECT 598.040 11.735 620.640 787.945 ;
        RECT 623.040 11.735 645.640 787.945 ;
        RECT 648.040 11.735 670.640 787.945 ;
        RECT 673.040 11.735 695.640 787.945 ;
        RECT 698.040 11.735 720.640 787.945 ;
        RECT 723.040 11.735 745.640 787.945 ;
        RECT 748.040 11.735 770.640 787.945 ;
        RECT 773.040 11.735 795.640 787.945 ;
        RECT 798.040 11.735 820.640 787.945 ;
        RECT 823.040 11.735 845.640 787.945 ;
        RECT 848.040 11.735 870.640 787.945 ;
        RECT 873.040 11.735 895.640 787.945 ;
        RECT 898.040 11.735 920.640 787.945 ;
        RECT 923.040 11.735 945.640 787.945 ;
        RECT 948.040 11.735 970.640 787.945 ;
        RECT 973.040 11.735 995.640 787.945 ;
        RECT 998.040 11.735 1020.640 787.945 ;
        RECT 1023.040 11.735 1045.640 787.945 ;
        RECT 1048.040 11.735 1070.640 787.945 ;
        RECT 1073.040 11.735 1095.640 787.945 ;
        RECT 1098.040 11.735 1120.640 787.945 ;
        RECT 1123.040 11.735 1145.640 787.945 ;
        RECT 1148.040 11.735 1170.640 787.945 ;
        RECT 1173.040 11.735 1180.490 787.945 ;
      LAYER met5 ;
        RECT 9.780 412.640 1180.700 475.100 ;
        RECT 9.780 336.050 1180.700 407.840 ;
        RECT 9.780 259.460 1180.700 331.250 ;
        RECT 9.780 182.870 1180.700 254.660 ;
        RECT 9.780 106.280 1180.700 178.070 ;
        RECT 9.780 72.300 1180.700 101.480 ;
  END
END core_sram
END LIBRARY

