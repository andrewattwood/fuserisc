VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wb_mem_split
  CLASS BLOCK ;
  FOREIGN wb_mem_split ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 150.000 ;
  PIN core_a_data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END core_a_data_addr_o[0]
  PIN core_a_data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 146.000 271.770 150.000 ;
    END
  END core_a_data_addr_o[1]
  PIN core_a_data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 146.000 218.870 150.000 ;
    END
  END core_a_data_addr_o[2]
  PIN core_a_data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END core_a_data_addr_o[3]
  PIN core_a_data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END core_a_data_addr_o[4]
  PIN core_a_data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 146.000 149.870 150.000 ;
    END
  END core_a_data_addr_o[5]
  PIN core_a_data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 146.000 53.270 150.000 ;
    END
  END core_a_data_addr_o[6]
  PIN core_a_data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END core_a_data_addr_o[7]
  PIN core_a_data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 146.000 276.370 150.000 ;
    END
  END core_a_data_addr_o[8]
  PIN core_a_data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 47.640 300.000 48.240 ;
    END
  END core_a_data_addr_o[9]
  PIN core_a_data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END core_a_data_be_o[0]
  PIN core_a_data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 146.000 119.970 150.000 ;
    END
  END core_a_data_be_o[1]
  PIN core_a_data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 146.000 69.370 150.000 ;
    END
  END core_a_data_be_o[2]
  PIN core_a_data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 95.240 300.000 95.840 ;
    END
  END core_a_data_be_o[3]
  PIN core_a_data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END core_a_data_rdata_i[0]
  PIN core_a_data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END core_a_data_rdata_i[10]
  PIN core_a_data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 112.240 300.000 112.840 ;
    END
  END core_a_data_rdata_i[11]
  PIN core_a_data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END core_a_data_rdata_i[12]
  PIN core_a_data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END core_a_data_rdata_i[13]
  PIN core_a_data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END core_a_data_rdata_i[14]
  PIN core_a_data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 146.000 260.270 150.000 ;
    END
  END core_a_data_rdata_i[15]
  PIN core_a_data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 146.000 290.170 150.000 ;
    END
  END core_a_data_rdata_i[16]
  PIN core_a_data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 13.640 300.000 14.240 ;
    END
  END core_a_data_rdata_i[17]
  PIN core_a_data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 132.640 300.000 133.240 ;
    END
  END core_a_data_rdata_i[18]
  PIN core_a_data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END core_a_data_rdata_i[19]
  PIN core_a_data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END core_a_data_rdata_i[1]
  PIN core_a_data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END core_a_data_rdata_i[20]
  PIN core_a_data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END core_a_data_rdata_i[21]
  PIN core_a_data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END core_a_data_rdata_i[22]
  PIN core_a_data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 146.000 142.970 150.000 ;
    END
  END core_a_data_rdata_i[23]
  PIN core_a_data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END core_a_data_rdata_i[24]
  PIN core_a_data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END core_a_data_rdata_i[25]
  PIN core_a_data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END core_a_data_rdata_i[26]
  PIN core_a_data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 146.000 159.070 150.000 ;
    END
  END core_a_data_rdata_i[27]
  PIN core_a_data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END core_a_data_rdata_i[28]
  PIN core_a_data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 146.000 207.370 150.000 ;
    END
  END core_a_data_rdata_i[29]
  PIN core_a_data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 146.000 60.170 150.000 ;
    END
  END core_a_data_rdata_i[2]
  PIN core_a_data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 146.000 193.570 150.000 ;
    END
  END core_a_data_rdata_i[30]
  PIN core_a_data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 146.000 133.770 150.000 ;
    END
  END core_a_data_rdata_i[31]
  PIN core_a_data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 146.000 78.570 150.000 ;
    END
  END core_a_data_rdata_i[3]
  PIN core_a_data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END core_a_data_rdata_i[4]
  PIN core_a_data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 71.440 300.000 72.040 ;
    END
  END core_a_data_rdata_i[5]
  PIN core_a_data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END core_a_data_rdata_i[6]
  PIN core_a_data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END core_a_data_rdata_i[7]
  PIN core_a_data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 146.000 225.770 150.000 ;
    END
  END core_a_data_rdata_i[8]
  PIN core_a_data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END core_a_data_rdata_i[9]
  PIN core_a_data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 146.000 122.270 150.000 ;
    END
  END core_a_data_req_o
  PIN core_a_data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END core_a_data_rvalid_i
  PIN core_a_data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END core_a_data_wdata_o[0]
  PIN core_a_data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END core_a_data_wdata_o[10]
  PIN core_a_data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END core_a_data_wdata_o[11]
  PIN core_a_data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 146.000 177.470 150.000 ;
    END
  END core_a_data_wdata_o[12]
  PIN core_a_data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 146.000 48.670 150.000 ;
    END
  END core_a_data_wdata_o[13]
  PIN core_a_data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 146.000 62.470 150.000 ;
    END
  END core_a_data_wdata_o[14]
  PIN core_a_data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 146.000 216.570 150.000 ;
    END
  END core_a_data_wdata_o[15]
  PIN core_a_data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 146.000 232.670 150.000 ;
    END
  END core_a_data_wdata_o[16]
  PIN core_a_data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 81.640 300.000 82.240 ;
    END
  END core_a_data_wdata_o[17]
  PIN core_a_data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 146.000 96.970 150.000 ;
    END
  END core_a_data_wdata_o[18]
  PIN core_a_data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END core_a_data_wdata_o[19]
  PIN core_a_data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 146.000 274.070 150.000 ;
    END
  END core_a_data_wdata_o[1]
  PIN core_a_data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 4.000 ;
    END
  END core_a_data_wdata_o[20]
  PIN core_a_data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 146.000 287.870 150.000 ;
    END
  END core_a_data_wdata_o[21]
  PIN core_a_data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 146.000 16.470 150.000 ;
    END
  END core_a_data_wdata_o[22]
  PIN core_a_data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END core_a_data_wdata_o[23]
  PIN core_a_data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 51.040 300.000 51.640 ;
    END
  END core_a_data_wdata_o[24]
  PIN core_a_data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END core_a_data_wdata_o[25]
  PIN core_a_data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END core_a_data_wdata_o[26]
  PIN core_a_data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 98.640 300.000 99.240 ;
    END
  END core_a_data_wdata_o[27]
  PIN core_a_data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 146.000 129.170 150.000 ;
    END
  END core_a_data_wdata_o[28]
  PIN core_a_data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 146.000 186.670 150.000 ;
    END
  END core_a_data_wdata_o[29]
  PIN core_a_data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END core_a_data_wdata_o[2]
  PIN core_a_data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END core_a_data_wdata_o[30]
  PIN core_a_data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 146.000 228.070 150.000 ;
    END
  END core_a_data_wdata_o[31]
  PIN core_a_data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END core_a_data_wdata_o[3]
  PIN core_a_data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END core_a_data_wdata_o[4]
  PIN core_a_data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END core_a_data_wdata_o[5]
  PIN core_a_data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END core_a_data_wdata_o[6]
  PIN core_a_data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END core_a_data_wdata_o[7]
  PIN core_a_data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 146.000 244.170 150.000 ;
    END
  END core_a_data_wdata_o[8]
  PIN core_a_data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 146.000 90.070 150.000 ;
    END
  END core_a_data_wdata_o[9]
  PIN core_a_data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 40.840 300.000 41.440 ;
    END
  END core_a_data_we_o
  PIN core_b_data_addr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END core_b_data_addr_o[0]
  PIN core_b_data_addr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 146.000 161.370 150.000 ;
    END
  END core_b_data_addr_o[1]
  PIN core_b_data_addr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 146.000 14.170 150.000 ;
    END
  END core_b_data_addr_o[2]
  PIN core_b_data_addr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END core_b_data_addr_o[3]
  PIN core_b_data_addr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 146.000 280.970 150.000 ;
    END
  END core_b_data_addr_o[4]
  PIN core_b_data_addr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 146.000 184.370 150.000 ;
    END
  END core_b_data_addr_o[5]
  PIN core_b_data_addr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END core_b_data_addr_o[6]
  PIN core_b_data_addr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END core_b_data_addr_o[7]
  PIN core_b_data_addr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END core_b_data_addr_o[8]
  PIN core_b_data_addr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END core_b_data_addr_o[9]
  PIN core_b_data_be_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END core_b_data_be_o[0]
  PIN core_b_data_be_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END core_b_data_be_o[1]
  PIN core_b_data_be_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.690 146.000 27.970 150.000 ;
    END
  END core_b_data_be_o[2]
  PIN core_b_data_be_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END core_b_data_be_o[3]
  PIN core_b_data_rdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END core_b_data_rdata_i[0]
  PIN core_b_data_rdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END core_b_data_rdata_i[10]
  PIN core_b_data_rdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END core_b_data_rdata_i[11]
  PIN core_b_data_rdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 146.000 85.470 150.000 ;
    END
  END core_b_data_rdata_i[12]
  PIN core_b_data_rdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 146.000 267.170 150.000 ;
    END
  END core_b_data_rdata_i[13]
  PIN core_b_data_rdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 146.000 168.270 150.000 ;
    END
  END core_b_data_rdata_i[14]
  PIN core_b_data_rdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END core_b_data_rdata_i[15]
  PIN core_b_data_rdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END core_b_data_rdata_i[16]
  PIN core_b_data_rdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 129.240 300.000 129.840 ;
    END
  END core_b_data_rdata_i[17]
  PIN core_b_data_rdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END core_b_data_rdata_i[18]
  PIN core_b_data_rdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 146.000 200.470 150.000 ;
    END
  END core_b_data_rdata_i[19]
  PIN core_b_data_rdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 146.000 4.970 150.000 ;
    END
  END core_b_data_rdata_i[1]
  PIN core_b_data_rdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 10.240 300.000 10.840 ;
    END
  END core_b_data_rdata_i[20]
  PIN core_b_data_rdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 20.440 300.000 21.040 ;
    END
  END core_b_data_rdata_i[21]
  PIN core_b_data_rdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 146.000 182.070 150.000 ;
    END
  END core_b_data_rdata_i[22]
  PIN core_b_data_rdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 88.440 300.000 89.040 ;
    END
  END core_b_data_rdata_i[23]
  PIN core_b_data_rdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 146.000 64.770 150.000 ;
    END
  END core_b_data_rdata_i[24]
  PIN core_b_data_rdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END core_b_data_rdata_i[25]
  PIN core_b_data_rdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 146.000 234.970 150.000 ;
    END
  END core_b_data_rdata_i[26]
  PIN core_b_data_rdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 146.000 23.370 150.000 ;
    END
  END core_b_data_rdata_i[27]
  PIN core_b_data_rdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END core_b_data_rdata_i[28]
  PIN core_b_data_rdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END core_b_data_rdata_i[29]
  PIN core_b_data_rdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END core_b_data_rdata_i[2]
  PIN core_b_data_rdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END core_b_data_rdata_i[30]
  PIN core_b_data_rdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 146.000 55.570 150.000 ;
    END
  END core_b_data_rdata_i[31]
  PIN core_b_data_rdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END core_b_data_rdata_i[3]
  PIN core_b_data_rdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 146.000 241.870 150.000 ;
    END
  END core_b_data_rdata_i[4]
  PIN core_b_data_rdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END core_b_data_rdata_i[5]
  PIN core_b_data_rdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END core_b_data_rdata_i[6]
  PIN core_b_data_rdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 23.840 300.000 24.440 ;
    END
  END core_b_data_rdata_i[7]
  PIN core_b_data_rdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 146.000 170.570 150.000 ;
    END
  END core_b_data_rdata_i[8]
  PIN core_b_data_rdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 105.440 300.000 106.040 ;
    END
  END core_b_data_rdata_i[9]
  PIN core_b_data_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 146.000 264.870 150.000 ;
    END
  END core_b_data_req_o
  PIN core_b_data_rvalid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 146.000 257.970 150.000 ;
    END
  END core_b_data_rvalid_i
  PIN core_b_data_wdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END core_b_data_wdata_o[0]
  PIN core_b_data_wdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END core_b_data_wdata_o[10]
  PIN core_b_data_wdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END core_b_data_wdata_o[11]
  PIN core_b_data_wdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END core_b_data_wdata_o[12]
  PIN core_b_data_wdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 146.000 251.070 150.000 ;
    END
  END core_b_data_wdata_o[13]
  PIN core_b_data_wdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END core_b_data_wdata_o[14]
  PIN core_b_data_wdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END core_b_data_wdata_o[15]
  PIN core_b_data_wdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END core_b_data_wdata_o[16]
  PIN core_b_data_wdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END core_b_data_wdata_o[17]
  PIN core_b_data_wdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 146.000 103.870 150.000 ;
    END
  END core_b_data_wdata_o[18]
  PIN core_b_data_wdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 146.000 154.470 150.000 ;
    END
  END core_b_data_wdata_o[19]
  PIN core_b_data_wdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 146.000 30.270 150.000 ;
    END
  END core_b_data_wdata_o[1]
  PIN core_b_data_wdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 146.000 138.370 150.000 ;
    END
  END core_b_data_wdata_o[20]
  PIN core_b_data_wdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END core_b_data_wdata_o[21]
  PIN core_b_data_wdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END core_b_data_wdata_o[22]
  PIN core_b_data_wdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 146.000 145.270 150.000 ;
    END
  END core_b_data_wdata_o[23]
  PIN core_b_data_wdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 146.000 113.070 150.000 ;
    END
  END core_b_data_wdata_o[24]
  PIN core_b_data_wdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END core_b_data_wdata_o[25]
  PIN core_b_data_wdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END core_b_data_wdata_o[26]
  PIN core_b_data_wdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 108.840 300.000 109.440 ;
    END
  END core_b_data_wdata_o[27]
  PIN core_b_data_wdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 142.840 300.000 143.440 ;
    END
  END core_b_data_wdata_o[28]
  PIN core_b_data_wdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END core_b_data_wdata_o[29]
  PIN core_b_data_wdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 146.000 248.770 150.000 ;
    END
  END core_b_data_wdata_o[2]
  PIN core_b_data_wdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 146.000 214.270 150.000 ;
    END
  END core_b_data_wdata_o[30]
  PIN core_b_data_wdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END core_b_data_wdata_o[31]
  PIN core_b_data_wdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 146.000 283.270 150.000 ;
    END
  END core_b_data_wdata_o[3]
  PIN core_b_data_wdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 150.000 ;
    END
  END core_b_data_wdata_o[4]
  PIN core_b_data_wdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END core_b_data_wdata_o[5]
  PIN core_b_data_wdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 146.000 223.470 150.000 ;
    END
  END core_b_data_wdata_o[6]
  PIN core_b_data_wdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 146.000 136.070 150.000 ;
    END
  END core_b_data_wdata_o[7]
  PIN core_b_data_wdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 146.000 32.570 150.000 ;
    END
  END core_b_data_wdata_o[8]
  PIN core_b_data_wdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END core_b_data_wdata_o[9]
  PIN core_b_data_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 146.000 255.670 150.000 ;
    END
  END core_b_data_we_o
  PIN wb_data_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 61.240 300.000 61.840 ;
    END
  END wb_data_addr_i[0]
  PIN wb_data_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_data_addr_i[10]
  PIN wb_data_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 146.000 11.870 150.000 ;
    END
  END wb_data_addr_i[1]
  PIN wb_data_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END wb_data_addr_i[2]
  PIN wb_data_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 74.840 300.000 75.440 ;
    END
  END wb_data_addr_i[3]
  PIN wb_data_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wb_data_addr_i[4]
  PIN wb_data_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wb_data_addr_i[5]
  PIN wb_data_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 146.000 37.170 150.000 ;
    END
  END wb_data_addr_i[6]
  PIN wb_data_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END wb_data_addr_i[7]
  PIN wb_data_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 146.000 39.470 150.000 ;
    END
  END wb_data_addr_i[8]
  PIN wb_data_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 4.000 ;
    END
  END wb_data_addr_i[9]
  PIN wb_data_be_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 0.000 278.670 4.000 ;
    END
  END wb_data_be_i[0]
  PIN wb_data_be_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 146.000 44.070 150.000 ;
    END
  END wb_data_be_i[1]
  PIN wb_data_be_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 146.000 87.770 150.000 ;
    END
  END wb_data_be_i[2]
  PIN wb_data_be_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END wb_data_be_i[3]
  PIN wb_data_rdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wb_data_rdata_o[0]
  PIN wb_data_rdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 146.000 73.970 150.000 ;
    END
  END wb_data_rdata_o[10]
  PIN wb_data_rdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 57.840 300.000 58.440 ;
    END
  END wb_data_rdata_o[11]
  PIN wb_data_rdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 146.000 292.470 150.000 ;
    END
  END wb_data_rdata_o[12]
  PIN wb_data_rdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wb_data_rdata_o[13]
  PIN wb_data_rdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END wb_data_rdata_o[14]
  PIN wb_data_rdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wb_data_rdata_o[15]
  PIN wb_data_rdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wb_data_rdata_o[16]
  PIN wb_data_rdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 146.000 198.170 150.000 ;
    END
  END wb_data_rdata_o[17]
  PIN wb_data_rdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 146.000 101.570 150.000 ;
    END
  END wb_data_rdata_o[18]
  PIN wb_data_rdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wb_data_rdata_o[19]
  PIN wb_data_rdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 27.240 300.000 27.840 ;
    END
  END wb_data_rdata_o[1]
  PIN wb_data_rdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 146.000 209.670 150.000 ;
    END
  END wb_data_rdata_o[20]
  PIN wb_data_rdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wb_data_rdata_o[21]
  PIN wb_data_rdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 146.000 7.270 150.000 ;
    END
  END wb_data_rdata_o[22]
  PIN wb_data_rdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wb_data_rdata_o[23]
  PIN wb_data_rdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 146.000 106.170 150.000 ;
    END
  END wb_data_rdata_o[24]
  PIN wb_data_rdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wb_data_rdata_o[25]
  PIN wb_data_rdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 146.000 46.370 150.000 ;
    END
  END wb_data_rdata_o[26]
  PIN wb_data_rdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wb_data_rdata_o[27]
  PIN wb_data_rdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 146.000 21.070 150.000 ;
    END
  END wb_data_rdata_o[28]
  PIN wb_data_rdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END wb_data_rdata_o[29]
  PIN wb_data_rdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 146.000 165.970 150.000 ;
    END
  END wb_data_rdata_o[2]
  PIN wb_data_rdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wb_data_rdata_o[30]
  PIN wb_data_rdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END wb_data_rdata_o[31]
  PIN wb_data_rdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END wb_data_rdata_o[3]
  PIN wb_data_rdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wb_data_rdata_o[4]
  PIN wb_data_rdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END wb_data_rdata_o[5]
  PIN wb_data_rdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wb_data_rdata_o[6]
  PIN wb_data_rdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wb_data_rdata_o[7]
  PIN wb_data_rdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wb_data_rdata_o[8]
  PIN wb_data_rdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 146.000 239.570 150.000 ;
    END
  END wb_data_rdata_o[9]
  PIN wb_data_rvalid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wb_data_rvalid_o
  PIN wb_data_wdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 85.040 300.000 85.640 ;
    END
  END wb_data_wdata_i[0]
  PIN wb_data_wdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END wb_data_wdata_i[10]
  PIN wb_data_wdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 37.440 300.000 38.040 ;
    END
  END wb_data_wdata_i[11]
  PIN wb_data_wdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END wb_data_wdata_i[12]
  PIN wb_data_wdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 146.000 71.670 150.000 ;
    END
  END wb_data_wdata_i[13]
  PIN wb_data_wdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END wb_data_wdata_i[14]
  PIN wb_data_wdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 3.440 300.000 4.040 ;
    END
  END wb_data_wdata_i[15]
  PIN wb_data_wdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END wb_data_wdata_i[16]
  PIN wb_data_wdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 136.040 300.000 136.640 ;
    END
  END wb_data_wdata_i[17]
  PIN wb_data_wdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wb_data_wdata_i[18]
  PIN wb_data_wdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wb_data_wdata_i[19]
  PIN wb_data_wdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 119.040 300.000 119.640 ;
    END
  END wb_data_wdata_i[1]
  PIN wb_data_wdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 146.000 126.870 150.000 ;
    END
  END wb_data_wdata_i[20]
  PIN wb_data_wdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END wb_data_wdata_i[21]
  PIN wb_data_wdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 146.000 117.670 150.000 ;
    END
  END wb_data_wdata_i[22]
  PIN wb_data_wdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 146.000 175.170 150.000 ;
    END
  END wb_data_wdata_i[23]
  PIN wb_data_wdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END wb_data_wdata_i[24]
  PIN wb_data_wdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END wb_data_wdata_i[25]
  PIN wb_data_wdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 146.000 202.770 150.000 ;
    END
  END wb_data_wdata_i[26]
  PIN wb_data_wdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wb_data_wdata_i[27]
  PIN wb_data_wdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 64.640 300.000 65.240 ;
    END
  END wb_data_wdata_i[28]
  PIN wb_data_wdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 146.000 110.770 150.000 ;
    END
  END wb_data_wdata_i[29]
  PIN wb_data_wdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END wb_data_wdata_i[2]
  PIN wb_data_wdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wb_data_wdata_i[30]
  PIN wb_data_wdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 122.440 300.000 123.040 ;
    END
  END wb_data_wdata_i[31]
  PIN wb_data_wdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END wb_data_wdata_i[3]
  PIN wb_data_wdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wb_data_wdata_i[4]
  PIN wb_data_wdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wb_data_wdata_i[5]
  PIN wb_data_wdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.000 34.040 300.000 34.640 ;
    END
  END wb_data_wdata_i[6]
  PIN wb_data_wdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END wb_data_wdata_i[7]
  PIN wb_data_wdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 146.000 152.170 150.000 ;
    END
  END wb_data_wdata_i[8]
  PIN wb_data_wdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 146.000 191.270 150.000 ;
    END
  END wb_data_wdata_i[9]
  PIN wb_data_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wb_data_we_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 146.000 94.670 150.000 ;
    END
  END wbs_cyc_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 146.000 297.070 150.000 ;
    END
  END wbs_stb_i
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 245.520 10.640 247.120 138.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 149.200 10.640 150.800 138.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 52.880 10.640 54.480 138.960 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 116.705 294.400 118.305 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 73.960 294.400 75.560 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 31.215 294.400 32.815 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 197.360 10.640 198.960 138.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.040 10.640 102.640 138.960 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 95.335 294.400 96.935 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 52.585 294.400 54.185 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 8.585 294.400 138.805 ;
      LAYER met1 ;
        RECT 2.370 7.520 297.090 140.720 ;
      LAYER met2 ;
        RECT 2.400 145.720 4.410 146.000 ;
        RECT 5.250 145.720 6.710 146.000 ;
        RECT 7.550 145.720 11.310 146.000 ;
        RECT 12.150 145.720 13.610 146.000 ;
        RECT 14.450 145.720 15.910 146.000 ;
        RECT 16.750 145.720 20.510 146.000 ;
        RECT 21.350 145.720 22.810 146.000 ;
        RECT 23.650 145.720 27.410 146.000 ;
        RECT 28.250 145.720 29.710 146.000 ;
        RECT 30.550 145.720 32.010 146.000 ;
        RECT 32.850 145.720 36.610 146.000 ;
        RECT 37.450 145.720 38.910 146.000 ;
        RECT 39.750 145.720 43.510 146.000 ;
        RECT 44.350 145.720 45.810 146.000 ;
        RECT 46.650 145.720 48.110 146.000 ;
        RECT 48.950 145.720 52.710 146.000 ;
        RECT 53.550 145.720 55.010 146.000 ;
        RECT 55.850 145.720 59.610 146.000 ;
        RECT 60.450 145.720 61.910 146.000 ;
        RECT 62.750 145.720 64.210 146.000 ;
        RECT 65.050 145.720 68.810 146.000 ;
        RECT 69.650 145.720 71.110 146.000 ;
        RECT 71.950 145.720 73.410 146.000 ;
        RECT 74.250 145.720 78.010 146.000 ;
        RECT 78.850 145.720 80.310 146.000 ;
        RECT 81.150 145.720 84.910 146.000 ;
        RECT 85.750 145.720 87.210 146.000 ;
        RECT 88.050 145.720 89.510 146.000 ;
        RECT 90.350 145.720 94.110 146.000 ;
        RECT 94.950 145.720 96.410 146.000 ;
        RECT 97.250 145.720 101.010 146.000 ;
        RECT 101.850 145.720 103.310 146.000 ;
        RECT 104.150 145.720 105.610 146.000 ;
        RECT 106.450 145.720 110.210 146.000 ;
        RECT 111.050 145.720 112.510 146.000 ;
        RECT 113.350 145.720 117.110 146.000 ;
        RECT 117.950 145.720 119.410 146.000 ;
        RECT 120.250 145.720 121.710 146.000 ;
        RECT 122.550 145.720 126.310 146.000 ;
        RECT 127.150 145.720 128.610 146.000 ;
        RECT 129.450 145.720 133.210 146.000 ;
        RECT 134.050 145.720 135.510 146.000 ;
        RECT 136.350 145.720 137.810 146.000 ;
        RECT 138.650 145.720 142.410 146.000 ;
        RECT 143.250 145.720 144.710 146.000 ;
        RECT 145.550 145.720 149.310 146.000 ;
        RECT 150.150 145.720 151.610 146.000 ;
        RECT 152.450 145.720 153.910 146.000 ;
        RECT 154.750 145.720 158.510 146.000 ;
        RECT 159.350 145.720 160.810 146.000 ;
        RECT 161.650 145.720 165.410 146.000 ;
        RECT 166.250 145.720 167.710 146.000 ;
        RECT 168.550 145.720 170.010 146.000 ;
        RECT 170.850 145.720 174.610 146.000 ;
        RECT 175.450 145.720 176.910 146.000 ;
        RECT 177.750 145.720 181.510 146.000 ;
        RECT 182.350 145.720 183.810 146.000 ;
        RECT 184.650 145.720 186.110 146.000 ;
        RECT 186.950 145.720 190.710 146.000 ;
        RECT 191.550 145.720 193.010 146.000 ;
        RECT 193.850 145.720 197.610 146.000 ;
        RECT 198.450 145.720 199.910 146.000 ;
        RECT 200.750 145.720 202.210 146.000 ;
        RECT 203.050 145.720 206.810 146.000 ;
        RECT 207.650 145.720 209.110 146.000 ;
        RECT 209.950 145.720 213.710 146.000 ;
        RECT 214.550 145.720 216.010 146.000 ;
        RECT 216.850 145.720 218.310 146.000 ;
        RECT 219.150 145.720 222.910 146.000 ;
        RECT 223.750 145.720 225.210 146.000 ;
        RECT 226.050 145.720 227.510 146.000 ;
        RECT 228.350 145.720 232.110 146.000 ;
        RECT 232.950 145.720 234.410 146.000 ;
        RECT 235.250 145.720 239.010 146.000 ;
        RECT 239.850 145.720 241.310 146.000 ;
        RECT 242.150 145.720 243.610 146.000 ;
        RECT 244.450 145.720 248.210 146.000 ;
        RECT 249.050 145.720 250.510 146.000 ;
        RECT 251.350 145.720 255.110 146.000 ;
        RECT 255.950 145.720 257.410 146.000 ;
        RECT 258.250 145.720 259.710 146.000 ;
        RECT 260.550 145.720 264.310 146.000 ;
        RECT 265.150 145.720 266.610 146.000 ;
        RECT 267.450 145.720 271.210 146.000 ;
        RECT 272.050 145.720 273.510 146.000 ;
        RECT 274.350 145.720 275.810 146.000 ;
        RECT 276.650 145.720 280.410 146.000 ;
        RECT 281.250 145.720 282.710 146.000 ;
        RECT 283.550 145.720 287.310 146.000 ;
        RECT 288.150 145.720 289.610 146.000 ;
        RECT 290.450 145.720 291.910 146.000 ;
        RECT 292.750 145.720 296.510 146.000 ;
        RECT 2.400 4.280 297.060 145.720 ;
        RECT 2.950 3.555 4.410 4.280 ;
        RECT 5.250 3.555 6.710 4.280 ;
        RECT 7.550 3.555 11.310 4.280 ;
        RECT 12.150 3.555 13.610 4.280 ;
        RECT 14.450 3.555 15.910 4.280 ;
        RECT 16.750 3.555 20.510 4.280 ;
        RECT 21.350 3.555 22.810 4.280 ;
        RECT 23.650 3.555 27.410 4.280 ;
        RECT 28.250 3.555 29.710 4.280 ;
        RECT 30.550 3.555 32.010 4.280 ;
        RECT 32.850 3.555 36.610 4.280 ;
        RECT 37.450 3.555 38.910 4.280 ;
        RECT 39.750 3.555 43.510 4.280 ;
        RECT 44.350 3.555 45.810 4.280 ;
        RECT 46.650 3.555 48.110 4.280 ;
        RECT 48.950 3.555 52.710 4.280 ;
        RECT 53.550 3.555 55.010 4.280 ;
        RECT 55.850 3.555 59.610 4.280 ;
        RECT 60.450 3.555 61.910 4.280 ;
        RECT 62.750 3.555 64.210 4.280 ;
        RECT 65.050 3.555 68.810 4.280 ;
        RECT 69.650 3.555 71.110 4.280 ;
        RECT 71.950 3.555 75.710 4.280 ;
        RECT 76.550 3.555 78.010 4.280 ;
        RECT 78.850 3.555 80.310 4.280 ;
        RECT 81.150 3.555 84.910 4.280 ;
        RECT 85.750 3.555 87.210 4.280 ;
        RECT 88.050 3.555 91.810 4.280 ;
        RECT 92.650 3.555 94.110 4.280 ;
        RECT 94.950 3.555 96.410 4.280 ;
        RECT 97.250 3.555 101.010 4.280 ;
        RECT 101.850 3.555 103.310 4.280 ;
        RECT 104.150 3.555 107.910 4.280 ;
        RECT 108.750 3.555 110.210 4.280 ;
        RECT 111.050 3.555 112.510 4.280 ;
        RECT 113.350 3.555 117.110 4.280 ;
        RECT 117.950 3.555 119.410 4.280 ;
        RECT 120.250 3.555 124.010 4.280 ;
        RECT 124.850 3.555 126.310 4.280 ;
        RECT 127.150 3.555 128.610 4.280 ;
        RECT 129.450 3.555 133.210 4.280 ;
        RECT 134.050 3.555 135.510 4.280 ;
        RECT 136.350 3.555 140.110 4.280 ;
        RECT 140.950 3.555 142.410 4.280 ;
        RECT 143.250 3.555 144.710 4.280 ;
        RECT 145.550 3.555 149.310 4.280 ;
        RECT 150.150 3.555 151.610 4.280 ;
        RECT 152.450 3.555 156.210 4.280 ;
        RECT 157.050 3.555 158.510 4.280 ;
        RECT 159.350 3.555 160.810 4.280 ;
        RECT 161.650 3.555 165.410 4.280 ;
        RECT 166.250 3.555 167.710 4.280 ;
        RECT 168.550 3.555 170.010 4.280 ;
        RECT 170.850 3.555 174.610 4.280 ;
        RECT 175.450 3.555 176.910 4.280 ;
        RECT 177.750 3.555 181.510 4.280 ;
        RECT 182.350 3.555 183.810 4.280 ;
        RECT 184.650 3.555 186.110 4.280 ;
        RECT 186.950 3.555 190.710 4.280 ;
        RECT 191.550 3.555 193.010 4.280 ;
        RECT 193.850 3.555 197.610 4.280 ;
        RECT 198.450 3.555 199.910 4.280 ;
        RECT 200.750 3.555 202.210 4.280 ;
        RECT 203.050 3.555 206.810 4.280 ;
        RECT 207.650 3.555 209.110 4.280 ;
        RECT 209.950 3.555 213.710 4.280 ;
        RECT 214.550 3.555 216.010 4.280 ;
        RECT 216.850 3.555 218.310 4.280 ;
        RECT 219.150 3.555 222.910 4.280 ;
        RECT 223.750 3.555 225.210 4.280 ;
        RECT 226.050 3.555 229.810 4.280 ;
        RECT 230.650 3.555 232.110 4.280 ;
        RECT 232.950 3.555 234.410 4.280 ;
        RECT 235.250 3.555 239.010 4.280 ;
        RECT 239.850 3.555 241.310 4.280 ;
        RECT 242.150 3.555 245.910 4.280 ;
        RECT 246.750 3.555 248.210 4.280 ;
        RECT 249.050 3.555 250.510 4.280 ;
        RECT 251.350 3.555 255.110 4.280 ;
        RECT 255.950 3.555 257.410 4.280 ;
        RECT 258.250 3.555 262.010 4.280 ;
        RECT 262.850 3.555 264.310 4.280 ;
        RECT 265.150 3.555 266.610 4.280 ;
        RECT 267.450 3.555 271.210 4.280 ;
        RECT 272.050 3.555 273.510 4.280 ;
        RECT 274.350 3.555 278.110 4.280 ;
        RECT 278.950 3.555 280.410 4.280 ;
        RECT 281.250 3.555 282.710 4.280 ;
        RECT 283.550 3.555 287.310 4.280 ;
        RECT 288.150 3.555 289.610 4.280 ;
        RECT 290.450 3.555 294.210 4.280 ;
        RECT 295.050 3.555 296.510 4.280 ;
      LAYER met3 ;
        RECT 4.400 142.440 295.600 143.305 ;
        RECT 4.000 140.440 296.000 142.440 ;
        RECT 4.400 139.040 296.000 140.440 ;
        RECT 4.000 137.040 296.000 139.040 ;
        RECT 4.400 135.640 295.600 137.040 ;
        RECT 4.000 133.640 296.000 135.640 ;
        RECT 4.000 132.240 295.600 133.640 ;
        RECT 4.000 130.240 296.000 132.240 ;
        RECT 4.400 128.840 295.600 130.240 ;
        RECT 4.000 126.840 296.000 128.840 ;
        RECT 4.400 125.440 296.000 126.840 ;
        RECT 4.000 123.440 296.000 125.440 ;
        RECT 4.000 122.040 295.600 123.440 ;
        RECT 4.000 120.040 296.000 122.040 ;
        RECT 4.400 118.640 295.600 120.040 ;
        RECT 4.000 116.640 296.000 118.640 ;
        RECT 4.400 115.240 296.000 116.640 ;
        RECT 4.000 113.240 296.000 115.240 ;
        RECT 4.400 111.840 295.600 113.240 ;
        RECT 4.000 109.840 296.000 111.840 ;
        RECT 4.000 108.440 295.600 109.840 ;
        RECT 4.000 106.440 296.000 108.440 ;
        RECT 4.400 105.040 295.600 106.440 ;
        RECT 4.000 103.040 296.000 105.040 ;
        RECT 4.400 101.640 296.000 103.040 ;
        RECT 4.000 99.640 296.000 101.640 ;
        RECT 4.000 98.240 295.600 99.640 ;
        RECT 4.000 96.240 296.000 98.240 ;
        RECT 4.400 94.840 295.600 96.240 ;
        RECT 4.000 92.840 296.000 94.840 ;
        RECT 4.400 91.440 296.000 92.840 ;
        RECT 4.000 89.440 296.000 91.440 ;
        RECT 4.400 88.040 295.600 89.440 ;
        RECT 4.000 86.040 296.000 88.040 ;
        RECT 4.000 84.640 295.600 86.040 ;
        RECT 4.000 82.640 296.000 84.640 ;
        RECT 4.400 81.240 295.600 82.640 ;
        RECT 4.000 79.240 296.000 81.240 ;
        RECT 4.400 77.840 296.000 79.240 ;
        RECT 4.000 75.840 296.000 77.840 ;
        RECT 4.000 74.440 295.600 75.840 ;
        RECT 4.000 72.440 296.000 74.440 ;
        RECT 4.400 71.040 295.600 72.440 ;
        RECT 4.000 69.040 296.000 71.040 ;
        RECT 4.400 67.640 296.000 69.040 ;
        RECT 4.000 65.640 296.000 67.640 ;
        RECT 4.400 64.240 295.600 65.640 ;
        RECT 4.000 62.240 296.000 64.240 ;
        RECT 4.000 60.840 295.600 62.240 ;
        RECT 4.000 58.840 296.000 60.840 ;
        RECT 4.400 57.440 295.600 58.840 ;
        RECT 4.000 55.440 296.000 57.440 ;
        RECT 4.400 54.040 296.000 55.440 ;
        RECT 4.000 52.040 296.000 54.040 ;
        RECT 4.000 50.640 295.600 52.040 ;
        RECT 4.000 48.640 296.000 50.640 ;
        RECT 4.400 47.240 295.600 48.640 ;
        RECT 4.000 45.240 296.000 47.240 ;
        RECT 4.400 43.840 296.000 45.240 ;
        RECT 4.000 41.840 296.000 43.840 ;
        RECT 4.400 40.440 295.600 41.840 ;
        RECT 4.000 38.440 296.000 40.440 ;
        RECT 4.000 37.040 295.600 38.440 ;
        RECT 4.000 35.040 296.000 37.040 ;
        RECT 4.400 33.640 295.600 35.040 ;
        RECT 4.000 31.640 296.000 33.640 ;
        RECT 4.400 30.240 296.000 31.640 ;
        RECT 4.000 28.240 296.000 30.240 ;
        RECT 4.000 26.840 295.600 28.240 ;
        RECT 4.000 24.840 296.000 26.840 ;
        RECT 4.400 23.440 295.600 24.840 ;
        RECT 4.000 21.440 296.000 23.440 ;
        RECT 4.400 20.040 295.600 21.440 ;
        RECT 4.000 18.040 296.000 20.040 ;
        RECT 4.400 16.640 296.000 18.040 ;
        RECT 4.000 14.640 296.000 16.640 ;
        RECT 4.000 13.240 295.600 14.640 ;
        RECT 4.000 11.240 296.000 13.240 ;
        RECT 4.400 9.840 295.600 11.240 ;
        RECT 4.000 7.840 296.000 9.840 ;
        RECT 4.400 6.440 296.000 7.840 ;
        RECT 4.000 4.440 296.000 6.440 ;
        RECT 4.000 3.575 295.600 4.440 ;
      LAYER met5 ;
        RECT 5.520 77.160 294.400 93.735 ;
        RECT 5.520 55.785 294.400 72.360 ;
        RECT 5.520 34.415 294.400 50.985 ;
  END
END wb_mem_split
END LIBRARY

