magic
tech sky130A
magscale 1 2
timestamp 1623315978
<< nwell >>
rect 1066 117221 178886 117542
rect 1066 116133 178886 116699
rect 1066 115045 178886 115611
rect 1066 113957 178886 114523
rect 1066 112869 178886 113435
rect 1066 111781 178886 112347
rect 1066 110693 178886 111259
rect 1066 109605 178886 110171
rect 1066 108517 178886 109083
rect 1066 107429 178886 107995
rect 1066 106341 178886 106907
rect 1066 105253 178886 105819
rect 1066 104165 178886 104731
rect 1066 103077 178886 103643
rect 1066 101989 178886 102555
rect 1066 100901 178886 101467
rect 1066 99813 178886 100379
rect 1066 98725 178886 99291
rect 1066 97637 178886 98203
rect 1066 96549 178886 97115
rect 1066 95461 178886 96027
rect 1066 94373 178886 94939
rect 1066 93285 178886 93851
rect 1066 92197 178886 92763
rect 1066 91109 178886 91675
rect 1066 90021 178886 90587
rect 1066 88933 178886 89499
rect 1066 87845 178886 88411
rect 1066 86757 178886 87323
rect 1066 85669 178886 86235
rect 1066 84581 178886 85147
rect 1066 83493 178886 84059
rect 1066 82405 178886 82971
rect 1066 81317 178886 81883
rect 1066 80229 178886 80795
rect 1066 79141 178886 79707
rect 1066 78053 178886 78619
rect 1066 76965 178886 77531
rect 1066 75877 178886 76443
rect 1066 74789 178886 75355
rect 1066 73701 178886 74267
rect 1066 72613 178886 73179
rect 1066 71525 178886 72091
rect 1066 70437 178886 71003
rect 1066 69349 178886 69915
rect 1066 68261 178886 68827
rect 1066 67173 178886 67739
rect 1066 66085 178886 66651
rect 1066 64997 178886 65563
rect 1066 63909 178886 64475
rect 1066 62821 178886 63387
rect 1066 61733 178886 62299
rect 1066 60645 178886 61211
rect 1066 59557 178886 60123
rect 1066 58469 178886 59035
rect 1066 57381 178886 57947
rect 1066 56293 178886 56859
rect 1066 55205 178886 55771
rect 1066 54117 178886 54683
rect 1066 53029 178886 53595
rect 1066 51941 178886 52507
rect 1066 50853 178886 51419
rect 1066 49765 178886 50331
rect 1066 48677 178886 49243
rect 1066 47589 178886 48155
rect 1066 46501 178886 47067
rect 1066 45413 178886 45979
rect 1066 44325 178886 44891
rect 1066 43237 178886 43803
rect 1066 42149 178886 42715
rect 1066 41061 178886 41627
rect 1066 39973 178886 40539
rect 1066 38885 178886 39451
rect 1066 37797 178886 38363
rect 1066 36709 178886 37275
rect 1066 35621 178886 36187
rect 1066 34533 178886 35099
rect 1066 33445 178886 34011
rect 1066 32357 178886 32923
rect 1066 31269 178886 31835
rect 1066 30181 178886 30747
rect 1066 29093 178886 29659
rect 1066 28005 178886 28571
rect 1066 26917 178886 27483
rect 1066 25829 178886 26395
rect 1066 24741 178886 25307
rect 1066 23653 178886 24219
rect 1066 22565 178886 23131
rect 1066 21477 178886 22043
rect 1066 20389 178886 20955
rect 1066 19301 178886 19867
rect 1066 18213 178886 18779
rect 1066 17125 178886 17691
rect 1066 16037 178886 16603
rect 1066 14949 178886 15515
rect 1066 13861 178886 14427
rect 1066 12773 178886 13339
rect 1066 11685 178886 12251
rect 1066 10597 178886 11163
rect 1066 9509 178886 10075
rect 1066 8421 178886 8987
rect 1066 7333 178886 7899
rect 1066 6245 178886 6811
rect 1066 5157 178886 5723
rect 1066 4069 178886 4635
rect 1066 2981 178886 3547
rect 1066 2138 178886 2459
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 1104 2128 178848 117552
<< metal2 >>
rect 7470 0 7526 800
rect 22466 0 22522 800
rect 37462 0 37518 800
rect 52458 0 52514 800
rect 67454 0 67510 800
rect 82450 0 82506 800
rect 97446 0 97502 800
rect 112442 0 112498 800
rect 127438 0 127494 800
rect 142434 0 142490 800
rect 157430 0 157486 800
rect 172426 0 172482 800
<< obsm2 >>
rect 4220 856 175978 117552
rect 4220 800 7414 856
rect 7582 800 22410 856
rect 22578 800 37406 856
rect 37574 800 52402 856
rect 52570 800 67398 856
rect 67566 800 82394 856
rect 82562 800 97390 856
rect 97558 800 112386 856
rect 112554 800 127382 856
rect 127550 800 142378 856
rect 142546 800 157374 856
rect 157542 800 172370 856
rect 172538 800 175978 856
<< metal3 >>
rect 179200 59984 180000 60104
<< obsm3 >>
rect 4208 60184 179200 117537
rect 4208 59904 179120 60184
rect 4208 2143 179200 59904
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 57283 10099 65568 47701
rect 66048 10099 66228 47701
rect 66708 10099 66888 47701
rect 67368 10099 67548 47701
rect 68028 10099 80928 47701
rect 81408 10099 81588 47701
rect 82068 10099 82248 47701
rect 82728 10099 82908 47701
rect 83388 10099 86789 47701
<< labels >>
rlabel metal3 s 179200 59984 180000 60104 6 clk
port 1 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_data_out[0]
port 2 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[10]
port 3 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 la_data_out[1]
port 4 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 la_data_out[2]
port 5 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 la_data_out[3]
port 6 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[4]
port 7 nsew signal output
rlabel metal2 s 97446 0 97502 800 6 la_data_out[5]
port 8 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 la_data_out[6]
port 9 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 la_data_out[7]
port 10 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[8]
port 11 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 la_data_out[9]
port 12 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 wb_rst_i
port 13 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 14 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 16 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 18 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 19 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 20 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 21 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 22 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 23 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 24 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 25 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 26 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 27 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 28 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 29 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 30 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 31 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 32 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 33 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 34 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 35 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 36 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 37 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 38 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 39 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 40 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 41 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 42 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 43 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 44 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 45 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 46 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 47 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 48 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 49 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 50 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 51 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 52 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 53 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 54 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 55 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 56 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 57 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 58 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 59 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 60 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 61 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 8738460
string GDS_START 611748
<< end >>

