VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1199.740 BY 1210.460 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END clk_i
  PIN debug_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 918.040 1199.740 918.640 ;
    END
  END debug_req_i
  PIN eFPGA_delay_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.490 1206.460 1168.770 1210.460 ;
    END
  END eFPGA_delay_o[0]
  PIN eFPGA_delay_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END eFPGA_delay_o[1]
  PIN eFPGA_delay_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END eFPGA_delay_o[2]
  PIN eFPGA_delay_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 1206.460 862.870 1210.460 ;
    END
  END eFPGA_delay_o[3]
  PIN eFPGA_en_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 1206.460 444.270 1210.460 ;
    END
  END eFPGA_en_o
  PIN eFPGA_fpga_done_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 0.000 517.870 4.000 ;
    END
  END eFPGA_fpga_done_i
  PIN eFPGA_operand_a_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 873.840 1199.740 874.440 ;
    END
  END eFPGA_operand_a_o[0]
  PIN eFPGA_operand_a_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END eFPGA_operand_a_o[10]
  PIN eFPGA_operand_a_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END eFPGA_operand_a_o[11]
  PIN eFPGA_operand_a_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 0.000 1173.370 4.000 ;
    END
  END eFPGA_operand_a_o[12]
  PIN eFPGA_operand_a_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END eFPGA_operand_a_o[13]
  PIN eFPGA_operand_a_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 0.000 740.970 4.000 ;
    END
  END eFPGA_operand_a_o[14]
  PIN eFPGA_operand_a_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 1206.460 1141.170 1210.460 ;
    END
  END eFPGA_operand_a_o[15]
  PIN eFPGA_operand_a_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 523.640 1199.740 524.240 ;
    END
  END eFPGA_operand_a_o[16]
  PIN eFPGA_operand_a_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 1206.460 1016.970 1210.460 ;
    END
  END eFPGA_operand_a_o[17]
  PIN eFPGA_operand_a_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END eFPGA_operand_a_o[18]
  PIN eFPGA_operand_a_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END eFPGA_operand_a_o[19]
  PIN eFPGA_operand_a_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 1206.460 80.870 1210.460 ;
    END
  END eFPGA_operand_a_o[1]
  PIN eFPGA_operand_a_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END eFPGA_operand_a_o[20]
  PIN eFPGA_operand_a_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 792.240 1199.740 792.840 ;
    END
  END eFPGA_operand_a_o[21]
  PIN eFPGA_operand_a_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 173.440 1199.740 174.040 ;
    END
  END eFPGA_operand_a_o[22]
  PIN eFPGA_operand_a_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 234.640 1199.740 235.240 ;
    END
  END eFPGA_operand_a_o[23]
  PIN eFPGA_operand_a_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END eFPGA_operand_a_o[24]
  PIN eFPGA_operand_a_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END eFPGA_operand_a_o[25]
  PIN eFPGA_operand_a_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1020.040 1199.740 1020.640 ;
    END
  END eFPGA_operand_a_o[26]
  PIN eFPGA_operand_a_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 979.240 1199.740 979.840 ;
    END
  END eFPGA_operand_a_o[27]
  PIN eFPGA_operand_a_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END eFPGA_operand_a_o[28]
  PIN eFPGA_operand_a_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.990 1206.460 835.270 1210.460 ;
    END
  END eFPGA_operand_a_o[29]
  PIN eFPGA_operand_a_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 319.640 1199.740 320.240 ;
    END
  END eFPGA_operand_a_o[2]
  PIN eFPGA_operand_a_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 0.000 1007.770 4.000 ;
    END
  END eFPGA_operand_a_o[30]
  PIN eFPGA_operand_a_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 1206.460 722.570 1210.460 ;
    END
  END eFPGA_operand_a_o[31]
  PIN eFPGA_operand_a_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.490 0.000 1145.770 4.000 ;
    END
  END eFPGA_operand_a_o[3]
  PIN eFPGA_operand_a_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 1206.460 1113.570 1210.460 ;
    END
  END eFPGA_operand_a_o[4]
  PIN eFPGA_operand_a_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END eFPGA_operand_a_o[5]
  PIN eFPGA_operand_a_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END eFPGA_operand_a_o[6]
  PIN eFPGA_operand_a_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END eFPGA_operand_a_o[7]
  PIN eFPGA_operand_a_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 0.000 867.470 4.000 ;
    END
  END eFPGA_operand_a_o[8]
  PIN eFPGA_operand_a_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 1206.460 554.670 1210.460 ;
    END
  END eFPGA_operand_a_o[9]
  PIN eFPGA_operand_b_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1060.840 1199.740 1061.440 ;
    END
  END eFPGA_operand_b_o[0]
  PIN eFPGA_operand_b_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1101.640 1199.740 1102.240 ;
    END
  END eFPGA_operand_b_o[10]
  PIN eFPGA_operand_b_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 1206.460 653.570 1210.460 ;
    END
  END eFPGA_operand_b_o[11]
  PIN eFPGA_operand_b_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END eFPGA_operand_b_o[12]
  PIN eFPGA_operand_b_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END eFPGA_operand_b_o[13]
  PIN eFPGA_operand_b_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 1206.460 750.170 1210.460 ;
    END
  END eFPGA_operand_b_o[14]
  PIN eFPGA_operand_b_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 1206.460 430.470 1210.460 ;
    END
  END eFPGA_operand_b_o[15]
  PIN eFPGA_operand_b_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END eFPGA_operand_b_o[16]
  PIN eFPGA_operand_b_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END eFPGA_operand_b_o[17]
  PIN eFPGA_operand_b_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.890 0.000 1118.170 4.000 ;
    END
  END eFPGA_operand_b_o[18]
  PIN eFPGA_operand_b_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 1206.460 207.370 1210.460 ;
    END
  END eFPGA_operand_b_o[19]
  PIN eFPGA_operand_b_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END eFPGA_operand_b_o[1]
  PIN eFPGA_operand_b_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END eFPGA_operand_b_o[20]
  PIN eFPGA_operand_b_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 584.840 1199.740 585.440 ;
    END
  END eFPGA_operand_b_o[21]
  PIN eFPGA_operand_b_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 1206.460 791.570 1210.460 ;
    END
  END eFPGA_operand_b_o[22]
  PIN eFPGA_operand_b_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 1206.460 568.470 1210.460 ;
    END
  END eFPGA_operand_b_o[23]
  PIN eFPGA_operand_b_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END eFPGA_operand_b_o[24]
  PIN eFPGA_operand_b_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.840 4.000 602.440 ;
    END
  END eFPGA_operand_b_o[25]
  PIN eFPGA_operand_b_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 0.000 812.270 4.000 ;
    END
  END eFPGA_operand_b_o[26]
  PIN eFPGA_operand_b_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END eFPGA_operand_b_o[27]
  PIN eFPGA_operand_b_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 1206.460 149.870 1210.460 ;
    END
  END eFPGA_operand_b_o[28]
  PIN eFPGA_operand_b_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.590 0.000 839.870 4.000 ;
    END
  END eFPGA_operand_b_o[29]
  PIN eFPGA_operand_b_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 731.040 1199.740 731.640 ;
    END
  END eFPGA_operand_b_o[2]
  PIN eFPGA_operand_b_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 340.040 1199.740 340.640 ;
    END
  END eFPGA_operand_b_o[30]
  PIN eFPGA_operand_b_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 0.000 448.870 4.000 ;
    END
  END eFPGA_operand_b_o[31]
  PIN eFPGA_operand_b_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END eFPGA_operand_b_o[3]
  PIN eFPGA_operand_b_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END eFPGA_operand_b_o[4]
  PIN eFPGA_operand_b_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END eFPGA_operand_b_o[5]
  PIN eFPGA_operand_b_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 1206.460 777.770 1210.460 ;
    END
  END eFPGA_operand_b_o[6]
  PIN eFPGA_operand_b_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END eFPGA_operand_b_o[7]
  PIN eFPGA_operand_b_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.590 1206.460 931.870 1210.460 ;
    END
  END eFPGA_operand_b_o[8]
  PIN eFPGA_operand_b_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END eFPGA_operand_b_o[9]
  PIN eFPGA_operator_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END eFPGA_operator_o[0]
  PIN eFPGA_operator_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 710.640 1199.740 711.240 ;
    END
  END eFPGA_operator_o[1]
  PIN eFPGA_result_a_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 1206.460 290.170 1210.460 ;
    END
  END eFPGA_result_a_i[0]
  PIN eFPGA_result_a_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END eFPGA_result_a_i[10]
  PIN eFPGA_result_a_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 1206.460 763.970 1210.460 ;
    END
  END eFPGA_result_a_i[11]
  PIN eFPGA_result_a_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END eFPGA_result_a_i[12]
  PIN eFPGA_result_a_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1081.240 1199.740 1081.840 ;
    END
  END eFPGA_result_a_i[13]
  PIN eFPGA_result_a_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END eFPGA_result_a_i[14]
  PIN eFPGA_result_a_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END eFPGA_result_a_i[15]
  PIN eFPGA_result_a_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 917.790 1206.460 918.070 1210.460 ;
    END
  END eFPGA_result_a_i[16]
  PIN eFPGA_result_a_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END eFPGA_result_a_i[17]
  PIN eFPGA_result_a_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 1206.460 276.370 1210.460 ;
    END
  END eFPGA_result_a_i[18]
  PIN eFPGA_result_a_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END eFPGA_result_a_i[19]
  PIN eFPGA_result_a_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END eFPGA_result_a_i[1]
  PIN eFPGA_result_a_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END eFPGA_result_a_i[20]
  PIN eFPGA_result_a_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 0.000 476.470 4.000 ;
    END
  END eFPGA_result_a_i[21]
  PIN eFPGA_result_a_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 91.840 1199.740 92.440 ;
    END
  END eFPGA_result_a_i[22]
  PIN eFPGA_result_a_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END eFPGA_result_a_i[23]
  PIN eFPGA_result_a_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END eFPGA_result_a_i[24]
  PIN eFPGA_result_a_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END eFPGA_result_a_i[25]
  PIN eFPGA_result_a_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END eFPGA_result_a_i[26]
  PIN eFPGA_result_a_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END eFPGA_result_a_i[27]
  PIN eFPGA_result_a_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 1206.460 598.370 1210.460 ;
    END
  END eFPGA_result_a_i[28]
  PIN eFPGA_result_a_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END eFPGA_result_a_i[29]
  PIN eFPGA_result_a_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END eFPGA_result_a_i[2]
  PIN eFPGA_result_a_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 938.440 1199.740 939.040 ;
    END
  END eFPGA_result_a_i[30]
  PIN eFPGA_result_a_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 1206.460 582.270 1210.460 ;
    END
  END eFPGA_result_a_i[31]
  PIN eFPGA_result_a_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 1206.460 945.670 1210.460 ;
    END
  END eFPGA_result_a_i[3]
  PIN eFPGA_result_a_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 1206.460 513.270 1210.460 ;
    END
  END eFPGA_result_a_i[4]
  PIN eFPGA_result_a_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END eFPGA_result_a_i[5]
  PIN eFPGA_result_a_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END eFPGA_result_a_i[6]
  PIN eFPGA_result_a_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END eFPGA_result_a_i[7]
  PIN eFPGA_result_a_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.690 1206.460 1085.970 1210.460 ;
    END
  END eFPGA_result_a_i[8]
  PIN eFPGA_result_a_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 1206.460 527.070 1210.460 ;
    END
  END eFPGA_result_a_i[9]
  PIN eFPGA_result_b_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 0.000 922.670 4.000 ;
    END
  END eFPGA_result_b_i[0]
  PIN eFPGA_result_b_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 564.440 1199.740 565.040 ;
    END
  END eFPGA_result_b_i[10]
  PIN eFPGA_result_b_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 1206.460 1003.170 1210.460 ;
    END
  END eFPGA_result_b_i[11]
  PIN eFPGA_result_b_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 503.240 1199.740 503.840 ;
    END
  END eFPGA_result_b_i[12]
  PIN eFPGA_result_b_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 1206.460 499.470 1210.460 ;
    END
  END eFPGA_result_b_i[13]
  PIN eFPGA_result_b_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END eFPGA_result_b_i[14]
  PIN eFPGA_result_b_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 1206.460 39.470 1210.460 ;
    END
  END eFPGA_result_b_i[15]
  PIN eFPGA_result_b_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1122.040 1199.740 1122.640 ;
    END
  END eFPGA_result_b_i[16]
  PIN eFPGA_result_b_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END eFPGA_result_b_i[17]
  PIN eFPGA_result_b_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END eFPGA_result_b_i[18]
  PIN eFPGA_result_b_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 1206.460 904.270 1210.460 ;
    END
  END eFPGA_result_b_i[19]
  PIN eFPGA_result_b_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 0.000 908.870 4.000 ;
    END
  END eFPGA_result_b_i[1]
  PIN eFPGA_result_b_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END eFPGA_result_b_i[20]
  PIN eFPGA_result_b_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 1206.460 694.970 1210.460 ;
    END
  END eFPGA_result_b_i[21]
  PIN eFPGA_result_b_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.240 4.000 1200.840 ;
    END
  END eFPGA_result_b_i[22]
  PIN eFPGA_result_b_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END eFPGA_result_b_i[23]
  PIN eFPGA_result_b_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END eFPGA_result_b_i[24]
  PIN eFPGA_result_b_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END eFPGA_result_b_i[25]
  PIN eFPGA_result_b_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 1206.460 625.970 1210.460 ;
    END
  END eFPGA_result_b_i[26]
  PIN eFPGA_result_b_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END eFPGA_result_b_i[27]
  PIN eFPGA_result_b_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 958.840 1199.740 959.440 ;
    END
  END eFPGA_result_b_i[28]
  PIN eFPGA_result_b_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 999.640 1199.740 1000.240 ;
    END
  END eFPGA_result_b_i[29]
  PIN eFPGA_result_b_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 1206.460 234.970 1210.460 ;
    END
  END eFPGA_result_b_i[2]
  PIN eFPGA_result_b_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 1206.460 53.270 1210.460 ;
    END
  END eFPGA_result_b_i[30]
  PIN eFPGA_result_b_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 0.000 1035.370 4.000 ;
    END
  END eFPGA_result_b_i[31]
  PIN eFPGA_result_b_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.490 1206.460 1099.770 1210.460 ;
    END
  END eFPGA_result_b_i[3]
  PIN eFPGA_result_b_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1040.440 1199.740 1041.040 ;
    END
  END eFPGA_result_b_i[4]
  PIN eFPGA_result_b_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END eFPGA_result_b_i[5]
  PIN eFPGA_result_b_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END eFPGA_result_b_i[6]
  PIN eFPGA_result_b_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 51.040 1199.740 51.640 ;
    END
  END eFPGA_result_b_i[7]
  PIN eFPGA_result_b_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 0.000 881.270 4.000 ;
    END
  END eFPGA_result_b_i[8]
  PIN eFPGA_result_b_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 1206.460 485.670 1210.460 ;
    END
  END eFPGA_result_b_i[9]
  PIN eFPGA_result_c_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 1206.460 667.370 1210.460 ;
    END
  END eFPGA_result_c_i[0]
  PIN eFPGA_result_c_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.190 1206.460 890.470 1210.460 ;
    END
  END eFPGA_result_c_i[10]
  PIN eFPGA_result_c_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END eFPGA_result_c_i[11]
  PIN eFPGA_result_c_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END eFPGA_result_c_i[12]
  PIN eFPGA_result_c_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 0.000 1049.170 4.000 ;
    END
  END eFPGA_result_c_i[13]
  PIN eFPGA_result_c_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 1206.460 736.370 1210.460 ;
    END
  END eFPGA_result_c_i[14]
  PIN eFPGA_result_c_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 214.240 1199.740 214.840 ;
    END
  END eFPGA_result_c_i[15]
  PIN eFPGA_result_c_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END eFPGA_result_c_i[16]
  PIN eFPGA_result_c_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END eFPGA_result_c_i[17]
  PIN eFPGA_result_c_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END eFPGA_result_c_i[18]
  PIN eFPGA_result_c_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 0.000 964.070 4.000 ;
    END
  END eFPGA_result_c_i[19]
  PIN eFPGA_result_c_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.490 0.000 1076.770 4.000 ;
    END
  END eFPGA_result_c_i[1]
  PIN eFPGA_result_c_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 132.640 1199.740 133.240 ;
    END
  END eFPGA_result_c_i[20]
  PIN eFPGA_result_c_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 275.440 1199.740 276.040 ;
    END
  END eFPGA_result_c_i[21]
  PIN eFPGA_result_c_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END eFPGA_result_c_i[22]
  PIN eFPGA_result_c_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END eFPGA_result_c_i[23]
  PIN eFPGA_result_c_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END eFPGA_result_c_i[24]
  PIN eFPGA_result_c_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END eFPGA_result_c_i[25]
  PIN eFPGA_result_c_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END eFPGA_result_c_i[26]
  PIN eFPGA_result_c_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END eFPGA_result_c_i[27]
  PIN eFPGA_result_c_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 1206.460 359.170 1210.460 ;
    END
  END eFPGA_result_c_i[28]
  PIN eFPGA_result_c_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 1206.460 163.670 1210.460 ;
    END
  END eFPGA_result_c_i[29]
  PIN eFPGA_result_c_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.790 0.000 895.070 4.000 ;
    END
  END eFPGA_result_c_i[2]
  PIN eFPGA_result_c_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.890 1206.460 1072.170 1210.460 ;
    END
  END eFPGA_result_c_i[30]
  PIN eFPGA_result_c_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END eFPGA_result_c_i[31]
  PIN eFPGA_result_c_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 1206.460 122.270 1210.460 ;
    END
  END eFPGA_result_c_i[3]
  PIN eFPGA_result_c_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 0.000 713.370 4.000 ;
    END
  END eFPGA_result_c_i[4]
  PIN eFPGA_result_c_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 482.840 1199.740 483.440 ;
    END
  END eFPGA_result_c_i[5]
  PIN eFPGA_result_c_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 1206.460 681.170 1210.460 ;
    END
  END eFPGA_result_c_i[6]
  PIN eFPGA_result_c_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.290 1206.460 1182.570 1210.460 ;
    END
  END eFPGA_result_c_i[7]
  PIN eFPGA_result_c_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END eFPGA_result_c_i[8]
  PIN eFPGA_result_c_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 421.640 1199.740 422.240 ;
    END
  END eFPGA_result_c_i[9]
  PIN eFPGA_write_strobe_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 1206.460 386.770 1210.460 ;
    END
  END eFPGA_write_strobe_o
  PIN ext_data_addr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1159.290 0.000 1159.570 4.000 ;
    END
  END ext_data_addr_i[0]
  PIN ext_data_addr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1183.240 1199.740 1183.840 ;
    END
  END ext_data_addr_i[10]
  PIN ext_data_addr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END ext_data_addr_i[11]
  PIN ext_data_addr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END ext_data_addr_i[12]
  PIN ext_data_addr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END ext_data_addr_i[13]
  PIN ext_data_addr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 0.000 1131.970 4.000 ;
    END
  END ext_data_addr_i[14]
  PIN ext_data_addr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END ext_data_addr_i[15]
  PIN ext_data_addr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END ext_data_addr_i[16]
  PIN ext_data_addr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 1206.460 402.870 1210.460 ;
    END
  END ext_data_addr_i[17]
  PIN ext_data_addr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.290 0.000 1021.570 4.000 ;
    END
  END ext_data_addr_i[18]
  PIN ext_data_addr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END ext_data_addr_i[19]
  PIN ext_data_addr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 605.240 1199.740 605.840 ;
    END
  END ext_data_addr_i[1]
  PIN ext_data_addr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 1206.460 94.670 1210.460 ;
    END
  END ext_data_addr_i[20]
  PIN ext_data_addr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 833.040 1199.740 833.640 ;
    END
  END ext_data_addr_i[21]
  PIN ext_data_addr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 1206.460 345.370 1210.460 ;
    END
  END ext_data_addr_i[22]
  PIN ext_data_addr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 295.840 1199.740 296.440 ;
    END
  END ext_data_addr_i[23]
  PIN ext_data_addr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.690 0.000 1062.970 4.000 ;
    END
  END ext_data_addr_i[24]
  PIN ext_data_addr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.090 0.000 253.370 4.000 ;
    END
  END ext_data_addr_i[25]
  PIN ext_data_addr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1162.840 1199.740 1163.440 ;
    END
  END ext_data_addr_i[26]
  PIN ext_data_addr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 1206.460 248.770 1210.460 ;
    END
  END ext_data_addr_i[27]
  PIN ext_data_addr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 1206.460 849.070 1210.460 ;
    END
  END ext_data_addr_i[28]
  PIN ext_data_addr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 1206.460 959.470 1210.460 ;
    END
  END ext_data_addr_i[29]
  PIN ext_data_addr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 991.390 0.000 991.670 4.000 ;
    END
  END ext_data_addr_i[2]
  PIN ext_data_addr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 1206.460 416.670 1210.460 ;
    END
  END ext_data_addr_i[30]
  PIN ext_data_addr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 1206.460 540.870 1210.460 ;
    END
  END ext_data_addr_i[31]
  PIN ext_data_addr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 1206.460 303.970 1210.460 ;
    END
  END ext_data_addr_i[3]
  PIN ext_data_addr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.090 1206.460 1127.370 1210.460 ;
    END
  END ext_data_addr_i[4]
  PIN ext_data_addr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 153.040 1199.740 153.640 ;
    END
  END ext_data_addr_i[5]
  PIN ext_data_addr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 1206.460 221.170 1210.460 ;
    END
  END ext_data_addr_i[6]
  PIN ext_data_addr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 1206.460 372.970 1210.460 ;
    END
  END ext_data_addr_i[7]
  PIN ext_data_addr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END ext_data_addr_i[8]
  PIN ext_data_addr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END ext_data_addr_i[9]
  PIN ext_data_be_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 1206.460 136.070 1210.460 ;
    END
  END ext_data_be_i[0]
  PIN ext_data_be_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 112.240 1199.740 112.840 ;
    END
  END ext_data_be_i[1]
  PIN ext_data_be_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 1206.460 67.070 1210.460 ;
    END
  END ext_data_be_i[2]
  PIN ext_data_be_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END ext_data_be_i[3]
  PIN ext_data_rdata_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END ext_data_rdata_o[0]
  PIN ext_data_rdata_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.090 0.000 1104.370 4.000 ;
    END
  END ext_data_rdata_o[10]
  PIN ext_data_rdata_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END ext_data_rdata_o[11]
  PIN ext_data_rdata_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 751.440 1199.740 752.040 ;
    END
  END ext_data_rdata_o[12]
  PIN ext_data_rdata_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 1206.460 612.170 1210.460 ;
    END
  END ext_data_rdata_o[13]
  PIN ext_data_rdata_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 812.640 1199.740 813.240 ;
    END
  END ext_data_rdata_o[14]
  PIN ext_data_rdata_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END ext_data_rdata_o[15]
  PIN ext_data_rdata_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END ext_data_rdata_o[16]
  PIN ext_data_rdata_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END ext_data_rdata_o[17]
  PIN ext_data_rdata_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END ext_data_rdata_o[18]
  PIN ext_data_rdata_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END ext_data_rdata_o[19]
  PIN ext_data_rdata_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 669.840 1199.740 670.440 ;
    END
  END ext_data_rdata_o[1]
  PIN ext_data_rdata_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END ext_data_rdata_o[20]
  PIN ext_data_rdata_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 30.640 1199.740 31.240 ;
    END
  END ext_data_rdata_o[21]
  PIN ext_data_rdata_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END ext_data_rdata_o[22]
  PIN ext_data_rdata_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 360.440 1199.740 361.040 ;
    END
  END ext_data_rdata_o[23]
  PIN ext_data_rdata_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END ext_data_rdata_o[24]
  PIN ext_data_rdata_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 972.990 1206.460 973.270 1210.460 ;
    END
  END ext_data_rdata_o[25]
  PIN ext_data_rdata_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END ext_data_rdata_o[26]
  PIN ext_data_rdata_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 1206.460 191.270 1210.460 ;
    END
  END ext_data_rdata_o[27]
  PIN ext_data_rdata_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.190 0.000 936.470 4.000 ;
    END
  END ext_data_rdata_o[28]
  PIN ext_data_rdata_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.090 1206.460 1196.370 1210.460 ;
    END
  END ext_data_rdata_o[29]
  PIN ext_data_rdata_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END ext_data_rdata_o[2]
  PIN ext_data_rdata_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.890 0.000 1187.170 4.000 ;
    END
  END ext_data_rdata_o[30]
  PIN ext_data_rdata_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 1206.460 108.470 1210.460 ;
    END
  END ext_data_rdata_o[31]
  PIN ext_data_rdata_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 193.840 1199.740 194.440 ;
    END
  END ext_data_rdata_o[3]
  PIN ext_data_rdata_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 690.240 1199.740 690.840 ;
    END
  END ext_data_rdata_o[4]
  PIN ext_data_rdata_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END ext_data_rdata_o[5]
  PIN ext_data_rdata_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 380.840 1199.740 381.440 ;
    END
  END ext_data_rdata_o[6]
  PIN ext_data_rdata_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END ext_data_rdata_o[7]
  PIN ext_data_rdata_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.390 1206.460 876.670 1210.460 ;
    END
  END ext_data_rdata_o[8]
  PIN ext_data_rdata_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 1206.460 821.470 1210.460 ;
    END
  END ext_data_rdata_o[9]
  PIN ext_data_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 1206.460 11.870 1210.460 ;
    END
  END ext_data_req_i
  PIN ext_data_rvalid_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 1206.460 331.570 1210.460 ;
    END
  END ext_data_rvalid_o
  PIN ext_data_wdata_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 1206.460 177.470 1210.460 ;
    END
  END ext_data_wdata_i[0]
  PIN ext_data_wdata_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 1142.440 1199.740 1143.040 ;
    END
  END ext_data_wdata_i[10]
  PIN ext_data_wdata_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END ext_data_wdata_i[11]
  PIN ext_data_wdata_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 544.040 1199.740 544.640 ;
    END
  END ext_data_wdata_i[12]
  PIN ext_data_wdata_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 401.240 1199.740 401.840 ;
    END
  END ext_data_wdata_i[13]
  PIN ext_data_wdata_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END ext_data_wdata_i[14]
  PIN ext_data_wdata_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END ext_data_wdata_i[15]
  PIN ext_data_wdata_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END ext_data_wdata_i[16]
  PIN ext_data_wdata_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.590 0.000 977.870 4.000 ;
    END
  END ext_data_wdata_i[17]
  PIN ext_data_wdata_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 649.440 1199.740 650.040 ;
    END
  END ext_data_wdata_i[18]
  PIN ext_data_wdata_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.490 1206.460 1030.770 1210.460 ;
    END
  END ext_data_wdata_i[19]
  PIN ext_data_wdata_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END ext_data_wdata_i[1]
  PIN ext_data_wdata_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END ext_data_wdata_i[20]
  PIN ext_data_wdata_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 853.440 1199.740 854.040 ;
    END
  END ext_data_wdata_i[21]
  PIN ext_data_wdata_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END ext_data_wdata_i[22]
  PIN ext_data_wdata_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END ext_data_wdata_i[23]
  PIN ext_data_wdata_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.690 1206.460 1154.970 1210.460 ;
    END
  END ext_data_wdata_i[24]
  PIN ext_data_wdata_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 1206.460 807.670 1210.460 ;
    END
  END ext_data_wdata_i[25]
  PIN ext_data_wdata_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 1206.460 639.770 1210.460 ;
    END
  END ext_data_wdata_i[26]
  PIN ext_data_wdata_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 0.000 1090.570 4.000 ;
    END
  END ext_data_wdata_i[27]
  PIN ext_data_wdata_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 629.040 1199.740 629.640 ;
    END
  END ext_data_wdata_i[28]
  PIN ext_data_wdata_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.040 4.000 663.640 ;
    END
  END ext_data_wdata_i[29]
  PIN ext_data_wdata_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 462.440 1199.740 463.040 ;
    END
  END ext_data_wdata_i[2]
  PIN ext_data_wdata_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 1206.460 1058.370 1210.460 ;
    END
  END ext_data_wdata_i[30]
  PIN ext_data_wdata_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 0.000 421.270 4.000 ;
    END
  END ext_data_wdata_i[31]
  PIN ext_data_wdata_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 1206.460 262.570 1210.460 ;
    END
  END ext_data_wdata_i[3]
  PIN ext_data_wdata_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END ext_data_wdata_i[4]
  PIN ext_data_wdata_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 894.240 1199.740 894.840 ;
    END
  END ext_data_wdata_i[5]
  PIN ext_data_wdata_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END ext_data_wdata_i[6]
  PIN ext_data_wdata_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 1206.460 25.670 1210.460 ;
    END
  END ext_data_wdata_i[7]
  PIN ext_data_wdata_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 394.440 4.000 395.040 ;
    END
  END ext_data_wdata_i[8]
  PIN ext_data_wdata_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 1206.460 317.770 1210.460 ;
    END
  END ext_data_wdata_i[9]
  PIN ext_data_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END ext_data_we_i
  PIN fetch_enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 6.840 1199.740 7.440 ;
    END
  END fetch_enable_i
  PIN irq_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 1206.460 458.070 1210.460 ;
    END
  END irq_ack_o
  PIN irq_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END irq_i
  PIN irq_id_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 1206.460 987.070 1210.460 ;
    END
  END irq_id_i[0]
  PIN irq_id_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END irq_id_i[1]
  PIN irq_id_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.590 1206.460 471.870 1210.460 ;
    END
  END irq_id_i[2]
  PIN irq_id_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 442.040 1199.740 442.640 ;
    END
  END irq_id_i[3]
  PIN irq_id_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 71.440 1199.740 72.040 ;
    END
  END irq_id_i[4]
  PIN irq_id_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 1206.460 708.770 1210.460 ;
    END
  END irq_id_o[0]
  PIN irq_id_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 255.040 1199.740 255.640 ;
    END
  END irq_id_o[1]
  PIN irq_id_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.290 1206.460 1044.570 1210.460 ;
    END
  END irq_id_o[2]
  PIN irq_id_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END irq_id_o[3]
  PIN irq_id_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1195.740 771.840 1199.740 772.440 ;
    END
  END irq_id_o[4]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END reset
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1171.040 10.640 1172.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1121.040 10.640 1122.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1071.040 10.640 1072.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1021.040 10.640 1022.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 971.040 10.640 972.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 921.040 10.640 922.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 871.040 10.640 872.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 821.040 10.640 822.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 771.040 10.640 772.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 721.040 10.640 722.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 671.040 10.640 672.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 621.040 10.640 622.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 502.260 572.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 502.260 522.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 502.260 472.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 502.260 422.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 502.260 372.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 502.260 322.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 502.260 272.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 502.260 222.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 502.260 172.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 502.260 122.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 71.040 10.640 72.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1199.760 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 571.040 10.640 572.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 521.040 10.640 522.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 471.040 10.640 472.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 421.040 10.640 422.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 371.040 10.640 372.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 321.040 10.640 322.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 271.040 10.640 272.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 221.040 10.640 222.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 171.040 10.640 172.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 121.040 10.640 122.640 95.240 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 1098.750 1194.160 1100.350 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 945.570 1194.160 947.170 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 792.390 1194.160 793.990 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 639.210 1194.160 640.810 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 1194.160 487.630 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 1194.160 334.450 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 1194.160 181.270 ;
    END
  END VPWR
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 1194.160 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1146.040 10.640 1147.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1096.040 10.640 1097.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1046.040 10.640 1047.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 996.040 10.640 997.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 946.040 10.640 947.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 896.040 10.640 897.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 846.040 10.640 847.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 796.040 10.640 797.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 746.040 10.640 747.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 696.040 10.640 697.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 646.040 10.640 647.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 596.040 10.640 597.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 502.260 547.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 502.260 497.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 502.260 447.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 502.260 397.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 502.260 347.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 502.260 297.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 502.260 247.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 502.260 197.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 502.260 147.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 502.260 97.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 46.040 10.640 47.640 1199.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 546.040 10.640 547.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 496.040 10.640 497.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 446.040 10.640 447.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 396.040 10.640 397.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 346.040 10.640 347.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 296.040 10.640 297.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 246.040 10.640 247.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 196.040 10.640 197.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 146.040 10.640 147.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.040 10.640 97.640 95.240 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1175.340 1194.160 1176.940 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 1022.160 1194.160 1023.760 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 868.980 1194.160 870.580 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 715.800 1194.160 717.400 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 1194.160 564.220 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 1194.160 411.040 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 1194.160 257.860 ;
    END
  END VGND
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 1194.160 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1199.605 ;
      LAYER met1 ;
        RECT 2.370 8.540 1196.390 1201.520 ;
      LAYER met2 ;
        RECT 2.400 1206.180 11.310 1206.460 ;
        RECT 12.150 1206.180 25.110 1206.460 ;
        RECT 25.950 1206.180 38.910 1206.460 ;
        RECT 39.750 1206.180 52.710 1206.460 ;
        RECT 53.550 1206.180 66.510 1206.460 ;
        RECT 67.350 1206.180 80.310 1206.460 ;
        RECT 81.150 1206.180 94.110 1206.460 ;
        RECT 94.950 1206.180 107.910 1206.460 ;
        RECT 108.750 1206.180 121.710 1206.460 ;
        RECT 122.550 1206.180 135.510 1206.460 ;
        RECT 136.350 1206.180 149.310 1206.460 ;
        RECT 150.150 1206.180 163.110 1206.460 ;
        RECT 163.950 1206.180 176.910 1206.460 ;
        RECT 177.750 1206.180 190.710 1206.460 ;
        RECT 191.550 1206.180 206.810 1206.460 ;
        RECT 207.650 1206.180 220.610 1206.460 ;
        RECT 221.450 1206.180 234.410 1206.460 ;
        RECT 235.250 1206.180 248.210 1206.460 ;
        RECT 249.050 1206.180 262.010 1206.460 ;
        RECT 262.850 1206.180 275.810 1206.460 ;
        RECT 276.650 1206.180 289.610 1206.460 ;
        RECT 290.450 1206.180 303.410 1206.460 ;
        RECT 304.250 1206.180 317.210 1206.460 ;
        RECT 318.050 1206.180 331.010 1206.460 ;
        RECT 331.850 1206.180 344.810 1206.460 ;
        RECT 345.650 1206.180 358.610 1206.460 ;
        RECT 359.450 1206.180 372.410 1206.460 ;
        RECT 373.250 1206.180 386.210 1206.460 ;
        RECT 387.050 1206.180 402.310 1206.460 ;
        RECT 403.150 1206.180 416.110 1206.460 ;
        RECT 416.950 1206.180 429.910 1206.460 ;
        RECT 430.750 1206.180 443.710 1206.460 ;
        RECT 444.550 1206.180 457.510 1206.460 ;
        RECT 458.350 1206.180 471.310 1206.460 ;
        RECT 472.150 1206.180 485.110 1206.460 ;
        RECT 485.950 1206.180 498.910 1206.460 ;
        RECT 499.750 1206.180 512.710 1206.460 ;
        RECT 513.550 1206.180 526.510 1206.460 ;
        RECT 527.350 1206.180 540.310 1206.460 ;
        RECT 541.150 1206.180 554.110 1206.460 ;
        RECT 554.950 1206.180 567.910 1206.460 ;
        RECT 568.750 1206.180 581.710 1206.460 ;
        RECT 582.550 1206.180 597.810 1206.460 ;
        RECT 598.650 1206.180 611.610 1206.460 ;
        RECT 612.450 1206.180 625.410 1206.460 ;
        RECT 626.250 1206.180 639.210 1206.460 ;
        RECT 640.050 1206.180 653.010 1206.460 ;
        RECT 653.850 1206.180 666.810 1206.460 ;
        RECT 667.650 1206.180 680.610 1206.460 ;
        RECT 681.450 1206.180 694.410 1206.460 ;
        RECT 695.250 1206.180 708.210 1206.460 ;
        RECT 709.050 1206.180 722.010 1206.460 ;
        RECT 722.850 1206.180 735.810 1206.460 ;
        RECT 736.650 1206.180 749.610 1206.460 ;
        RECT 750.450 1206.180 763.410 1206.460 ;
        RECT 764.250 1206.180 777.210 1206.460 ;
        RECT 778.050 1206.180 791.010 1206.460 ;
        RECT 791.850 1206.180 807.110 1206.460 ;
        RECT 807.950 1206.180 820.910 1206.460 ;
        RECT 821.750 1206.180 834.710 1206.460 ;
        RECT 835.550 1206.180 848.510 1206.460 ;
        RECT 849.350 1206.180 862.310 1206.460 ;
        RECT 863.150 1206.180 876.110 1206.460 ;
        RECT 876.950 1206.180 889.910 1206.460 ;
        RECT 890.750 1206.180 903.710 1206.460 ;
        RECT 904.550 1206.180 917.510 1206.460 ;
        RECT 918.350 1206.180 931.310 1206.460 ;
        RECT 932.150 1206.180 945.110 1206.460 ;
        RECT 945.950 1206.180 958.910 1206.460 ;
        RECT 959.750 1206.180 972.710 1206.460 ;
        RECT 973.550 1206.180 986.510 1206.460 ;
        RECT 987.350 1206.180 1002.610 1206.460 ;
        RECT 1003.450 1206.180 1016.410 1206.460 ;
        RECT 1017.250 1206.180 1030.210 1206.460 ;
        RECT 1031.050 1206.180 1044.010 1206.460 ;
        RECT 1044.850 1206.180 1057.810 1206.460 ;
        RECT 1058.650 1206.180 1071.610 1206.460 ;
        RECT 1072.450 1206.180 1085.410 1206.460 ;
        RECT 1086.250 1206.180 1099.210 1206.460 ;
        RECT 1100.050 1206.180 1113.010 1206.460 ;
        RECT 1113.850 1206.180 1126.810 1206.460 ;
        RECT 1127.650 1206.180 1140.610 1206.460 ;
        RECT 1141.450 1206.180 1154.410 1206.460 ;
        RECT 1155.250 1206.180 1168.210 1206.460 ;
        RECT 1169.050 1206.180 1182.010 1206.460 ;
        RECT 1182.850 1206.180 1195.810 1206.460 ;
        RECT 2.400 4.280 1196.360 1206.180 ;
        RECT 2.950 4.000 15.910 4.280 ;
        RECT 16.750 4.000 29.710 4.280 ;
        RECT 30.550 4.000 43.510 4.280 ;
        RECT 44.350 4.000 57.310 4.280 ;
        RECT 58.150 4.000 71.110 4.280 ;
        RECT 71.950 4.000 84.910 4.280 ;
        RECT 85.750 4.000 98.710 4.280 ;
        RECT 99.550 4.000 112.510 4.280 ;
        RECT 113.350 4.000 126.310 4.280 ;
        RECT 127.150 4.000 140.110 4.280 ;
        RECT 140.950 4.000 153.910 4.280 ;
        RECT 154.750 4.000 167.710 4.280 ;
        RECT 168.550 4.000 181.510 4.280 ;
        RECT 182.350 4.000 195.310 4.280 ;
        RECT 196.150 4.000 211.410 4.280 ;
        RECT 212.250 4.000 225.210 4.280 ;
        RECT 226.050 4.000 239.010 4.280 ;
        RECT 239.850 4.000 252.810 4.280 ;
        RECT 253.650 4.000 266.610 4.280 ;
        RECT 267.450 4.000 280.410 4.280 ;
        RECT 281.250 4.000 294.210 4.280 ;
        RECT 295.050 4.000 308.010 4.280 ;
        RECT 308.850 4.000 321.810 4.280 ;
        RECT 322.650 4.000 335.610 4.280 ;
        RECT 336.450 4.000 349.410 4.280 ;
        RECT 350.250 4.000 363.210 4.280 ;
        RECT 364.050 4.000 377.010 4.280 ;
        RECT 377.850 4.000 390.810 4.280 ;
        RECT 391.650 4.000 406.910 4.280 ;
        RECT 407.750 4.000 420.710 4.280 ;
        RECT 421.550 4.000 434.510 4.280 ;
        RECT 435.350 4.000 448.310 4.280 ;
        RECT 449.150 4.000 462.110 4.280 ;
        RECT 462.950 4.000 475.910 4.280 ;
        RECT 476.750 4.000 489.710 4.280 ;
        RECT 490.550 4.000 503.510 4.280 ;
        RECT 504.350 4.000 517.310 4.280 ;
        RECT 518.150 4.000 531.110 4.280 ;
        RECT 531.950 4.000 544.910 4.280 ;
        RECT 545.750 4.000 558.710 4.280 ;
        RECT 559.550 4.000 572.510 4.280 ;
        RECT 573.350 4.000 586.310 4.280 ;
        RECT 587.150 4.000 600.110 4.280 ;
        RECT 600.950 4.000 616.210 4.280 ;
        RECT 617.050 4.000 630.010 4.280 ;
        RECT 630.850 4.000 643.810 4.280 ;
        RECT 644.650 4.000 657.610 4.280 ;
        RECT 658.450 4.000 671.410 4.280 ;
        RECT 672.250 4.000 685.210 4.280 ;
        RECT 686.050 4.000 699.010 4.280 ;
        RECT 699.850 4.000 712.810 4.280 ;
        RECT 713.650 4.000 726.610 4.280 ;
        RECT 727.450 4.000 740.410 4.280 ;
        RECT 741.250 4.000 754.210 4.280 ;
        RECT 755.050 4.000 768.010 4.280 ;
        RECT 768.850 4.000 781.810 4.280 ;
        RECT 782.650 4.000 795.610 4.280 ;
        RECT 796.450 4.000 811.710 4.280 ;
        RECT 812.550 4.000 825.510 4.280 ;
        RECT 826.350 4.000 839.310 4.280 ;
        RECT 840.150 4.000 853.110 4.280 ;
        RECT 853.950 4.000 866.910 4.280 ;
        RECT 867.750 4.000 880.710 4.280 ;
        RECT 881.550 4.000 894.510 4.280 ;
        RECT 895.350 4.000 908.310 4.280 ;
        RECT 909.150 4.000 922.110 4.280 ;
        RECT 922.950 4.000 935.910 4.280 ;
        RECT 936.750 4.000 949.710 4.280 ;
        RECT 950.550 4.000 963.510 4.280 ;
        RECT 964.350 4.000 977.310 4.280 ;
        RECT 978.150 4.000 991.110 4.280 ;
        RECT 991.950 4.000 1007.210 4.280 ;
        RECT 1008.050 4.000 1021.010 4.280 ;
        RECT 1021.850 4.000 1034.810 4.280 ;
        RECT 1035.650 4.000 1048.610 4.280 ;
        RECT 1049.450 4.000 1062.410 4.280 ;
        RECT 1063.250 4.000 1076.210 4.280 ;
        RECT 1077.050 4.000 1090.010 4.280 ;
        RECT 1090.850 4.000 1103.810 4.280 ;
        RECT 1104.650 4.000 1117.610 4.280 ;
        RECT 1118.450 4.000 1131.410 4.280 ;
        RECT 1132.250 4.000 1145.210 4.280 ;
        RECT 1146.050 4.000 1159.010 4.280 ;
        RECT 1159.850 4.000 1172.810 4.280 ;
        RECT 1173.650 4.000 1186.610 4.280 ;
        RECT 1187.450 4.000 1196.360 4.280 ;
      LAYER met3 ;
        RECT 4.000 1201.240 1195.740 1202.745 ;
        RECT 4.400 1199.840 1195.740 1201.240 ;
        RECT 4.000 1184.240 1195.740 1199.840 ;
        RECT 4.000 1182.840 1195.340 1184.240 ;
        RECT 4.000 1177.440 1195.740 1182.840 ;
        RECT 4.400 1176.040 1195.740 1177.440 ;
        RECT 4.000 1163.840 1195.740 1176.040 ;
        RECT 4.000 1162.440 1195.340 1163.840 ;
        RECT 4.000 1157.040 1195.740 1162.440 ;
        RECT 4.400 1155.640 1195.740 1157.040 ;
        RECT 4.000 1143.440 1195.740 1155.640 ;
        RECT 4.000 1142.040 1195.340 1143.440 ;
        RECT 4.000 1136.640 1195.740 1142.040 ;
        RECT 4.400 1135.240 1195.740 1136.640 ;
        RECT 4.000 1123.040 1195.740 1135.240 ;
        RECT 4.000 1121.640 1195.340 1123.040 ;
        RECT 4.000 1116.240 1195.740 1121.640 ;
        RECT 4.400 1114.840 1195.740 1116.240 ;
        RECT 4.000 1102.640 1195.740 1114.840 ;
        RECT 4.000 1101.240 1195.340 1102.640 ;
        RECT 4.000 1095.840 1195.740 1101.240 ;
        RECT 4.400 1094.440 1195.740 1095.840 ;
        RECT 4.000 1082.240 1195.740 1094.440 ;
        RECT 4.000 1080.840 1195.340 1082.240 ;
        RECT 4.000 1075.440 1195.740 1080.840 ;
        RECT 4.400 1074.040 1195.740 1075.440 ;
        RECT 4.000 1061.840 1195.740 1074.040 ;
        RECT 4.000 1060.440 1195.340 1061.840 ;
        RECT 4.000 1055.040 1195.740 1060.440 ;
        RECT 4.400 1053.640 1195.740 1055.040 ;
        RECT 4.000 1041.440 1195.740 1053.640 ;
        RECT 4.000 1040.040 1195.340 1041.440 ;
        RECT 4.000 1034.640 1195.740 1040.040 ;
        RECT 4.400 1033.240 1195.740 1034.640 ;
        RECT 4.000 1021.040 1195.740 1033.240 ;
        RECT 4.000 1019.640 1195.340 1021.040 ;
        RECT 4.000 1014.240 1195.740 1019.640 ;
        RECT 4.400 1012.840 1195.740 1014.240 ;
        RECT 4.000 1000.640 1195.740 1012.840 ;
        RECT 4.000 999.240 1195.340 1000.640 ;
        RECT 4.000 993.840 1195.740 999.240 ;
        RECT 4.400 992.440 1195.740 993.840 ;
        RECT 4.000 980.240 1195.740 992.440 ;
        RECT 4.000 978.840 1195.340 980.240 ;
        RECT 4.000 973.440 1195.740 978.840 ;
        RECT 4.400 972.040 1195.740 973.440 ;
        RECT 4.000 959.840 1195.740 972.040 ;
        RECT 4.000 958.440 1195.340 959.840 ;
        RECT 4.000 953.040 1195.740 958.440 ;
        RECT 4.400 951.640 1195.740 953.040 ;
        RECT 4.000 939.440 1195.740 951.640 ;
        RECT 4.000 938.040 1195.340 939.440 ;
        RECT 4.000 932.640 1195.740 938.040 ;
        RECT 4.400 931.240 1195.740 932.640 ;
        RECT 4.000 919.040 1195.740 931.240 ;
        RECT 4.000 917.640 1195.340 919.040 ;
        RECT 4.000 912.240 1195.740 917.640 ;
        RECT 4.400 910.840 1195.740 912.240 ;
        RECT 4.000 895.240 1195.740 910.840 ;
        RECT 4.000 893.840 1195.340 895.240 ;
        RECT 4.000 888.440 1195.740 893.840 ;
        RECT 4.400 887.040 1195.740 888.440 ;
        RECT 4.000 874.840 1195.740 887.040 ;
        RECT 4.000 873.440 1195.340 874.840 ;
        RECT 4.000 868.040 1195.740 873.440 ;
        RECT 4.400 866.640 1195.740 868.040 ;
        RECT 4.000 854.440 1195.740 866.640 ;
        RECT 4.000 853.040 1195.340 854.440 ;
        RECT 4.000 847.640 1195.740 853.040 ;
        RECT 4.400 846.240 1195.740 847.640 ;
        RECT 4.000 834.040 1195.740 846.240 ;
        RECT 4.000 832.640 1195.340 834.040 ;
        RECT 4.000 827.240 1195.740 832.640 ;
        RECT 4.400 825.840 1195.740 827.240 ;
        RECT 4.000 813.640 1195.740 825.840 ;
        RECT 4.000 812.240 1195.340 813.640 ;
        RECT 4.000 806.840 1195.740 812.240 ;
        RECT 4.400 805.440 1195.740 806.840 ;
        RECT 4.000 793.240 1195.740 805.440 ;
        RECT 4.000 791.840 1195.340 793.240 ;
        RECT 4.000 786.440 1195.740 791.840 ;
        RECT 4.400 785.040 1195.740 786.440 ;
        RECT 4.000 772.840 1195.740 785.040 ;
        RECT 4.000 771.440 1195.340 772.840 ;
        RECT 4.000 766.040 1195.740 771.440 ;
        RECT 4.400 764.640 1195.740 766.040 ;
        RECT 4.000 752.440 1195.740 764.640 ;
        RECT 4.000 751.040 1195.340 752.440 ;
        RECT 4.000 745.640 1195.740 751.040 ;
        RECT 4.400 744.240 1195.740 745.640 ;
        RECT 4.000 732.040 1195.740 744.240 ;
        RECT 4.000 730.640 1195.340 732.040 ;
        RECT 4.000 725.240 1195.740 730.640 ;
        RECT 4.400 723.840 1195.740 725.240 ;
        RECT 4.000 711.640 1195.740 723.840 ;
        RECT 4.000 710.240 1195.340 711.640 ;
        RECT 4.000 704.840 1195.740 710.240 ;
        RECT 4.400 703.440 1195.740 704.840 ;
        RECT 4.000 691.240 1195.740 703.440 ;
        RECT 4.000 689.840 1195.340 691.240 ;
        RECT 4.000 684.440 1195.740 689.840 ;
        RECT 4.400 683.040 1195.740 684.440 ;
        RECT 4.000 670.840 1195.740 683.040 ;
        RECT 4.000 669.440 1195.340 670.840 ;
        RECT 4.000 664.040 1195.740 669.440 ;
        RECT 4.400 662.640 1195.740 664.040 ;
        RECT 4.000 650.440 1195.740 662.640 ;
        RECT 4.000 649.040 1195.340 650.440 ;
        RECT 4.000 643.640 1195.740 649.040 ;
        RECT 4.400 642.240 1195.740 643.640 ;
        RECT 4.000 630.040 1195.740 642.240 ;
        RECT 4.000 628.640 1195.340 630.040 ;
        RECT 4.000 623.240 1195.740 628.640 ;
        RECT 4.400 621.840 1195.740 623.240 ;
        RECT 4.000 606.240 1195.740 621.840 ;
        RECT 4.000 604.840 1195.340 606.240 ;
        RECT 4.000 602.840 1195.740 604.840 ;
        RECT 4.400 601.440 1195.740 602.840 ;
        RECT 4.000 585.840 1195.740 601.440 ;
        RECT 4.000 584.440 1195.340 585.840 ;
        RECT 4.000 579.040 1195.740 584.440 ;
        RECT 4.400 577.640 1195.740 579.040 ;
        RECT 4.000 565.440 1195.740 577.640 ;
        RECT 4.000 564.040 1195.340 565.440 ;
        RECT 4.000 558.640 1195.740 564.040 ;
        RECT 4.400 557.240 1195.740 558.640 ;
        RECT 4.000 545.040 1195.740 557.240 ;
        RECT 4.000 543.640 1195.340 545.040 ;
        RECT 4.000 538.240 1195.740 543.640 ;
        RECT 4.400 536.840 1195.740 538.240 ;
        RECT 4.000 524.640 1195.740 536.840 ;
        RECT 4.000 523.240 1195.340 524.640 ;
        RECT 4.000 517.840 1195.740 523.240 ;
        RECT 4.400 516.440 1195.740 517.840 ;
        RECT 4.000 504.240 1195.740 516.440 ;
        RECT 4.000 502.840 1195.340 504.240 ;
        RECT 4.000 497.440 1195.740 502.840 ;
        RECT 4.400 496.040 1195.740 497.440 ;
        RECT 4.000 483.840 1195.740 496.040 ;
        RECT 4.000 482.440 1195.340 483.840 ;
        RECT 4.000 477.040 1195.740 482.440 ;
        RECT 4.400 475.640 1195.740 477.040 ;
        RECT 4.000 463.440 1195.740 475.640 ;
        RECT 4.000 462.040 1195.340 463.440 ;
        RECT 4.000 456.640 1195.740 462.040 ;
        RECT 4.400 455.240 1195.740 456.640 ;
        RECT 4.000 443.040 1195.740 455.240 ;
        RECT 4.000 441.640 1195.340 443.040 ;
        RECT 4.000 436.240 1195.740 441.640 ;
        RECT 4.400 434.840 1195.740 436.240 ;
        RECT 4.000 422.640 1195.740 434.840 ;
        RECT 4.000 421.240 1195.340 422.640 ;
        RECT 4.000 415.840 1195.740 421.240 ;
        RECT 4.400 414.440 1195.740 415.840 ;
        RECT 4.000 402.240 1195.740 414.440 ;
        RECT 4.000 400.840 1195.340 402.240 ;
        RECT 4.000 395.440 1195.740 400.840 ;
        RECT 4.400 394.040 1195.740 395.440 ;
        RECT 4.000 381.840 1195.740 394.040 ;
        RECT 4.000 380.440 1195.340 381.840 ;
        RECT 4.000 375.040 1195.740 380.440 ;
        RECT 4.400 373.640 1195.740 375.040 ;
        RECT 4.000 361.440 1195.740 373.640 ;
        RECT 4.000 360.040 1195.340 361.440 ;
        RECT 4.000 354.640 1195.740 360.040 ;
        RECT 4.400 353.240 1195.740 354.640 ;
        RECT 4.000 341.040 1195.740 353.240 ;
        RECT 4.000 339.640 1195.340 341.040 ;
        RECT 4.000 334.240 1195.740 339.640 ;
        RECT 4.400 332.840 1195.740 334.240 ;
        RECT 4.000 320.640 1195.740 332.840 ;
        RECT 4.000 319.240 1195.340 320.640 ;
        RECT 4.000 313.840 1195.740 319.240 ;
        RECT 4.400 312.440 1195.740 313.840 ;
        RECT 4.000 296.840 1195.740 312.440 ;
        RECT 4.000 295.440 1195.340 296.840 ;
        RECT 4.000 290.040 1195.740 295.440 ;
        RECT 4.400 288.640 1195.740 290.040 ;
        RECT 4.000 276.440 1195.740 288.640 ;
        RECT 4.000 275.040 1195.340 276.440 ;
        RECT 4.000 269.640 1195.740 275.040 ;
        RECT 4.400 268.240 1195.740 269.640 ;
        RECT 4.000 256.040 1195.740 268.240 ;
        RECT 4.000 254.640 1195.340 256.040 ;
        RECT 4.000 249.240 1195.740 254.640 ;
        RECT 4.400 247.840 1195.740 249.240 ;
        RECT 4.000 235.640 1195.740 247.840 ;
        RECT 4.000 234.240 1195.340 235.640 ;
        RECT 4.000 228.840 1195.740 234.240 ;
        RECT 4.400 227.440 1195.740 228.840 ;
        RECT 4.000 215.240 1195.740 227.440 ;
        RECT 4.000 213.840 1195.340 215.240 ;
        RECT 4.000 208.440 1195.740 213.840 ;
        RECT 4.400 207.040 1195.740 208.440 ;
        RECT 4.000 194.840 1195.740 207.040 ;
        RECT 4.000 193.440 1195.340 194.840 ;
        RECT 4.000 188.040 1195.740 193.440 ;
        RECT 4.400 186.640 1195.740 188.040 ;
        RECT 4.000 174.440 1195.740 186.640 ;
        RECT 4.000 173.040 1195.340 174.440 ;
        RECT 4.000 167.640 1195.740 173.040 ;
        RECT 4.400 166.240 1195.740 167.640 ;
        RECT 4.000 154.040 1195.740 166.240 ;
        RECT 4.000 152.640 1195.340 154.040 ;
        RECT 4.000 147.240 1195.740 152.640 ;
        RECT 4.400 145.840 1195.740 147.240 ;
        RECT 4.000 133.640 1195.740 145.840 ;
        RECT 4.000 132.240 1195.340 133.640 ;
        RECT 4.000 126.840 1195.740 132.240 ;
        RECT 4.400 125.440 1195.740 126.840 ;
        RECT 4.000 113.240 1195.740 125.440 ;
        RECT 4.000 111.840 1195.340 113.240 ;
        RECT 4.000 106.440 1195.740 111.840 ;
        RECT 4.400 105.040 1195.740 106.440 ;
        RECT 4.000 92.840 1195.740 105.040 ;
        RECT 4.000 91.440 1195.340 92.840 ;
        RECT 4.000 86.040 1195.740 91.440 ;
        RECT 4.400 84.640 1195.740 86.040 ;
        RECT 4.000 72.440 1195.740 84.640 ;
        RECT 4.000 71.040 1195.340 72.440 ;
        RECT 4.000 65.640 1195.740 71.040 ;
        RECT 4.400 64.240 1195.740 65.640 ;
        RECT 4.000 52.040 1195.740 64.240 ;
        RECT 4.000 50.640 1195.340 52.040 ;
        RECT 4.000 45.240 1195.740 50.640 ;
        RECT 4.400 43.840 1195.740 45.240 ;
        RECT 4.000 31.640 1195.740 43.840 ;
        RECT 4.000 30.240 1195.340 31.640 ;
        RECT 4.000 24.840 1195.740 30.240 ;
        RECT 4.400 23.440 1195.740 24.840 ;
        RECT 4.000 7.840 1195.740 23.440 ;
        RECT 4.000 6.975 1195.340 7.840 ;
      LAYER met4 ;
        RECT 95.055 1200.160 1076.105 1202.745 ;
        RECT 95.055 501.860 95.640 1200.160 ;
        RECT 98.040 501.860 120.640 1200.160 ;
        RECT 123.040 501.860 145.640 1200.160 ;
        RECT 148.040 501.860 170.640 1200.160 ;
        RECT 173.040 501.860 195.640 1200.160 ;
        RECT 198.040 501.860 220.640 1200.160 ;
        RECT 223.040 501.860 245.640 1200.160 ;
        RECT 248.040 501.860 270.640 1200.160 ;
        RECT 273.040 501.860 295.640 1200.160 ;
        RECT 298.040 501.860 320.640 1200.160 ;
        RECT 323.040 501.860 345.640 1200.160 ;
        RECT 348.040 501.860 370.640 1200.160 ;
        RECT 373.040 501.860 395.640 1200.160 ;
        RECT 398.040 501.860 420.640 1200.160 ;
        RECT 423.040 501.860 445.640 1200.160 ;
        RECT 448.040 501.860 470.640 1200.160 ;
        RECT 473.040 501.860 495.640 1200.160 ;
        RECT 498.040 501.860 520.640 1200.160 ;
        RECT 523.040 501.860 545.640 1200.160 ;
        RECT 548.040 501.860 570.640 1200.160 ;
        RECT 573.040 501.860 595.640 1200.160 ;
        RECT 95.055 95.640 595.640 501.860 ;
        RECT 95.055 10.240 95.640 95.640 ;
        RECT 98.040 10.240 120.640 95.640 ;
        RECT 123.040 10.240 145.640 95.640 ;
        RECT 148.040 10.240 170.640 95.640 ;
        RECT 173.040 10.240 195.640 95.640 ;
        RECT 198.040 10.240 220.640 95.640 ;
        RECT 223.040 10.240 245.640 95.640 ;
        RECT 248.040 10.240 270.640 95.640 ;
        RECT 273.040 10.240 295.640 95.640 ;
        RECT 298.040 10.240 320.640 95.640 ;
        RECT 323.040 10.240 345.640 95.640 ;
        RECT 348.040 10.240 370.640 95.640 ;
        RECT 373.040 10.240 395.640 95.640 ;
        RECT 398.040 10.240 420.640 95.640 ;
        RECT 423.040 10.240 445.640 95.640 ;
        RECT 448.040 10.240 470.640 95.640 ;
        RECT 473.040 10.240 495.640 95.640 ;
        RECT 498.040 10.240 520.640 95.640 ;
        RECT 523.040 10.240 545.640 95.640 ;
        RECT 548.040 10.240 570.640 95.640 ;
        RECT 573.040 10.240 595.640 95.640 ;
        RECT 598.040 10.240 620.640 1200.160 ;
        RECT 623.040 10.240 645.640 1200.160 ;
        RECT 648.040 10.240 670.640 1200.160 ;
        RECT 673.040 10.240 695.640 1200.160 ;
        RECT 698.040 10.240 720.640 1200.160 ;
        RECT 723.040 10.240 745.640 1200.160 ;
        RECT 748.040 10.240 770.640 1200.160 ;
        RECT 773.040 10.240 795.640 1200.160 ;
        RECT 798.040 10.240 820.640 1200.160 ;
        RECT 823.040 10.240 845.640 1200.160 ;
        RECT 848.040 10.240 870.640 1200.160 ;
        RECT 873.040 10.240 895.640 1200.160 ;
        RECT 898.040 10.240 920.640 1200.160 ;
        RECT 923.040 10.240 945.640 1200.160 ;
        RECT 948.040 10.240 970.640 1200.160 ;
        RECT 973.040 10.240 995.640 1200.160 ;
        RECT 998.040 10.240 1020.640 1200.160 ;
        RECT 1023.040 10.240 1045.640 1200.160 ;
        RECT 1048.040 10.240 1070.640 1200.160 ;
        RECT 1073.040 10.240 1076.105 1200.160 ;
        RECT 95.055 9.015 1076.105 10.240 ;
  END
END user_proj_example
END LIBRARY

